module fpga (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    VPWR,
    VGND,
    gpio_east,
    gpio_north,
    gpio_south,
    gpio_west,
    wbs_addr_i,
    wbs_data_i,
    wbs_data_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input VPWR;
 input VGND;
 inout [9:0] gpio_east;
 inout [9:0] gpio_north;
 inout [7:0] gpio_south;
 inout [9:0] gpio_west;
 input [31:0] wbs_addr_i;
 input [31:0] wbs_data_i;
 output [31:0] wbs_data_o;
 input [3:0] wbs_sel_i;

 clb_tile \X[0].Y[0].clb  (.carry_in(_000_),
    .carry_out(\carry[1][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[0][0] ),
    .set_out_hard(\col_set[1][0] ),
    .shift_in_hard(\wb_shift_out[0][0] ),
    .shift_out_hard(\col_shift[1][0] ),
    .cb_east_in({\dc_ew[1][4] ,
    \dc_ew[1][3] ,
    \dc_ew[1][2] ,
    \dc_ew[1][1] ,
    \dc_ew[1][0] }),
    .cb_east_out({\dc_we[1][9] ,
    \dc_we[1][8] ,
    \dc_we[1][7] ,
    \dc_we[1][6] ,
    \dc_we[1][5] ,
    \dc_we[1][4] ,
    \dc_we[1][3] ,
    \dc_we[1][2] ,
    \dc_we[1][1] ,
    \dc_we[1][0] }),
    .cb_north_in({\dc_ns[7][4] ,
    \dc_ns[7][3] ,
    \dc_ns[7][2] ,
    \dc_ns[7][1] ,
    \dc_ns[7][0] }),
    .cb_north_out({\dc_sn[7][9] ,
    \dc_sn[7][8] ,
    \dc_sn[7][7] ,
    \dc_sn[7][6] ,
    \dc_sn[7][5] ,
    \dc_sn[7][4] ,
    \dc_sn[7][3] ,
    \dc_sn[7][2] ,
    \dc_sn[7][1] ,
    \dc_sn[7][0] }),
    .clb_south_in({_010_,
    _009_,
    _008_,
    _007_,
    _006_,
    _005_,
    _004_,
    _003_,
    _002_,
    _001_}),
    .clb_south_out({\dc_ns[0][4] ,
    \dc_ns[0][3] ,
    \dc_ns[0][2] ,
    \dc_ns[0][1] ,
    \dc_ns[0][0] }),
    .clb_west_in({_020_,
    _019_,
    _018_,
    _017_,
    _016_,
    _015_,
    _014_,
    _013_,
    _012_,
    _011_}),
    .clb_west_out({\dc_ew[0][4] ,
    \dc_ew[0][3] ,
    \dc_ew[0][2] ,
    \dc_ew[0][1] ,
    \dc_ew[0][0] }),
    .east_double({\ix_double_ew[1][7] ,
    \ix_double_ew[1][6] ,
    \ix_double_ew[1][5] ,
    \ix_double_ew[1][4] ,
    \ix_double_ew[1][3] ,
    \ix_double_ew[1][2] ,
    \ix_double_ew[1][1] ,
    \ix_double_ew[1][0] }),
    .east_single({\ix_single_ew[1][3] ,
    \ix_single_ew[1][2] ,
    \ix_single_ew[1][1] ,
    \ix_single_ew[1][0] }),
    .north_double({\ix_double_ns[7][7] ,
    \ix_double_ns[7][6] ,
    \ix_double_ns[7][5] ,
    \ix_double_ns[7][4] ,
    \ix_double_ns[7][3] ,
    \ix_double_ns[7][2] ,
    \ix_double_ns[7][1] ,
    \ix_double_ns[7][0] }),
    .north_single({\ix_single_ns[7][3] ,
    \ix_single_ns[7][2] ,
    \ix_single_ns[7][1] ,
    \ix_single_ns[7][0] }),
    .south_double({\ix_double_ns[0][7] ,
    \ix_double_ns[0][6] ,
    \ix_double_ns[0][5] ,
    \ix_double_ns[0][4] ,
    \ix_double_ns[0][3] ,
    \ix_double_ns[0][2] ,
    \ix_double_ns[0][1] ,
    \ix_double_ns[0][0] }),
    .south_single({\ix_single_ns[0][3] ,
    \ix_single_ns[0][2] ,
    \ix_single_ns[0][1] ,
    gpio_south[0]}),
    .west_double({\ix_double_ew[0][7] ,
    \ix_double_ew[0][6] ,
    \ix_double_ew[0][5] ,
    \ix_double_ew[0][4] ,
    \ix_double_ew[0][3] ,
    \ix_double_ew[0][2] ,
    \ix_double_ew[0][1] ,
    \ix_double_ew[0][0] }),
    .west_single({\ix_single_ew[0][3] ,
    \ix_single_ew[0][2] ,
    \ix_single_ew[0][1] ,
    gpio_west[0]}));
 clb_tile \X[0].Y[1].clb  (.carry_in(\carry[1][0] ),
    .carry_out(\carry[2][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][0] ),
    .set_out_hard(\col_set[2][0] ),
    .shift_in_hard(\col_shift[1][0] ),
    .shift_out_hard(\col_shift[2][0] ),
    .cb_east_in({\dc_ew[9][4] ,
    \dc_ew[9][3] ,
    \dc_ew[9][2] ,
    \dc_ew[9][1] ,
    \dc_ew[9][0] }),
    .cb_east_out({\dc_we[9][9] ,
    \dc_we[9][8] ,
    \dc_we[9][7] ,
    \dc_we[9][6] ,
    \dc_we[9][5] ,
    \dc_we[9][4] ,
    \dc_we[9][3] ,
    \dc_we[9][2] ,
    \dc_we[9][1] ,
    \dc_we[9][0] }),
    .cb_north_in({\dc_ns[14][4] ,
    \dc_ns[14][3] ,
    \dc_ns[14][2] ,
    \dc_ns[14][1] ,
    \dc_ns[14][0] }),
    .cb_north_out({\dc_sn[14][9] ,
    \dc_sn[14][8] ,
    \dc_sn[14][7] ,
    \dc_sn[14][6] ,
    \dc_sn[14][5] ,
    \dc_sn[14][4] ,
    \dc_sn[14][3] ,
    \dc_sn[14][2] ,
    \dc_sn[14][1] ,
    \dc_sn[14][0] }),
    .clb_south_in({\dc_sn[7][9] ,
    \dc_sn[7][8] ,
    \dc_sn[7][7] ,
    \dc_sn[7][6] ,
    \dc_sn[7][5] ,
    \dc_sn[7][4] ,
    \dc_sn[7][3] ,
    \dc_sn[7][2] ,
    \dc_sn[7][1] ,
    \dc_sn[7][0] }),
    .clb_south_out({\dc_ns[7][4] ,
    \dc_ns[7][3] ,
    \dc_ns[7][2] ,
    \dc_ns[7][1] ,
    \dc_ns[7][0] }),
    .clb_west_in({_030_,
    _029_,
    _028_,
    _027_,
    _026_,
    _025_,
    _024_,
    _023_,
    _022_,
    _021_}),
    .clb_west_out({\dc_ew[8][4] ,
    \dc_ew[8][3] ,
    \dc_ew[8][2] ,
    \dc_ew[8][1] ,
    \dc_ew[8][0] }),
    .east_double({\ix_double_ew[9][7] ,
    \ix_double_ew[9][6] ,
    \ix_double_ew[9][5] ,
    \ix_double_ew[9][4] ,
    \ix_double_ew[9][3] ,
    \ix_double_ew[9][2] ,
    \ix_double_ew[9][1] ,
    \ix_double_ew[9][0] }),
    .east_single({\ix_single_ew[9][3] ,
    \ix_single_ew[9][2] ,
    \ix_single_ew[9][1] ,
    \ix_single_ew[9][0] }),
    .north_double({\ix_double_ns[14][7] ,
    \ix_double_ns[14][6] ,
    \ix_double_ns[14][5] ,
    \ix_double_ns[14][4] ,
    \ix_double_ns[14][3] ,
    \ix_double_ns[14][2] ,
    \ix_double_ns[14][1] ,
    \ix_double_ns[14][0] }),
    .north_single({\ix_single_ns[14][3] ,
    \ix_single_ns[14][2] ,
    \ix_single_ns[14][1] ,
    \ix_single_ns[14][0] }),
    .south_double({\ix_double_ns[7][7] ,
    \ix_double_ns[7][6] ,
    \ix_double_ns[7][5] ,
    \ix_double_ns[7][4] ,
    \ix_double_ns[7][3] ,
    \ix_double_ns[7][2] ,
    \ix_double_ns[7][1] ,
    \ix_double_ns[7][0] }),
    .south_single({\ix_single_ns[7][3] ,
    \ix_single_ns[7][2] ,
    \ix_single_ns[7][1] ,
    \ix_single_ns[7][0] }),
    .west_double({\ix_double_ew[8][7] ,
    \ix_double_ew[8][6] ,
    \ix_double_ew[8][5] ,
    \ix_double_ew[8][4] ,
    \ix_double_ew[8][3] ,
    \ix_double_ew[8][2] ,
    \ix_double_ew[8][1] ,
    \ix_double_ew[8][0] }),
    .west_single({\ix_single_ew[8][3] ,
    \ix_single_ew[8][2] ,
    \ix_single_ew[8][1] ,
    gpio_west[1]}));
 clb_tile \X[0].Y[2].clb  (.carry_in(\carry[2][0] ),
    .carry_out(\carry[3][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][0] ),
    .set_out_hard(\col_set[3][0] ),
    .shift_in_hard(\col_shift[2][0] ),
    .shift_out_hard(\col_shift[3][0] ),
    .cb_east_in({\dc_ew[17][4] ,
    \dc_ew[17][3] ,
    \dc_ew[17][2] ,
    \dc_ew[17][1] ,
    \dc_ew[17][0] }),
    .cb_east_out({\dc_we[17][9] ,
    \dc_we[17][8] ,
    \dc_we[17][7] ,
    \dc_we[17][6] ,
    \dc_we[17][5] ,
    \dc_we[17][4] ,
    \dc_we[17][3] ,
    \dc_we[17][2] ,
    \dc_we[17][1] ,
    \dc_we[17][0] }),
    .cb_north_in({\dc_ns[21][4] ,
    \dc_ns[21][3] ,
    \dc_ns[21][2] ,
    \dc_ns[21][1] ,
    \dc_ns[21][0] }),
    .cb_north_out({\dc_sn[21][9] ,
    \dc_sn[21][8] ,
    \dc_sn[21][7] ,
    \dc_sn[21][6] ,
    \dc_sn[21][5] ,
    \dc_sn[21][4] ,
    \dc_sn[21][3] ,
    \dc_sn[21][2] ,
    \dc_sn[21][1] ,
    \dc_sn[21][0] }),
    .clb_south_in({\dc_sn[14][9] ,
    \dc_sn[14][8] ,
    \dc_sn[14][7] ,
    \dc_sn[14][6] ,
    \dc_sn[14][5] ,
    \dc_sn[14][4] ,
    \dc_sn[14][3] ,
    \dc_sn[14][2] ,
    \dc_sn[14][1] ,
    \dc_sn[14][0] }),
    .clb_south_out({\dc_ns[14][4] ,
    \dc_ns[14][3] ,
    \dc_ns[14][2] ,
    \dc_ns[14][1] ,
    \dc_ns[14][0] }),
    .clb_west_in({_040_,
    _039_,
    _038_,
    _037_,
    _036_,
    _035_,
    _034_,
    _033_,
    _032_,
    _031_}),
    .clb_west_out({\dc_ew[16][4] ,
    \dc_ew[16][3] ,
    \dc_ew[16][2] ,
    \dc_ew[16][1] ,
    \dc_ew[16][0] }),
    .east_double({\ix_double_ew[17][7] ,
    \ix_double_ew[17][6] ,
    \ix_double_ew[17][5] ,
    \ix_double_ew[17][4] ,
    \ix_double_ew[17][3] ,
    \ix_double_ew[17][2] ,
    \ix_double_ew[17][1] ,
    \ix_double_ew[17][0] }),
    .east_single({\ix_single_ew[17][3] ,
    \ix_single_ew[17][2] ,
    \ix_single_ew[17][1] ,
    \ix_single_ew[17][0] }),
    .north_double({\ix_double_ns[21][7] ,
    \ix_double_ns[21][6] ,
    \ix_double_ns[21][5] ,
    \ix_double_ns[21][4] ,
    \ix_double_ns[21][3] ,
    \ix_double_ns[21][2] ,
    \ix_double_ns[21][1] ,
    \ix_double_ns[21][0] }),
    .north_single({\ix_single_ns[21][3] ,
    \ix_single_ns[21][2] ,
    \ix_single_ns[21][1] ,
    \ix_single_ns[21][0] }),
    .south_double({\ix_double_ns[14][7] ,
    \ix_double_ns[14][6] ,
    \ix_double_ns[14][5] ,
    \ix_double_ns[14][4] ,
    \ix_double_ns[14][3] ,
    \ix_double_ns[14][2] ,
    \ix_double_ns[14][1] ,
    \ix_double_ns[14][0] }),
    .south_single({\ix_single_ns[14][3] ,
    \ix_single_ns[14][2] ,
    \ix_single_ns[14][1] ,
    \ix_single_ns[14][0] }),
    .west_double({\ix_double_ew[16][7] ,
    \ix_double_ew[16][6] ,
    \ix_double_ew[16][5] ,
    \ix_double_ew[16][4] ,
    \ix_double_ew[16][3] ,
    \ix_double_ew[16][2] ,
    \ix_double_ew[16][1] ,
    \ix_double_ew[16][0] }),
    .west_single({\ix_single_ew[16][3] ,
    \ix_single_ew[16][2] ,
    \ix_single_ew[16][1] ,
    gpio_west[2]}));
 clb_tile \X[0].Y[3].clb  (.carry_in(\carry[3][0] ),
    .carry_out(\carry[4][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][0] ),
    .set_out_hard(\col_set[4][0] ),
    .shift_in_hard(\col_shift[3][0] ),
    .shift_out_hard(\col_shift[4][0] ),
    .cb_east_in({\dc_ew[25][4] ,
    \dc_ew[25][3] ,
    \dc_ew[25][2] ,
    \dc_ew[25][1] ,
    \dc_ew[25][0] }),
    .cb_east_out({\dc_we[25][9] ,
    \dc_we[25][8] ,
    \dc_we[25][7] ,
    \dc_we[25][6] ,
    \dc_we[25][5] ,
    \dc_we[25][4] ,
    \dc_we[25][3] ,
    \dc_we[25][2] ,
    \dc_we[25][1] ,
    \dc_we[25][0] }),
    .cb_north_in({\dc_ns[28][4] ,
    \dc_ns[28][3] ,
    \dc_ns[28][2] ,
    \dc_ns[28][1] ,
    \dc_ns[28][0] }),
    .cb_north_out({\dc_sn[28][9] ,
    \dc_sn[28][8] ,
    \dc_sn[28][7] ,
    \dc_sn[28][6] ,
    \dc_sn[28][5] ,
    \dc_sn[28][4] ,
    \dc_sn[28][3] ,
    \dc_sn[28][2] ,
    \dc_sn[28][1] ,
    \dc_sn[28][0] }),
    .clb_south_in({\dc_sn[21][9] ,
    \dc_sn[21][8] ,
    \dc_sn[21][7] ,
    \dc_sn[21][6] ,
    \dc_sn[21][5] ,
    \dc_sn[21][4] ,
    \dc_sn[21][3] ,
    \dc_sn[21][2] ,
    \dc_sn[21][1] ,
    \dc_sn[21][0] }),
    .clb_south_out({\dc_ns[21][4] ,
    \dc_ns[21][3] ,
    \dc_ns[21][2] ,
    \dc_ns[21][1] ,
    \dc_ns[21][0] }),
    .clb_west_in({_050_,
    _049_,
    _048_,
    _047_,
    _046_,
    _045_,
    _044_,
    _043_,
    _042_,
    _041_}),
    .clb_west_out({\dc_ew[24][4] ,
    \dc_ew[24][3] ,
    \dc_ew[24][2] ,
    \dc_ew[24][1] ,
    \dc_ew[24][0] }),
    .east_double({\ix_double_ew[25][7] ,
    \ix_double_ew[25][6] ,
    \ix_double_ew[25][5] ,
    \ix_double_ew[25][4] ,
    \ix_double_ew[25][3] ,
    \ix_double_ew[25][2] ,
    \ix_double_ew[25][1] ,
    \ix_double_ew[25][0] }),
    .east_single({\ix_single_ew[25][3] ,
    \ix_single_ew[25][2] ,
    \ix_single_ew[25][1] ,
    \ix_single_ew[25][0] }),
    .north_double({\ix_double_ns[28][7] ,
    \ix_double_ns[28][6] ,
    \ix_double_ns[28][5] ,
    \ix_double_ns[28][4] ,
    \ix_double_ns[28][3] ,
    \ix_double_ns[28][2] ,
    \ix_double_ns[28][1] ,
    \ix_double_ns[28][0] }),
    .north_single({\ix_single_ns[28][3] ,
    \ix_single_ns[28][2] ,
    \ix_single_ns[28][1] ,
    \ix_single_ns[28][0] }),
    .south_double({\ix_double_ns[21][7] ,
    \ix_double_ns[21][6] ,
    \ix_double_ns[21][5] ,
    \ix_double_ns[21][4] ,
    \ix_double_ns[21][3] ,
    \ix_double_ns[21][2] ,
    \ix_double_ns[21][1] ,
    \ix_double_ns[21][0] }),
    .south_single({\ix_single_ns[21][3] ,
    \ix_single_ns[21][2] ,
    \ix_single_ns[21][1] ,
    \ix_single_ns[21][0] }),
    .west_double({\ix_double_ew[24][7] ,
    \ix_double_ew[24][6] ,
    \ix_double_ew[24][5] ,
    \ix_double_ew[24][4] ,
    \ix_double_ew[24][3] ,
    \ix_double_ew[24][2] ,
    \ix_double_ew[24][1] ,
    \ix_double_ew[24][0] }),
    .west_single({\ix_single_ew[24][3] ,
    \ix_single_ew[24][2] ,
    \ix_single_ew[24][1] ,
    gpio_west[3]}));
 clb_tile \X[0].Y[4].clb  (.carry_in(\carry[4][0] ),
    .carry_out(\carry[5][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][0] ),
    .set_out_hard(\col_set[5][0] ),
    .shift_in_hard(\col_shift[4][0] ),
    .shift_out_hard(\col_shift[5][0] ),
    .cb_east_in({\dc_ew[33][4] ,
    \dc_ew[33][3] ,
    \dc_ew[33][2] ,
    \dc_ew[33][1] ,
    \dc_ew[33][0] }),
    .cb_east_out({\dc_we[33][9] ,
    \dc_we[33][8] ,
    \dc_we[33][7] ,
    \dc_we[33][6] ,
    \dc_we[33][5] ,
    \dc_we[33][4] ,
    \dc_we[33][3] ,
    \dc_we[33][2] ,
    \dc_we[33][1] ,
    \dc_we[33][0] }),
    .cb_north_in({\dc_ns[35][4] ,
    \dc_ns[35][3] ,
    \dc_ns[35][2] ,
    \dc_ns[35][1] ,
    \dc_ns[35][0] }),
    .cb_north_out({\dc_sn[35][9] ,
    \dc_sn[35][8] ,
    \dc_sn[35][7] ,
    \dc_sn[35][6] ,
    \dc_sn[35][5] ,
    \dc_sn[35][4] ,
    \dc_sn[35][3] ,
    \dc_sn[35][2] ,
    \dc_sn[35][1] ,
    \dc_sn[35][0] }),
    .clb_south_in({\dc_sn[28][9] ,
    \dc_sn[28][8] ,
    \dc_sn[28][7] ,
    \dc_sn[28][6] ,
    \dc_sn[28][5] ,
    \dc_sn[28][4] ,
    \dc_sn[28][3] ,
    \dc_sn[28][2] ,
    \dc_sn[28][1] ,
    \dc_sn[28][0] }),
    .clb_south_out({\dc_ns[28][4] ,
    \dc_ns[28][3] ,
    \dc_ns[28][2] ,
    \dc_ns[28][1] ,
    \dc_ns[28][0] }),
    .clb_west_in({_060_,
    _059_,
    _058_,
    _057_,
    _056_,
    _055_,
    _054_,
    _053_,
    _052_,
    _051_}),
    .clb_west_out({\dc_ew[32][4] ,
    \dc_ew[32][3] ,
    \dc_ew[32][2] ,
    \dc_ew[32][1] ,
    \dc_ew[32][0] }),
    .east_double({\ix_double_ew[33][7] ,
    \ix_double_ew[33][6] ,
    \ix_double_ew[33][5] ,
    \ix_double_ew[33][4] ,
    \ix_double_ew[33][3] ,
    \ix_double_ew[33][2] ,
    \ix_double_ew[33][1] ,
    \ix_double_ew[33][0] }),
    .east_single({\ix_single_ew[33][3] ,
    \ix_single_ew[33][2] ,
    \ix_single_ew[33][1] ,
    \ix_single_ew[33][0] }),
    .north_double({\ix_double_ns[35][7] ,
    \ix_double_ns[35][6] ,
    \ix_double_ns[35][5] ,
    \ix_double_ns[35][4] ,
    \ix_double_ns[35][3] ,
    \ix_double_ns[35][2] ,
    \ix_double_ns[35][1] ,
    \ix_double_ns[35][0] }),
    .north_single({\ix_single_ns[35][3] ,
    \ix_single_ns[35][2] ,
    \ix_single_ns[35][1] ,
    \ix_single_ns[35][0] }),
    .south_double({\ix_double_ns[28][7] ,
    \ix_double_ns[28][6] ,
    \ix_double_ns[28][5] ,
    \ix_double_ns[28][4] ,
    \ix_double_ns[28][3] ,
    \ix_double_ns[28][2] ,
    \ix_double_ns[28][1] ,
    \ix_double_ns[28][0] }),
    .south_single({\ix_single_ns[28][3] ,
    \ix_single_ns[28][2] ,
    \ix_single_ns[28][1] ,
    \ix_single_ns[28][0] }),
    .west_double({\ix_double_ew[32][7] ,
    \ix_double_ew[32][6] ,
    \ix_double_ew[32][5] ,
    \ix_double_ew[32][4] ,
    \ix_double_ew[32][3] ,
    \ix_double_ew[32][2] ,
    \ix_double_ew[32][1] ,
    \ix_double_ew[32][0] }),
    .west_single({\ix_single_ew[32][3] ,
    \ix_single_ew[32][2] ,
    \ix_single_ew[32][1] ,
    gpio_west[4]}));
 clb_tile \X[0].Y[5].clb  (.carry_in(\carry[5][0] ),
    .carry_out(\carry[6][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][0] ),
    .set_out_hard(\col_set[6][0] ),
    .shift_in_hard(\col_shift[5][0] ),
    .shift_out_hard(\col_shift[6][0] ),
    .cb_east_in({\dc_ew[41][4] ,
    \dc_ew[41][3] ,
    \dc_ew[41][2] ,
    \dc_ew[41][1] ,
    \dc_ew[41][0] }),
    .cb_east_out({\dc_we[41][9] ,
    \dc_we[41][8] ,
    \dc_we[41][7] ,
    \dc_we[41][6] ,
    \dc_we[41][5] ,
    \dc_we[41][4] ,
    \dc_we[41][3] ,
    \dc_we[41][2] ,
    \dc_we[41][1] ,
    \dc_we[41][0] }),
    .cb_north_in({\dc_ns[42][4] ,
    \dc_ns[42][3] ,
    \dc_ns[42][2] ,
    \dc_ns[42][1] ,
    \dc_ns[42][0] }),
    .cb_north_out({\dc_sn[42][9] ,
    \dc_sn[42][8] ,
    \dc_sn[42][7] ,
    \dc_sn[42][6] ,
    \dc_sn[42][5] ,
    \dc_sn[42][4] ,
    \dc_sn[42][3] ,
    \dc_sn[42][2] ,
    \dc_sn[42][1] ,
    \dc_sn[42][0] }),
    .clb_south_in({\dc_sn[35][9] ,
    \dc_sn[35][8] ,
    \dc_sn[35][7] ,
    \dc_sn[35][6] ,
    \dc_sn[35][5] ,
    \dc_sn[35][4] ,
    \dc_sn[35][3] ,
    \dc_sn[35][2] ,
    \dc_sn[35][1] ,
    \dc_sn[35][0] }),
    .clb_south_out({\dc_ns[35][4] ,
    \dc_ns[35][3] ,
    \dc_ns[35][2] ,
    \dc_ns[35][1] ,
    \dc_ns[35][0] }),
    .clb_west_in({_070_,
    _069_,
    _068_,
    _067_,
    _066_,
    _065_,
    _064_,
    _063_,
    _062_,
    _061_}),
    .clb_west_out({\dc_ew[40][4] ,
    \dc_ew[40][3] ,
    \dc_ew[40][2] ,
    \dc_ew[40][1] ,
    \dc_ew[40][0] }),
    .east_double({\ix_double_ew[41][7] ,
    \ix_double_ew[41][6] ,
    \ix_double_ew[41][5] ,
    \ix_double_ew[41][4] ,
    \ix_double_ew[41][3] ,
    \ix_double_ew[41][2] ,
    \ix_double_ew[41][1] ,
    \ix_double_ew[41][0] }),
    .east_single({\ix_single_ew[41][3] ,
    \ix_single_ew[41][2] ,
    \ix_single_ew[41][1] ,
    \ix_single_ew[41][0] }),
    .north_double({\ix_double_ns[42][7] ,
    \ix_double_ns[42][6] ,
    \ix_double_ns[42][5] ,
    \ix_double_ns[42][4] ,
    \ix_double_ns[42][3] ,
    \ix_double_ns[42][2] ,
    \ix_double_ns[42][1] ,
    \ix_double_ns[42][0] }),
    .north_single({\ix_single_ns[42][3] ,
    \ix_single_ns[42][2] ,
    \ix_single_ns[42][1] ,
    \ix_single_ns[42][0] }),
    .south_double({\ix_double_ns[35][7] ,
    \ix_double_ns[35][6] ,
    \ix_double_ns[35][5] ,
    \ix_double_ns[35][4] ,
    \ix_double_ns[35][3] ,
    \ix_double_ns[35][2] ,
    \ix_double_ns[35][1] ,
    \ix_double_ns[35][0] }),
    .south_single({\ix_single_ns[35][3] ,
    \ix_single_ns[35][2] ,
    \ix_single_ns[35][1] ,
    \ix_single_ns[35][0] }),
    .west_double({\ix_double_ew[40][7] ,
    \ix_double_ew[40][6] ,
    \ix_double_ew[40][5] ,
    \ix_double_ew[40][4] ,
    \ix_double_ew[40][3] ,
    \ix_double_ew[40][2] ,
    \ix_double_ew[40][1] ,
    \ix_double_ew[40][0] }),
    .west_single({\ix_single_ew[40][3] ,
    \ix_single_ew[40][2] ,
    \ix_single_ew[40][1] ,
    gpio_west[5]}));
 clb_tile \X[0].Y[6].clb  (.carry_in(\carry[6][0] ),
    .carry_out(\carry[7][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][0] ),
    .set_out_hard(\col_set[7][0] ),
    .shift_in_hard(\col_shift[6][0] ),
    .shift_out_hard(\col_shift[7][0] ),
    .cb_east_in({\dc_ew[49][4] ,
    \dc_ew[49][3] ,
    \dc_ew[49][2] ,
    \dc_ew[49][1] ,
    \dc_ew[49][0] }),
    .cb_east_out({\dc_we[49][9] ,
    \dc_we[49][8] ,
    \dc_we[49][7] ,
    \dc_we[49][6] ,
    \dc_we[49][5] ,
    \dc_we[49][4] ,
    \dc_we[49][3] ,
    \dc_we[49][2] ,
    \dc_we[49][1] ,
    \dc_we[49][0] }),
    .cb_north_in({\dc_ns[49][4] ,
    \dc_ns[49][3] ,
    \dc_ns[49][2] ,
    \dc_ns[49][1] ,
    \dc_ns[49][0] }),
    .cb_north_out({\dc_sn[49][9] ,
    \dc_sn[49][8] ,
    \dc_sn[49][7] ,
    \dc_sn[49][6] ,
    \dc_sn[49][5] ,
    \dc_sn[49][4] ,
    \dc_sn[49][3] ,
    \dc_sn[49][2] ,
    \dc_sn[49][1] ,
    \dc_sn[49][0] }),
    .clb_south_in({\dc_sn[42][9] ,
    \dc_sn[42][8] ,
    \dc_sn[42][7] ,
    \dc_sn[42][6] ,
    \dc_sn[42][5] ,
    \dc_sn[42][4] ,
    \dc_sn[42][3] ,
    \dc_sn[42][2] ,
    \dc_sn[42][1] ,
    \dc_sn[42][0] }),
    .clb_south_out({\dc_ns[42][4] ,
    \dc_ns[42][3] ,
    \dc_ns[42][2] ,
    \dc_ns[42][1] ,
    \dc_ns[42][0] }),
    .clb_west_in({_080_,
    _079_,
    _078_,
    _077_,
    _076_,
    _075_,
    _074_,
    _073_,
    _072_,
    _071_}),
    .clb_west_out({\dc_ew[48][4] ,
    \dc_ew[48][3] ,
    \dc_ew[48][2] ,
    \dc_ew[48][1] ,
    \dc_ew[48][0] }),
    .east_double({\ix_double_ew[49][7] ,
    \ix_double_ew[49][6] ,
    \ix_double_ew[49][5] ,
    \ix_double_ew[49][4] ,
    \ix_double_ew[49][3] ,
    \ix_double_ew[49][2] ,
    \ix_double_ew[49][1] ,
    \ix_double_ew[49][0] }),
    .east_single({\ix_single_ew[49][3] ,
    \ix_single_ew[49][2] ,
    \ix_single_ew[49][1] ,
    \ix_single_ew[49][0] }),
    .north_double({\ix_double_ns[49][7] ,
    \ix_double_ns[49][6] ,
    \ix_double_ns[49][5] ,
    \ix_double_ns[49][4] ,
    \ix_double_ns[49][3] ,
    \ix_double_ns[49][2] ,
    \ix_double_ns[49][1] ,
    \ix_double_ns[49][0] }),
    .north_single({\ix_single_ns[49][3] ,
    \ix_single_ns[49][2] ,
    \ix_single_ns[49][1] ,
    \ix_single_ns[49][0] }),
    .south_double({\ix_double_ns[42][7] ,
    \ix_double_ns[42][6] ,
    \ix_double_ns[42][5] ,
    \ix_double_ns[42][4] ,
    \ix_double_ns[42][3] ,
    \ix_double_ns[42][2] ,
    \ix_double_ns[42][1] ,
    \ix_double_ns[42][0] }),
    .south_single({\ix_single_ns[42][3] ,
    \ix_single_ns[42][2] ,
    \ix_single_ns[42][1] ,
    \ix_single_ns[42][0] }),
    .west_double({\ix_double_ew[48][7] ,
    \ix_double_ew[48][6] ,
    \ix_double_ew[48][5] ,
    \ix_double_ew[48][4] ,
    \ix_double_ew[48][3] ,
    \ix_double_ew[48][2] ,
    \ix_double_ew[48][1] ,
    \ix_double_ew[48][0] }),
    .west_single({\ix_single_ew[48][3] ,
    \ix_single_ew[48][2] ,
    \ix_single_ew[48][1] ,
    gpio_west[6]}));
 clb_tile \X[0].Y[7].clb  (.carry_in(\carry[7][0] ),
    .carry_out(\carry[8][0] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][0] ),
    .set_out_hard(\col_set[8][0] ),
    .shift_in_hard(\col_shift[7][0] ),
    .shift_out_hard(\col_shift[8][0] ),
    .cb_east_in({\dc_ew[57][4] ,
    \dc_ew[57][3] ,
    \dc_ew[57][2] ,
    \dc_ew[57][1] ,
    \dc_ew[57][0] }),
    .cb_east_out({\dc_we[57][9] ,
    \dc_we[57][8] ,
    \dc_we[57][7] ,
    \dc_we[57][6] ,
    \dc_we[57][5] ,
    \dc_we[57][4] ,
    \dc_we[57][3] ,
    \dc_we[57][2] ,
    \dc_we[57][1] ,
    \dc_we[57][0] }),
    .cb_north_in({_085_,
    _084_,
    _083_,
    _082_,
    _081_}),
    .cb_north_out({\dc_sn[56][9] ,
    \dc_sn[56][8] ,
    \dc_sn[56][7] ,
    \dc_sn[56][6] ,
    \dc_sn[56][5] ,
    \dc_sn[56][4] ,
    \dc_sn[56][3] ,
    \dc_sn[56][2] ,
    \dc_sn[56][1] ,
    \dc_sn[56][0] }),
    .clb_south_in({\dc_sn[49][9] ,
    \dc_sn[49][8] ,
    \dc_sn[49][7] ,
    \dc_sn[49][6] ,
    \dc_sn[49][5] ,
    \dc_sn[49][4] ,
    \dc_sn[49][3] ,
    \dc_sn[49][2] ,
    \dc_sn[49][1] ,
    \dc_sn[49][0] }),
    .clb_south_out({\dc_ns[49][4] ,
    \dc_ns[49][3] ,
    \dc_ns[49][2] ,
    \dc_ns[49][1] ,
    \dc_ns[49][0] }),
    .clb_west_in({_095_,
    _094_,
    _093_,
    _092_,
    _091_,
    _090_,
    _089_,
    _088_,
    _087_,
    _086_}),
    .clb_west_out({\dc_ew[56][4] ,
    \dc_ew[56][3] ,
    \dc_ew[56][2] ,
    \dc_ew[56][1] ,
    \dc_ew[56][0] }),
    .east_double({\ix_double_ew[57][7] ,
    \ix_double_ew[57][6] ,
    \ix_double_ew[57][5] ,
    \ix_double_ew[57][4] ,
    \ix_double_ew[57][3] ,
    \ix_double_ew[57][2] ,
    \ix_double_ew[57][1] ,
    \ix_double_ew[57][0] }),
    .east_single({\ix_single_ew[57][3] ,
    \ix_single_ew[57][2] ,
    \ix_single_ew[57][1] ,
    \ix_single_ew[57][0] }),
    .north_double({\ix_double_ns[56][7] ,
    \ix_double_ns[56][6] ,
    \ix_double_ns[56][5] ,
    \ix_double_ns[56][4] ,
    \ix_double_ns[56][3] ,
    \ix_double_ns[56][2] ,
    \ix_double_ns[56][1] ,
    \ix_double_ns[56][0] }),
    .north_single({\ix_single_ns[56][3] ,
    \ix_single_ns[56][2] ,
    \ix_single_ns[56][1] ,
    gpio_north[0]}),
    .south_double({\ix_double_ns[49][7] ,
    \ix_double_ns[49][6] ,
    \ix_double_ns[49][5] ,
    \ix_double_ns[49][4] ,
    \ix_double_ns[49][3] ,
    \ix_double_ns[49][2] ,
    \ix_double_ns[49][1] ,
    \ix_double_ns[49][0] }),
    .south_single({\ix_single_ns[49][3] ,
    \ix_single_ns[49][2] ,
    \ix_single_ns[49][1] ,
    \ix_single_ns[49][0] }),
    .west_double({\ix_double_ew[56][7] ,
    \ix_double_ew[56][6] ,
    \ix_double_ew[56][5] ,
    \ix_double_ew[56][4] ,
    \ix_double_ew[56][3] ,
    \ix_double_ew[56][2] ,
    \ix_double_ew[56][1] ,
    \ix_double_ew[56][0] }),
    .west_single({\ix_single_ew[56][3] ,
    \ix_single_ew[56][2] ,
    \ix_single_ew[56][1] ,
    gpio_west[7]}));
 clb_tile \X[1].Y[0].clb  (.carry_in(_096_),
    .carry_out(\carry[1][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[0][1] ),
    .set_out_hard(\col_set[1][1] ),
    .shift_in_hard(\wb_shift_out[0][1] ),
    .shift_out_hard(\col_shift[1][1] ),
    .cb_east_in({\dc_ew[2][4] ,
    \dc_ew[2][3] ,
    \dc_ew[2][2] ,
    \dc_ew[2][1] ,
    \dc_ew[2][0] }),
    .cb_east_out({\dc_we[2][9] ,
    \dc_we[2][8] ,
    \dc_we[2][7] ,
    \dc_we[2][6] ,
    \dc_we[2][5] ,
    \dc_we[2][4] ,
    \dc_we[2][3] ,
    \dc_we[2][2] ,
    \dc_we[2][1] ,
    \dc_we[2][0] }),
    .cb_north_in({\dc_ns[8][4] ,
    \dc_ns[8][3] ,
    \dc_ns[8][2] ,
    \dc_ns[8][1] ,
    \dc_ns[8][0] }),
    .cb_north_out({\dc_sn[8][9] ,
    \dc_sn[8][8] ,
    \dc_sn[8][7] ,
    \dc_sn[8][6] ,
    \dc_sn[8][5] ,
    \dc_sn[8][4] ,
    \dc_sn[8][3] ,
    \dc_sn[8][2] ,
    \dc_sn[8][1] ,
    \dc_sn[8][0] }),
    .clb_south_in({_106_,
    _105_,
    _104_,
    _103_,
    _102_,
    _101_,
    _100_,
    _099_,
    _098_,
    _097_}),
    .clb_south_out({\dc_ns[1][4] ,
    \dc_ns[1][3] ,
    \dc_ns[1][2] ,
    \dc_ns[1][1] ,
    \dc_ns[1][0] }),
    .clb_west_in({\dc_we[1][9] ,
    \dc_we[1][8] ,
    \dc_we[1][7] ,
    \dc_we[1][6] ,
    \dc_we[1][5] ,
    \dc_we[1][4] ,
    \dc_we[1][3] ,
    \dc_we[1][2] ,
    \dc_we[1][1] ,
    \dc_we[1][0] }),
    .clb_west_out({\dc_ew[1][4] ,
    \dc_ew[1][3] ,
    \dc_ew[1][2] ,
    \dc_ew[1][1] ,
    \dc_ew[1][0] }),
    .east_double({\ix_double_ew[2][7] ,
    \ix_double_ew[2][6] ,
    \ix_double_ew[2][5] ,
    \ix_double_ew[2][4] ,
    \ix_double_ew[2][3] ,
    \ix_double_ew[2][2] ,
    \ix_double_ew[2][1] ,
    \ix_double_ew[2][0] }),
    .east_single({\ix_single_ew[2][3] ,
    \ix_single_ew[2][2] ,
    \ix_single_ew[2][1] ,
    \ix_single_ew[2][0] }),
    .north_double({\ix_double_ns[8][7] ,
    \ix_double_ns[8][6] ,
    \ix_double_ns[8][5] ,
    \ix_double_ns[8][4] ,
    \ix_double_ns[8][3] ,
    \ix_double_ns[8][2] ,
    \ix_double_ns[8][1] ,
    \ix_double_ns[8][0] }),
    .north_single({\ix_single_ns[8][3] ,
    \ix_single_ns[8][2] ,
    \ix_single_ns[8][1] ,
    \ix_single_ns[8][0] }),
    .south_double({\ix_double_ns[1][7] ,
    \ix_double_ns[1][6] ,
    \ix_double_ns[1][5] ,
    \ix_double_ns[1][4] ,
    \ix_double_ns[1][3] ,
    \ix_double_ns[1][2] ,
    \ix_double_ns[1][1] ,
    \ix_double_ns[1][0] }),
    .south_single({\ix_single_ns[1][3] ,
    \ix_single_ns[1][2] ,
    \ix_single_ns[1][1] ,
    gpio_south[1]}),
    .west_double({\ix_double_ew[1][7] ,
    \ix_double_ew[1][6] ,
    \ix_double_ew[1][5] ,
    \ix_double_ew[1][4] ,
    \ix_double_ew[1][3] ,
    \ix_double_ew[1][2] ,
    \ix_double_ew[1][1] ,
    \ix_double_ew[1][0] }),
    .west_single({\ix_single_ew[1][3] ,
    \ix_single_ew[1][2] ,
    \ix_single_ew[1][1] ,
    \ix_single_ew[1][0] }));
 clb_tile \X[1].Y[1].clb  (.carry_in(\carry[1][1] ),
    .carry_out(\carry[2][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][1] ),
    .set_out_hard(\col_set[2][1] ),
    .shift_in_hard(\col_shift[1][1] ),
    .shift_out_hard(\col_shift[2][1] ),
    .cb_east_in({\dc_ew[10][4] ,
    \dc_ew[10][3] ,
    \dc_ew[10][2] ,
    \dc_ew[10][1] ,
    \dc_ew[10][0] }),
    .cb_east_out({\dc_we[10][9] ,
    \dc_we[10][8] ,
    \dc_we[10][7] ,
    \dc_we[10][6] ,
    \dc_we[10][5] ,
    \dc_we[10][4] ,
    \dc_we[10][3] ,
    \dc_we[10][2] ,
    \dc_we[10][1] ,
    \dc_we[10][0] }),
    .cb_north_in({\dc_ns[15][4] ,
    \dc_ns[15][3] ,
    \dc_ns[15][2] ,
    \dc_ns[15][1] ,
    \dc_ns[15][0] }),
    .cb_north_out({\dc_sn[15][9] ,
    \dc_sn[15][8] ,
    \dc_sn[15][7] ,
    \dc_sn[15][6] ,
    \dc_sn[15][5] ,
    \dc_sn[15][4] ,
    \dc_sn[15][3] ,
    \dc_sn[15][2] ,
    \dc_sn[15][1] ,
    \dc_sn[15][0] }),
    .clb_south_in({\dc_sn[8][9] ,
    \dc_sn[8][8] ,
    \dc_sn[8][7] ,
    \dc_sn[8][6] ,
    \dc_sn[8][5] ,
    \dc_sn[8][4] ,
    \dc_sn[8][3] ,
    \dc_sn[8][2] ,
    \dc_sn[8][1] ,
    \dc_sn[8][0] }),
    .clb_south_out({\dc_ns[8][4] ,
    \dc_ns[8][3] ,
    \dc_ns[8][2] ,
    \dc_ns[8][1] ,
    \dc_ns[8][0] }),
    .clb_west_in({\dc_we[9][9] ,
    \dc_we[9][8] ,
    \dc_we[9][7] ,
    \dc_we[9][6] ,
    \dc_we[9][5] ,
    \dc_we[9][4] ,
    \dc_we[9][3] ,
    \dc_we[9][2] ,
    \dc_we[9][1] ,
    \dc_we[9][0] }),
    .clb_west_out({\dc_ew[9][4] ,
    \dc_ew[9][3] ,
    \dc_ew[9][2] ,
    \dc_ew[9][1] ,
    \dc_ew[9][0] }),
    .east_double({\ix_double_ew[10][7] ,
    \ix_double_ew[10][6] ,
    \ix_double_ew[10][5] ,
    \ix_double_ew[10][4] ,
    \ix_double_ew[10][3] ,
    \ix_double_ew[10][2] ,
    \ix_double_ew[10][1] ,
    \ix_double_ew[10][0] }),
    .east_single({\ix_single_ew[10][3] ,
    \ix_single_ew[10][2] ,
    \ix_single_ew[10][1] ,
    \ix_single_ew[10][0] }),
    .north_double({\ix_double_ns[15][7] ,
    \ix_double_ns[15][6] ,
    \ix_double_ns[15][5] ,
    \ix_double_ns[15][4] ,
    \ix_double_ns[15][3] ,
    \ix_double_ns[15][2] ,
    \ix_double_ns[15][1] ,
    \ix_double_ns[15][0] }),
    .north_single({\ix_single_ns[15][3] ,
    \ix_single_ns[15][2] ,
    \ix_single_ns[15][1] ,
    \ix_single_ns[15][0] }),
    .south_double({\ix_double_ns[8][7] ,
    \ix_double_ns[8][6] ,
    \ix_double_ns[8][5] ,
    \ix_double_ns[8][4] ,
    \ix_double_ns[8][3] ,
    \ix_double_ns[8][2] ,
    \ix_double_ns[8][1] ,
    \ix_double_ns[8][0] }),
    .south_single({\ix_single_ns[8][3] ,
    \ix_single_ns[8][2] ,
    \ix_single_ns[8][1] ,
    \ix_single_ns[8][0] }),
    .west_double({\ix_double_ew[9][7] ,
    \ix_double_ew[9][6] ,
    \ix_double_ew[9][5] ,
    \ix_double_ew[9][4] ,
    \ix_double_ew[9][3] ,
    \ix_double_ew[9][2] ,
    \ix_double_ew[9][1] ,
    \ix_double_ew[9][0] }),
    .west_single({\ix_single_ew[9][3] ,
    \ix_single_ew[9][2] ,
    \ix_single_ew[9][1] ,
    \ix_single_ew[9][0] }));
 clb_tile \X[1].Y[2].clb  (.carry_in(\carry[2][1] ),
    .carry_out(\carry[3][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][1] ),
    .set_out_hard(\col_set[3][1] ),
    .shift_in_hard(\col_shift[2][1] ),
    .shift_out_hard(\col_shift[3][1] ),
    .cb_east_in({\dc_ew[18][4] ,
    \dc_ew[18][3] ,
    \dc_ew[18][2] ,
    \dc_ew[18][1] ,
    \dc_ew[18][0] }),
    .cb_east_out({\dc_we[18][9] ,
    \dc_we[18][8] ,
    \dc_we[18][7] ,
    \dc_we[18][6] ,
    \dc_we[18][5] ,
    \dc_we[18][4] ,
    \dc_we[18][3] ,
    \dc_we[18][2] ,
    \dc_we[18][1] ,
    \dc_we[18][0] }),
    .cb_north_in({\dc_ns[22][4] ,
    \dc_ns[22][3] ,
    \dc_ns[22][2] ,
    \dc_ns[22][1] ,
    \dc_ns[22][0] }),
    .cb_north_out({\dc_sn[22][9] ,
    \dc_sn[22][8] ,
    \dc_sn[22][7] ,
    \dc_sn[22][6] ,
    \dc_sn[22][5] ,
    \dc_sn[22][4] ,
    \dc_sn[22][3] ,
    \dc_sn[22][2] ,
    \dc_sn[22][1] ,
    \dc_sn[22][0] }),
    .clb_south_in({\dc_sn[15][9] ,
    \dc_sn[15][8] ,
    \dc_sn[15][7] ,
    \dc_sn[15][6] ,
    \dc_sn[15][5] ,
    \dc_sn[15][4] ,
    \dc_sn[15][3] ,
    \dc_sn[15][2] ,
    \dc_sn[15][1] ,
    \dc_sn[15][0] }),
    .clb_south_out({\dc_ns[15][4] ,
    \dc_ns[15][3] ,
    \dc_ns[15][2] ,
    \dc_ns[15][1] ,
    \dc_ns[15][0] }),
    .clb_west_in({\dc_we[17][9] ,
    \dc_we[17][8] ,
    \dc_we[17][7] ,
    \dc_we[17][6] ,
    \dc_we[17][5] ,
    \dc_we[17][4] ,
    \dc_we[17][3] ,
    \dc_we[17][2] ,
    \dc_we[17][1] ,
    \dc_we[17][0] }),
    .clb_west_out({\dc_ew[17][4] ,
    \dc_ew[17][3] ,
    \dc_ew[17][2] ,
    \dc_ew[17][1] ,
    \dc_ew[17][0] }),
    .east_double({\ix_double_ew[18][7] ,
    \ix_double_ew[18][6] ,
    \ix_double_ew[18][5] ,
    \ix_double_ew[18][4] ,
    \ix_double_ew[18][3] ,
    \ix_double_ew[18][2] ,
    \ix_double_ew[18][1] ,
    \ix_double_ew[18][0] }),
    .east_single({\ix_single_ew[18][3] ,
    \ix_single_ew[18][2] ,
    \ix_single_ew[18][1] ,
    \ix_single_ew[18][0] }),
    .north_double({\ix_double_ns[22][7] ,
    \ix_double_ns[22][6] ,
    \ix_double_ns[22][5] ,
    \ix_double_ns[22][4] ,
    \ix_double_ns[22][3] ,
    \ix_double_ns[22][2] ,
    \ix_double_ns[22][1] ,
    \ix_double_ns[22][0] }),
    .north_single({\ix_single_ns[22][3] ,
    \ix_single_ns[22][2] ,
    \ix_single_ns[22][1] ,
    \ix_single_ns[22][0] }),
    .south_double({\ix_double_ns[15][7] ,
    \ix_double_ns[15][6] ,
    \ix_double_ns[15][5] ,
    \ix_double_ns[15][4] ,
    \ix_double_ns[15][3] ,
    \ix_double_ns[15][2] ,
    \ix_double_ns[15][1] ,
    \ix_double_ns[15][0] }),
    .south_single({\ix_single_ns[15][3] ,
    \ix_single_ns[15][2] ,
    \ix_single_ns[15][1] ,
    \ix_single_ns[15][0] }),
    .west_double({\ix_double_ew[17][7] ,
    \ix_double_ew[17][6] ,
    \ix_double_ew[17][5] ,
    \ix_double_ew[17][4] ,
    \ix_double_ew[17][3] ,
    \ix_double_ew[17][2] ,
    \ix_double_ew[17][1] ,
    \ix_double_ew[17][0] }),
    .west_single({\ix_single_ew[17][3] ,
    \ix_single_ew[17][2] ,
    \ix_single_ew[17][1] ,
    \ix_single_ew[17][0] }));
 clb_tile \X[1].Y[3].clb  (.carry_in(\carry[3][1] ),
    .carry_out(\carry[4][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][1] ),
    .set_out_hard(\col_set[4][1] ),
    .shift_in_hard(\col_shift[3][1] ),
    .shift_out_hard(\col_shift[4][1] ),
    .cb_east_in({\dc_ew[26][4] ,
    \dc_ew[26][3] ,
    \dc_ew[26][2] ,
    \dc_ew[26][1] ,
    \dc_ew[26][0] }),
    .cb_east_out({\dc_we[26][9] ,
    \dc_we[26][8] ,
    \dc_we[26][7] ,
    \dc_we[26][6] ,
    \dc_we[26][5] ,
    \dc_we[26][4] ,
    \dc_we[26][3] ,
    \dc_we[26][2] ,
    \dc_we[26][1] ,
    \dc_we[26][0] }),
    .cb_north_in({\dc_ns[29][4] ,
    \dc_ns[29][3] ,
    \dc_ns[29][2] ,
    \dc_ns[29][1] ,
    \dc_ns[29][0] }),
    .cb_north_out({\dc_sn[29][9] ,
    \dc_sn[29][8] ,
    \dc_sn[29][7] ,
    \dc_sn[29][6] ,
    \dc_sn[29][5] ,
    \dc_sn[29][4] ,
    \dc_sn[29][3] ,
    \dc_sn[29][2] ,
    \dc_sn[29][1] ,
    \dc_sn[29][0] }),
    .clb_south_in({\dc_sn[22][9] ,
    \dc_sn[22][8] ,
    \dc_sn[22][7] ,
    \dc_sn[22][6] ,
    \dc_sn[22][5] ,
    \dc_sn[22][4] ,
    \dc_sn[22][3] ,
    \dc_sn[22][2] ,
    \dc_sn[22][1] ,
    \dc_sn[22][0] }),
    .clb_south_out({\dc_ns[22][4] ,
    \dc_ns[22][3] ,
    \dc_ns[22][2] ,
    \dc_ns[22][1] ,
    \dc_ns[22][0] }),
    .clb_west_in({\dc_we[25][9] ,
    \dc_we[25][8] ,
    \dc_we[25][7] ,
    \dc_we[25][6] ,
    \dc_we[25][5] ,
    \dc_we[25][4] ,
    \dc_we[25][3] ,
    \dc_we[25][2] ,
    \dc_we[25][1] ,
    \dc_we[25][0] }),
    .clb_west_out({\dc_ew[25][4] ,
    \dc_ew[25][3] ,
    \dc_ew[25][2] ,
    \dc_ew[25][1] ,
    \dc_ew[25][0] }),
    .east_double({\ix_double_ew[26][7] ,
    \ix_double_ew[26][6] ,
    \ix_double_ew[26][5] ,
    \ix_double_ew[26][4] ,
    \ix_double_ew[26][3] ,
    \ix_double_ew[26][2] ,
    \ix_double_ew[26][1] ,
    \ix_double_ew[26][0] }),
    .east_single({\ix_single_ew[26][3] ,
    \ix_single_ew[26][2] ,
    \ix_single_ew[26][1] ,
    \ix_single_ew[26][0] }),
    .north_double({\ix_double_ns[29][7] ,
    \ix_double_ns[29][6] ,
    \ix_double_ns[29][5] ,
    \ix_double_ns[29][4] ,
    \ix_double_ns[29][3] ,
    \ix_double_ns[29][2] ,
    \ix_double_ns[29][1] ,
    \ix_double_ns[29][0] }),
    .north_single({\ix_single_ns[29][3] ,
    \ix_single_ns[29][2] ,
    \ix_single_ns[29][1] ,
    \ix_single_ns[29][0] }),
    .south_double({\ix_double_ns[22][7] ,
    \ix_double_ns[22][6] ,
    \ix_double_ns[22][5] ,
    \ix_double_ns[22][4] ,
    \ix_double_ns[22][3] ,
    \ix_double_ns[22][2] ,
    \ix_double_ns[22][1] ,
    \ix_double_ns[22][0] }),
    .south_single({\ix_single_ns[22][3] ,
    \ix_single_ns[22][2] ,
    \ix_single_ns[22][1] ,
    \ix_single_ns[22][0] }),
    .west_double({\ix_double_ew[25][7] ,
    \ix_double_ew[25][6] ,
    \ix_double_ew[25][5] ,
    \ix_double_ew[25][4] ,
    \ix_double_ew[25][3] ,
    \ix_double_ew[25][2] ,
    \ix_double_ew[25][1] ,
    \ix_double_ew[25][0] }),
    .west_single({\ix_single_ew[25][3] ,
    \ix_single_ew[25][2] ,
    \ix_single_ew[25][1] ,
    \ix_single_ew[25][0] }));
 clb_tile \X[1].Y[4].clb  (.carry_in(\carry[4][1] ),
    .carry_out(\carry[5][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][1] ),
    .set_out_hard(\col_set[5][1] ),
    .shift_in_hard(\col_shift[4][1] ),
    .shift_out_hard(\col_shift[5][1] ),
    .cb_east_in({\dc_ew[34][4] ,
    \dc_ew[34][3] ,
    \dc_ew[34][2] ,
    \dc_ew[34][1] ,
    \dc_ew[34][0] }),
    .cb_east_out({\dc_we[34][9] ,
    \dc_we[34][8] ,
    \dc_we[34][7] ,
    \dc_we[34][6] ,
    \dc_we[34][5] ,
    \dc_we[34][4] ,
    \dc_we[34][3] ,
    \dc_we[34][2] ,
    \dc_we[34][1] ,
    \dc_we[34][0] }),
    .cb_north_in({\dc_ns[36][4] ,
    \dc_ns[36][3] ,
    \dc_ns[36][2] ,
    \dc_ns[36][1] ,
    \dc_ns[36][0] }),
    .cb_north_out({\dc_sn[36][9] ,
    \dc_sn[36][8] ,
    \dc_sn[36][7] ,
    \dc_sn[36][6] ,
    \dc_sn[36][5] ,
    \dc_sn[36][4] ,
    \dc_sn[36][3] ,
    \dc_sn[36][2] ,
    \dc_sn[36][1] ,
    \dc_sn[36][0] }),
    .clb_south_in({\dc_sn[29][9] ,
    \dc_sn[29][8] ,
    \dc_sn[29][7] ,
    \dc_sn[29][6] ,
    \dc_sn[29][5] ,
    \dc_sn[29][4] ,
    \dc_sn[29][3] ,
    \dc_sn[29][2] ,
    \dc_sn[29][1] ,
    \dc_sn[29][0] }),
    .clb_south_out({\dc_ns[29][4] ,
    \dc_ns[29][3] ,
    \dc_ns[29][2] ,
    \dc_ns[29][1] ,
    \dc_ns[29][0] }),
    .clb_west_in({\dc_we[33][9] ,
    \dc_we[33][8] ,
    \dc_we[33][7] ,
    \dc_we[33][6] ,
    \dc_we[33][5] ,
    \dc_we[33][4] ,
    \dc_we[33][3] ,
    \dc_we[33][2] ,
    \dc_we[33][1] ,
    \dc_we[33][0] }),
    .clb_west_out({\dc_ew[33][4] ,
    \dc_ew[33][3] ,
    \dc_ew[33][2] ,
    \dc_ew[33][1] ,
    \dc_ew[33][0] }),
    .east_double({\ix_double_ew[34][7] ,
    \ix_double_ew[34][6] ,
    \ix_double_ew[34][5] ,
    \ix_double_ew[34][4] ,
    \ix_double_ew[34][3] ,
    \ix_double_ew[34][2] ,
    \ix_double_ew[34][1] ,
    \ix_double_ew[34][0] }),
    .east_single({\ix_single_ew[34][3] ,
    \ix_single_ew[34][2] ,
    \ix_single_ew[34][1] ,
    \ix_single_ew[34][0] }),
    .north_double({\ix_double_ns[36][7] ,
    \ix_double_ns[36][6] ,
    \ix_double_ns[36][5] ,
    \ix_double_ns[36][4] ,
    \ix_double_ns[36][3] ,
    \ix_double_ns[36][2] ,
    \ix_double_ns[36][1] ,
    \ix_double_ns[36][0] }),
    .north_single({\ix_single_ns[36][3] ,
    \ix_single_ns[36][2] ,
    \ix_single_ns[36][1] ,
    \ix_single_ns[36][0] }),
    .south_double({\ix_double_ns[29][7] ,
    \ix_double_ns[29][6] ,
    \ix_double_ns[29][5] ,
    \ix_double_ns[29][4] ,
    \ix_double_ns[29][3] ,
    \ix_double_ns[29][2] ,
    \ix_double_ns[29][1] ,
    \ix_double_ns[29][0] }),
    .south_single({\ix_single_ns[29][3] ,
    \ix_single_ns[29][2] ,
    \ix_single_ns[29][1] ,
    \ix_single_ns[29][0] }),
    .west_double({\ix_double_ew[33][7] ,
    \ix_double_ew[33][6] ,
    \ix_double_ew[33][5] ,
    \ix_double_ew[33][4] ,
    \ix_double_ew[33][3] ,
    \ix_double_ew[33][2] ,
    \ix_double_ew[33][1] ,
    \ix_double_ew[33][0] }),
    .west_single({\ix_single_ew[33][3] ,
    \ix_single_ew[33][2] ,
    \ix_single_ew[33][1] ,
    \ix_single_ew[33][0] }));
 clb_tile \X[1].Y[5].clb  (.carry_in(\carry[5][1] ),
    .carry_out(\carry[6][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][1] ),
    .set_out_hard(\col_set[6][1] ),
    .shift_in_hard(\col_shift[5][1] ),
    .shift_out_hard(\col_shift[6][1] ),
    .cb_east_in({\dc_ew[42][4] ,
    \dc_ew[42][3] ,
    \dc_ew[42][2] ,
    \dc_ew[42][1] ,
    \dc_ew[42][0] }),
    .cb_east_out({\dc_we[42][9] ,
    \dc_we[42][8] ,
    \dc_we[42][7] ,
    \dc_we[42][6] ,
    \dc_we[42][5] ,
    \dc_we[42][4] ,
    \dc_we[42][3] ,
    \dc_we[42][2] ,
    \dc_we[42][1] ,
    \dc_we[42][0] }),
    .cb_north_in({\dc_ns[43][4] ,
    \dc_ns[43][3] ,
    \dc_ns[43][2] ,
    \dc_ns[43][1] ,
    \dc_ns[43][0] }),
    .cb_north_out({\dc_sn[43][9] ,
    \dc_sn[43][8] ,
    \dc_sn[43][7] ,
    \dc_sn[43][6] ,
    \dc_sn[43][5] ,
    \dc_sn[43][4] ,
    \dc_sn[43][3] ,
    \dc_sn[43][2] ,
    \dc_sn[43][1] ,
    \dc_sn[43][0] }),
    .clb_south_in({\dc_sn[36][9] ,
    \dc_sn[36][8] ,
    \dc_sn[36][7] ,
    \dc_sn[36][6] ,
    \dc_sn[36][5] ,
    \dc_sn[36][4] ,
    \dc_sn[36][3] ,
    \dc_sn[36][2] ,
    \dc_sn[36][1] ,
    \dc_sn[36][0] }),
    .clb_south_out({\dc_ns[36][4] ,
    \dc_ns[36][3] ,
    \dc_ns[36][2] ,
    \dc_ns[36][1] ,
    \dc_ns[36][0] }),
    .clb_west_in({\dc_we[41][9] ,
    \dc_we[41][8] ,
    \dc_we[41][7] ,
    \dc_we[41][6] ,
    \dc_we[41][5] ,
    \dc_we[41][4] ,
    \dc_we[41][3] ,
    \dc_we[41][2] ,
    \dc_we[41][1] ,
    \dc_we[41][0] }),
    .clb_west_out({\dc_ew[41][4] ,
    \dc_ew[41][3] ,
    \dc_ew[41][2] ,
    \dc_ew[41][1] ,
    \dc_ew[41][0] }),
    .east_double({\ix_double_ew[42][7] ,
    \ix_double_ew[42][6] ,
    \ix_double_ew[42][5] ,
    \ix_double_ew[42][4] ,
    \ix_double_ew[42][3] ,
    \ix_double_ew[42][2] ,
    \ix_double_ew[42][1] ,
    \ix_double_ew[42][0] }),
    .east_single({\ix_single_ew[42][3] ,
    \ix_single_ew[42][2] ,
    \ix_single_ew[42][1] ,
    \ix_single_ew[42][0] }),
    .north_double({\ix_double_ns[43][7] ,
    \ix_double_ns[43][6] ,
    \ix_double_ns[43][5] ,
    \ix_double_ns[43][4] ,
    \ix_double_ns[43][3] ,
    \ix_double_ns[43][2] ,
    \ix_double_ns[43][1] ,
    \ix_double_ns[43][0] }),
    .north_single({\ix_single_ns[43][3] ,
    \ix_single_ns[43][2] ,
    \ix_single_ns[43][1] ,
    \ix_single_ns[43][0] }),
    .south_double({\ix_double_ns[36][7] ,
    \ix_double_ns[36][6] ,
    \ix_double_ns[36][5] ,
    \ix_double_ns[36][4] ,
    \ix_double_ns[36][3] ,
    \ix_double_ns[36][2] ,
    \ix_double_ns[36][1] ,
    \ix_double_ns[36][0] }),
    .south_single({\ix_single_ns[36][3] ,
    \ix_single_ns[36][2] ,
    \ix_single_ns[36][1] ,
    \ix_single_ns[36][0] }),
    .west_double({\ix_double_ew[41][7] ,
    \ix_double_ew[41][6] ,
    \ix_double_ew[41][5] ,
    \ix_double_ew[41][4] ,
    \ix_double_ew[41][3] ,
    \ix_double_ew[41][2] ,
    \ix_double_ew[41][1] ,
    \ix_double_ew[41][0] }),
    .west_single({\ix_single_ew[41][3] ,
    \ix_single_ew[41][2] ,
    \ix_single_ew[41][1] ,
    \ix_single_ew[41][0] }));
 clb_tile \X[1].Y[6].clb  (.carry_in(\carry[6][1] ),
    .carry_out(\carry[7][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][1] ),
    .set_out_hard(\col_set[7][1] ),
    .shift_in_hard(\col_shift[6][1] ),
    .shift_out_hard(\col_shift[7][1] ),
    .cb_east_in({\dc_ew[50][4] ,
    \dc_ew[50][3] ,
    \dc_ew[50][2] ,
    \dc_ew[50][1] ,
    \dc_ew[50][0] }),
    .cb_east_out({\dc_we[50][9] ,
    \dc_we[50][8] ,
    \dc_we[50][7] ,
    \dc_we[50][6] ,
    \dc_we[50][5] ,
    \dc_we[50][4] ,
    \dc_we[50][3] ,
    \dc_we[50][2] ,
    \dc_we[50][1] ,
    \dc_we[50][0] }),
    .cb_north_in({\dc_ns[50][4] ,
    \dc_ns[50][3] ,
    \dc_ns[50][2] ,
    \dc_ns[50][1] ,
    \dc_ns[50][0] }),
    .cb_north_out({\dc_sn[50][9] ,
    \dc_sn[50][8] ,
    \dc_sn[50][7] ,
    \dc_sn[50][6] ,
    \dc_sn[50][5] ,
    \dc_sn[50][4] ,
    \dc_sn[50][3] ,
    \dc_sn[50][2] ,
    \dc_sn[50][1] ,
    \dc_sn[50][0] }),
    .clb_south_in({\dc_sn[43][9] ,
    \dc_sn[43][8] ,
    \dc_sn[43][7] ,
    \dc_sn[43][6] ,
    \dc_sn[43][5] ,
    \dc_sn[43][4] ,
    \dc_sn[43][3] ,
    \dc_sn[43][2] ,
    \dc_sn[43][1] ,
    \dc_sn[43][0] }),
    .clb_south_out({\dc_ns[43][4] ,
    \dc_ns[43][3] ,
    \dc_ns[43][2] ,
    \dc_ns[43][1] ,
    \dc_ns[43][0] }),
    .clb_west_in({\dc_we[49][9] ,
    \dc_we[49][8] ,
    \dc_we[49][7] ,
    \dc_we[49][6] ,
    \dc_we[49][5] ,
    \dc_we[49][4] ,
    \dc_we[49][3] ,
    \dc_we[49][2] ,
    \dc_we[49][1] ,
    \dc_we[49][0] }),
    .clb_west_out({\dc_ew[49][4] ,
    \dc_ew[49][3] ,
    \dc_ew[49][2] ,
    \dc_ew[49][1] ,
    \dc_ew[49][0] }),
    .east_double({\ix_double_ew[50][7] ,
    \ix_double_ew[50][6] ,
    \ix_double_ew[50][5] ,
    \ix_double_ew[50][4] ,
    \ix_double_ew[50][3] ,
    \ix_double_ew[50][2] ,
    \ix_double_ew[50][1] ,
    \ix_double_ew[50][0] }),
    .east_single({\ix_single_ew[50][3] ,
    \ix_single_ew[50][2] ,
    \ix_single_ew[50][1] ,
    \ix_single_ew[50][0] }),
    .north_double({\ix_double_ns[50][7] ,
    \ix_double_ns[50][6] ,
    \ix_double_ns[50][5] ,
    \ix_double_ns[50][4] ,
    \ix_double_ns[50][3] ,
    \ix_double_ns[50][2] ,
    \ix_double_ns[50][1] ,
    \ix_double_ns[50][0] }),
    .north_single({\ix_single_ns[50][3] ,
    \ix_single_ns[50][2] ,
    \ix_single_ns[50][1] ,
    \ix_single_ns[50][0] }),
    .south_double({\ix_double_ns[43][7] ,
    \ix_double_ns[43][6] ,
    \ix_double_ns[43][5] ,
    \ix_double_ns[43][4] ,
    \ix_double_ns[43][3] ,
    \ix_double_ns[43][2] ,
    \ix_double_ns[43][1] ,
    \ix_double_ns[43][0] }),
    .south_single({\ix_single_ns[43][3] ,
    \ix_single_ns[43][2] ,
    \ix_single_ns[43][1] ,
    \ix_single_ns[43][0] }),
    .west_double({\ix_double_ew[49][7] ,
    \ix_double_ew[49][6] ,
    \ix_double_ew[49][5] ,
    \ix_double_ew[49][4] ,
    \ix_double_ew[49][3] ,
    \ix_double_ew[49][2] ,
    \ix_double_ew[49][1] ,
    \ix_double_ew[49][0] }),
    .west_single({\ix_single_ew[49][3] ,
    \ix_single_ew[49][2] ,
    \ix_single_ew[49][1] ,
    \ix_single_ew[49][0] }));
 clb_tile \X[1].Y[7].clb  (.carry_in(\carry[7][1] ),
    .carry_out(\carry[8][1] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][1] ),
    .set_out_hard(\col_set[8][1] ),
    .shift_in_hard(\col_shift[7][1] ),
    .shift_out_hard(\col_shift[8][1] ),
    .cb_east_in({\dc_ew[58][4] ,
    \dc_ew[58][3] ,
    \dc_ew[58][2] ,
    \dc_ew[58][1] ,
    \dc_ew[58][0] }),
    .cb_east_out({\dc_we[58][9] ,
    \dc_we[58][8] ,
    \dc_we[58][7] ,
    \dc_we[58][6] ,
    \dc_we[58][5] ,
    \dc_we[58][4] ,
    \dc_we[58][3] ,
    \dc_we[58][2] ,
    \dc_we[58][1] ,
    \dc_we[58][0] }),
    .cb_north_in({_111_,
    _110_,
    _109_,
    _108_,
    _107_}),
    .cb_north_out({\dc_sn[57][9] ,
    \dc_sn[57][8] ,
    \dc_sn[57][7] ,
    \dc_sn[57][6] ,
    \dc_sn[57][5] ,
    \dc_sn[57][4] ,
    \dc_sn[57][3] ,
    \dc_sn[57][2] ,
    \dc_sn[57][1] ,
    \dc_sn[57][0] }),
    .clb_south_in({\dc_sn[50][9] ,
    \dc_sn[50][8] ,
    \dc_sn[50][7] ,
    \dc_sn[50][6] ,
    \dc_sn[50][5] ,
    \dc_sn[50][4] ,
    \dc_sn[50][3] ,
    \dc_sn[50][2] ,
    \dc_sn[50][1] ,
    \dc_sn[50][0] }),
    .clb_south_out({\dc_ns[50][4] ,
    \dc_ns[50][3] ,
    \dc_ns[50][2] ,
    \dc_ns[50][1] ,
    \dc_ns[50][0] }),
    .clb_west_in({\dc_we[57][9] ,
    \dc_we[57][8] ,
    \dc_we[57][7] ,
    \dc_we[57][6] ,
    \dc_we[57][5] ,
    \dc_we[57][4] ,
    \dc_we[57][3] ,
    \dc_we[57][2] ,
    \dc_we[57][1] ,
    \dc_we[57][0] }),
    .clb_west_out({\dc_ew[57][4] ,
    \dc_ew[57][3] ,
    \dc_ew[57][2] ,
    \dc_ew[57][1] ,
    \dc_ew[57][0] }),
    .east_double({\ix_double_ew[58][7] ,
    \ix_double_ew[58][6] ,
    \ix_double_ew[58][5] ,
    \ix_double_ew[58][4] ,
    \ix_double_ew[58][3] ,
    \ix_double_ew[58][2] ,
    \ix_double_ew[58][1] ,
    \ix_double_ew[58][0] }),
    .east_single({\ix_single_ew[58][3] ,
    \ix_single_ew[58][2] ,
    \ix_single_ew[58][1] ,
    \ix_single_ew[58][0] }),
    .north_double({\ix_double_ns[57][7] ,
    \ix_double_ns[57][6] ,
    \ix_double_ns[57][5] ,
    \ix_double_ns[57][4] ,
    \ix_double_ns[57][3] ,
    \ix_double_ns[57][2] ,
    \ix_double_ns[57][1] ,
    \ix_double_ns[57][0] }),
    .north_single({\ix_single_ns[57][3] ,
    \ix_single_ns[57][2] ,
    \ix_single_ns[57][1] ,
    gpio_north[1]}),
    .south_double({\ix_double_ns[50][7] ,
    \ix_double_ns[50][6] ,
    \ix_double_ns[50][5] ,
    \ix_double_ns[50][4] ,
    \ix_double_ns[50][3] ,
    \ix_double_ns[50][2] ,
    \ix_double_ns[50][1] ,
    \ix_double_ns[50][0] }),
    .south_single({\ix_single_ns[50][3] ,
    \ix_single_ns[50][2] ,
    \ix_single_ns[50][1] ,
    \ix_single_ns[50][0] }),
    .west_double({\ix_double_ew[57][7] ,
    \ix_double_ew[57][6] ,
    \ix_double_ew[57][5] ,
    \ix_double_ew[57][4] ,
    \ix_double_ew[57][3] ,
    \ix_double_ew[57][2] ,
    \ix_double_ew[57][1] ,
    \ix_double_ew[57][0] }),
    .west_single({\ix_single_ew[57][3] ,
    \ix_single_ew[57][2] ,
    \ix_single_ew[57][1] ,
    \ix_single_ew[57][0] }));
 clb_tile \X[2].Y[0].clb  (.carry_in(_112_),
    .carry_out(\carry[1][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[0][2] ),
    .set_out_hard(\col_set[1][2] ),
    .shift_in_hard(\wb_shift_out[0][2] ),
    .shift_out_hard(\col_shift[1][2] ),
    .cb_east_in({\dc_ew[3][4] ,
    \dc_ew[3][3] ,
    \dc_ew[3][2] ,
    \dc_ew[3][1] ,
    \dc_ew[3][0] }),
    .cb_east_out({\dc_we[3][9] ,
    \dc_we[3][8] ,
    \dc_we[3][7] ,
    \dc_we[3][6] ,
    \dc_we[3][5] ,
    \dc_we[3][4] ,
    \dc_we[3][3] ,
    \dc_we[3][2] ,
    \dc_we[3][1] ,
    \dc_we[3][0] }),
    .cb_north_in({\dc_ns[9][4] ,
    \dc_ns[9][3] ,
    \dc_ns[9][2] ,
    \dc_ns[9][1] ,
    \dc_ns[9][0] }),
    .cb_north_out({\dc_sn[9][9] ,
    \dc_sn[9][8] ,
    \dc_sn[9][7] ,
    \dc_sn[9][6] ,
    \dc_sn[9][5] ,
    \dc_sn[9][4] ,
    \dc_sn[9][3] ,
    \dc_sn[9][2] ,
    \dc_sn[9][1] ,
    \dc_sn[9][0] }),
    .clb_south_in({_122_,
    _121_,
    _120_,
    _119_,
    _118_,
    _117_,
    _116_,
    _115_,
    _114_,
    _113_}),
    .clb_south_out({\dc_ns[2][4] ,
    \dc_ns[2][3] ,
    \dc_ns[2][2] ,
    \dc_ns[2][1] ,
    \dc_ns[2][0] }),
    .clb_west_in({\dc_we[2][9] ,
    \dc_we[2][8] ,
    \dc_we[2][7] ,
    \dc_we[2][6] ,
    \dc_we[2][5] ,
    \dc_we[2][4] ,
    \dc_we[2][3] ,
    \dc_we[2][2] ,
    \dc_we[2][1] ,
    \dc_we[2][0] }),
    .clb_west_out({\dc_ew[2][4] ,
    \dc_ew[2][3] ,
    \dc_ew[2][2] ,
    \dc_ew[2][1] ,
    \dc_ew[2][0] }),
    .east_double({\ix_double_ew[3][7] ,
    \ix_double_ew[3][6] ,
    \ix_double_ew[3][5] ,
    \ix_double_ew[3][4] ,
    \ix_double_ew[3][3] ,
    \ix_double_ew[3][2] ,
    \ix_double_ew[3][1] ,
    \ix_double_ew[3][0] }),
    .east_single({\ix_single_ew[3][3] ,
    \ix_single_ew[3][2] ,
    \ix_single_ew[3][1] ,
    \ix_single_ew[3][0] }),
    .north_double({\ix_double_ns[9][7] ,
    \ix_double_ns[9][6] ,
    \ix_double_ns[9][5] ,
    \ix_double_ns[9][4] ,
    \ix_double_ns[9][3] ,
    \ix_double_ns[9][2] ,
    \ix_double_ns[9][1] ,
    \ix_double_ns[9][0] }),
    .north_single({\ix_single_ns[9][3] ,
    \ix_single_ns[9][2] ,
    \ix_single_ns[9][1] ,
    \ix_single_ns[9][0] }),
    .south_double({\ix_double_ns[2][7] ,
    \ix_double_ns[2][6] ,
    \ix_double_ns[2][5] ,
    \ix_double_ns[2][4] ,
    \ix_double_ns[2][3] ,
    \ix_double_ns[2][2] ,
    \ix_double_ns[2][1] ,
    \ix_double_ns[2][0] }),
    .south_single({\ix_single_ns[2][3] ,
    \ix_single_ns[2][2] ,
    \ix_single_ns[2][1] ,
    gpio_south[2]}),
    .west_double({\ix_double_ew[2][7] ,
    \ix_double_ew[2][6] ,
    \ix_double_ew[2][5] ,
    \ix_double_ew[2][4] ,
    \ix_double_ew[2][3] ,
    \ix_double_ew[2][2] ,
    \ix_double_ew[2][1] ,
    \ix_double_ew[2][0] }),
    .west_single({\ix_single_ew[2][3] ,
    \ix_single_ew[2][2] ,
    \ix_single_ew[2][1] ,
    \ix_single_ew[2][0] }));
 clb_tile \X[2].Y[1].clb  (.carry_in(\carry[1][2] ),
    .carry_out(\carry[2][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][2] ),
    .set_out_hard(\col_set[2][2] ),
    .shift_in_hard(\col_shift[1][2] ),
    .shift_out_hard(\col_shift[2][2] ),
    .cb_east_in({\dc_ew[11][4] ,
    \dc_ew[11][3] ,
    \dc_ew[11][2] ,
    \dc_ew[11][1] ,
    \dc_ew[11][0] }),
    .cb_east_out({\dc_we[11][9] ,
    \dc_we[11][8] ,
    \dc_we[11][7] ,
    \dc_we[11][6] ,
    \dc_we[11][5] ,
    \dc_we[11][4] ,
    \dc_we[11][3] ,
    \dc_we[11][2] ,
    \dc_we[11][1] ,
    \dc_we[11][0] }),
    .cb_north_in({\dc_ns[16][4] ,
    \dc_ns[16][3] ,
    \dc_ns[16][2] ,
    \dc_ns[16][1] ,
    \dc_ns[16][0] }),
    .cb_north_out({\dc_sn[16][9] ,
    \dc_sn[16][8] ,
    \dc_sn[16][7] ,
    \dc_sn[16][6] ,
    \dc_sn[16][5] ,
    \dc_sn[16][4] ,
    \dc_sn[16][3] ,
    \dc_sn[16][2] ,
    \dc_sn[16][1] ,
    \dc_sn[16][0] }),
    .clb_south_in({\dc_sn[9][9] ,
    \dc_sn[9][8] ,
    \dc_sn[9][7] ,
    \dc_sn[9][6] ,
    \dc_sn[9][5] ,
    \dc_sn[9][4] ,
    \dc_sn[9][3] ,
    \dc_sn[9][2] ,
    \dc_sn[9][1] ,
    \dc_sn[9][0] }),
    .clb_south_out({\dc_ns[9][4] ,
    \dc_ns[9][3] ,
    \dc_ns[9][2] ,
    \dc_ns[9][1] ,
    \dc_ns[9][0] }),
    .clb_west_in({\dc_we[10][9] ,
    \dc_we[10][8] ,
    \dc_we[10][7] ,
    \dc_we[10][6] ,
    \dc_we[10][5] ,
    \dc_we[10][4] ,
    \dc_we[10][3] ,
    \dc_we[10][2] ,
    \dc_we[10][1] ,
    \dc_we[10][0] }),
    .clb_west_out({\dc_ew[10][4] ,
    \dc_ew[10][3] ,
    \dc_ew[10][2] ,
    \dc_ew[10][1] ,
    \dc_ew[10][0] }),
    .east_double({\ix_double_ew[11][7] ,
    \ix_double_ew[11][6] ,
    \ix_double_ew[11][5] ,
    \ix_double_ew[11][4] ,
    \ix_double_ew[11][3] ,
    \ix_double_ew[11][2] ,
    \ix_double_ew[11][1] ,
    \ix_double_ew[11][0] }),
    .east_single({\ix_single_ew[11][3] ,
    \ix_single_ew[11][2] ,
    \ix_single_ew[11][1] ,
    \ix_single_ew[11][0] }),
    .north_double({\ix_double_ns[16][7] ,
    \ix_double_ns[16][6] ,
    \ix_double_ns[16][5] ,
    \ix_double_ns[16][4] ,
    \ix_double_ns[16][3] ,
    \ix_double_ns[16][2] ,
    \ix_double_ns[16][1] ,
    \ix_double_ns[16][0] }),
    .north_single({\ix_single_ns[16][3] ,
    \ix_single_ns[16][2] ,
    \ix_single_ns[16][1] ,
    \ix_single_ns[16][0] }),
    .south_double({\ix_double_ns[9][7] ,
    \ix_double_ns[9][6] ,
    \ix_double_ns[9][5] ,
    \ix_double_ns[9][4] ,
    \ix_double_ns[9][3] ,
    \ix_double_ns[9][2] ,
    \ix_double_ns[9][1] ,
    \ix_double_ns[9][0] }),
    .south_single({\ix_single_ns[9][3] ,
    \ix_single_ns[9][2] ,
    \ix_single_ns[9][1] ,
    \ix_single_ns[9][0] }),
    .west_double({\ix_double_ew[10][7] ,
    \ix_double_ew[10][6] ,
    \ix_double_ew[10][5] ,
    \ix_double_ew[10][4] ,
    \ix_double_ew[10][3] ,
    \ix_double_ew[10][2] ,
    \ix_double_ew[10][1] ,
    \ix_double_ew[10][0] }),
    .west_single({\ix_single_ew[10][3] ,
    \ix_single_ew[10][2] ,
    \ix_single_ew[10][1] ,
    \ix_single_ew[10][0] }));
 clb_tile \X[2].Y[2].clb  (.carry_in(\carry[2][2] ),
    .carry_out(\carry[3][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][2] ),
    .set_out_hard(\col_set[3][2] ),
    .shift_in_hard(\col_shift[2][2] ),
    .shift_out_hard(\col_shift[3][2] ),
    .cb_east_in({\dc_ew[19][4] ,
    \dc_ew[19][3] ,
    \dc_ew[19][2] ,
    \dc_ew[19][1] ,
    \dc_ew[19][0] }),
    .cb_east_out({\dc_we[19][9] ,
    \dc_we[19][8] ,
    \dc_we[19][7] ,
    \dc_we[19][6] ,
    \dc_we[19][5] ,
    \dc_we[19][4] ,
    \dc_we[19][3] ,
    \dc_we[19][2] ,
    \dc_we[19][1] ,
    \dc_we[19][0] }),
    .cb_north_in({\dc_ns[23][4] ,
    \dc_ns[23][3] ,
    \dc_ns[23][2] ,
    \dc_ns[23][1] ,
    \dc_ns[23][0] }),
    .cb_north_out({\dc_sn[23][9] ,
    \dc_sn[23][8] ,
    \dc_sn[23][7] ,
    \dc_sn[23][6] ,
    \dc_sn[23][5] ,
    \dc_sn[23][4] ,
    \dc_sn[23][3] ,
    \dc_sn[23][2] ,
    \dc_sn[23][1] ,
    \dc_sn[23][0] }),
    .clb_south_in({\dc_sn[16][9] ,
    \dc_sn[16][8] ,
    \dc_sn[16][7] ,
    \dc_sn[16][6] ,
    \dc_sn[16][5] ,
    \dc_sn[16][4] ,
    \dc_sn[16][3] ,
    \dc_sn[16][2] ,
    \dc_sn[16][1] ,
    \dc_sn[16][0] }),
    .clb_south_out({\dc_ns[16][4] ,
    \dc_ns[16][3] ,
    \dc_ns[16][2] ,
    \dc_ns[16][1] ,
    \dc_ns[16][0] }),
    .clb_west_in({\dc_we[18][9] ,
    \dc_we[18][8] ,
    \dc_we[18][7] ,
    \dc_we[18][6] ,
    \dc_we[18][5] ,
    \dc_we[18][4] ,
    \dc_we[18][3] ,
    \dc_we[18][2] ,
    \dc_we[18][1] ,
    \dc_we[18][0] }),
    .clb_west_out({\dc_ew[18][4] ,
    \dc_ew[18][3] ,
    \dc_ew[18][2] ,
    \dc_ew[18][1] ,
    \dc_ew[18][0] }),
    .east_double({\ix_double_ew[19][7] ,
    \ix_double_ew[19][6] ,
    \ix_double_ew[19][5] ,
    \ix_double_ew[19][4] ,
    \ix_double_ew[19][3] ,
    \ix_double_ew[19][2] ,
    \ix_double_ew[19][1] ,
    \ix_double_ew[19][0] }),
    .east_single({\ix_single_ew[19][3] ,
    \ix_single_ew[19][2] ,
    \ix_single_ew[19][1] ,
    \ix_single_ew[19][0] }),
    .north_double({\ix_double_ns[23][7] ,
    \ix_double_ns[23][6] ,
    \ix_double_ns[23][5] ,
    \ix_double_ns[23][4] ,
    \ix_double_ns[23][3] ,
    \ix_double_ns[23][2] ,
    \ix_double_ns[23][1] ,
    \ix_double_ns[23][0] }),
    .north_single({\ix_single_ns[23][3] ,
    \ix_single_ns[23][2] ,
    \ix_single_ns[23][1] ,
    \ix_single_ns[23][0] }),
    .south_double({\ix_double_ns[16][7] ,
    \ix_double_ns[16][6] ,
    \ix_double_ns[16][5] ,
    \ix_double_ns[16][4] ,
    \ix_double_ns[16][3] ,
    \ix_double_ns[16][2] ,
    \ix_double_ns[16][1] ,
    \ix_double_ns[16][0] }),
    .south_single({\ix_single_ns[16][3] ,
    \ix_single_ns[16][2] ,
    \ix_single_ns[16][1] ,
    \ix_single_ns[16][0] }),
    .west_double({\ix_double_ew[18][7] ,
    \ix_double_ew[18][6] ,
    \ix_double_ew[18][5] ,
    \ix_double_ew[18][4] ,
    \ix_double_ew[18][3] ,
    \ix_double_ew[18][2] ,
    \ix_double_ew[18][1] ,
    \ix_double_ew[18][0] }),
    .west_single({\ix_single_ew[18][3] ,
    \ix_single_ew[18][2] ,
    \ix_single_ew[18][1] ,
    \ix_single_ew[18][0] }));
 clb_tile \X[2].Y[3].clb  (.carry_in(\carry[3][2] ),
    .carry_out(\carry[4][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][2] ),
    .set_out_hard(\col_set[4][2] ),
    .shift_in_hard(\col_shift[3][2] ),
    .shift_out_hard(\col_shift[4][2] ),
    .cb_east_in({\dc_ew[27][4] ,
    \dc_ew[27][3] ,
    \dc_ew[27][2] ,
    \dc_ew[27][1] ,
    \dc_ew[27][0] }),
    .cb_east_out({\dc_we[27][9] ,
    \dc_we[27][8] ,
    \dc_we[27][7] ,
    \dc_we[27][6] ,
    \dc_we[27][5] ,
    \dc_we[27][4] ,
    \dc_we[27][3] ,
    \dc_we[27][2] ,
    \dc_we[27][1] ,
    \dc_we[27][0] }),
    .cb_north_in({\dc_ns[30][4] ,
    \dc_ns[30][3] ,
    \dc_ns[30][2] ,
    \dc_ns[30][1] ,
    \dc_ns[30][0] }),
    .cb_north_out({\dc_sn[30][9] ,
    \dc_sn[30][8] ,
    \dc_sn[30][7] ,
    \dc_sn[30][6] ,
    \dc_sn[30][5] ,
    \dc_sn[30][4] ,
    \dc_sn[30][3] ,
    \dc_sn[30][2] ,
    \dc_sn[30][1] ,
    \dc_sn[30][0] }),
    .clb_south_in({\dc_sn[23][9] ,
    \dc_sn[23][8] ,
    \dc_sn[23][7] ,
    \dc_sn[23][6] ,
    \dc_sn[23][5] ,
    \dc_sn[23][4] ,
    \dc_sn[23][3] ,
    \dc_sn[23][2] ,
    \dc_sn[23][1] ,
    \dc_sn[23][0] }),
    .clb_south_out({\dc_ns[23][4] ,
    \dc_ns[23][3] ,
    \dc_ns[23][2] ,
    \dc_ns[23][1] ,
    \dc_ns[23][0] }),
    .clb_west_in({\dc_we[26][9] ,
    \dc_we[26][8] ,
    \dc_we[26][7] ,
    \dc_we[26][6] ,
    \dc_we[26][5] ,
    \dc_we[26][4] ,
    \dc_we[26][3] ,
    \dc_we[26][2] ,
    \dc_we[26][1] ,
    \dc_we[26][0] }),
    .clb_west_out({\dc_ew[26][4] ,
    \dc_ew[26][3] ,
    \dc_ew[26][2] ,
    \dc_ew[26][1] ,
    \dc_ew[26][0] }),
    .east_double({\ix_double_ew[27][7] ,
    \ix_double_ew[27][6] ,
    \ix_double_ew[27][5] ,
    \ix_double_ew[27][4] ,
    \ix_double_ew[27][3] ,
    \ix_double_ew[27][2] ,
    \ix_double_ew[27][1] ,
    \ix_double_ew[27][0] }),
    .east_single({\ix_single_ew[27][3] ,
    \ix_single_ew[27][2] ,
    \ix_single_ew[27][1] ,
    \ix_single_ew[27][0] }),
    .north_double({\ix_double_ns[30][7] ,
    \ix_double_ns[30][6] ,
    \ix_double_ns[30][5] ,
    \ix_double_ns[30][4] ,
    \ix_double_ns[30][3] ,
    \ix_double_ns[30][2] ,
    \ix_double_ns[30][1] ,
    \ix_double_ns[30][0] }),
    .north_single({\ix_single_ns[30][3] ,
    \ix_single_ns[30][2] ,
    \ix_single_ns[30][1] ,
    \ix_single_ns[30][0] }),
    .south_double({\ix_double_ns[23][7] ,
    \ix_double_ns[23][6] ,
    \ix_double_ns[23][5] ,
    \ix_double_ns[23][4] ,
    \ix_double_ns[23][3] ,
    \ix_double_ns[23][2] ,
    \ix_double_ns[23][1] ,
    \ix_double_ns[23][0] }),
    .south_single({\ix_single_ns[23][3] ,
    \ix_single_ns[23][2] ,
    \ix_single_ns[23][1] ,
    \ix_single_ns[23][0] }),
    .west_double({\ix_double_ew[26][7] ,
    \ix_double_ew[26][6] ,
    \ix_double_ew[26][5] ,
    \ix_double_ew[26][4] ,
    \ix_double_ew[26][3] ,
    \ix_double_ew[26][2] ,
    \ix_double_ew[26][1] ,
    \ix_double_ew[26][0] }),
    .west_single({\ix_single_ew[26][3] ,
    \ix_single_ew[26][2] ,
    \ix_single_ew[26][1] ,
    \ix_single_ew[26][0] }));
 clb_tile \X[2].Y[4].clb  (.carry_in(\carry[4][2] ),
    .carry_out(\carry[5][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][2] ),
    .set_out_hard(\col_set[5][2] ),
    .shift_in_hard(\col_shift[4][2] ),
    .shift_out_hard(\col_shift[5][2] ),
    .cb_east_in({\dc_ew[35][4] ,
    \dc_ew[35][3] ,
    \dc_ew[35][2] ,
    \dc_ew[35][1] ,
    \dc_ew[35][0] }),
    .cb_east_out({\dc_we[35][9] ,
    \dc_we[35][8] ,
    \dc_we[35][7] ,
    \dc_we[35][6] ,
    \dc_we[35][5] ,
    \dc_we[35][4] ,
    \dc_we[35][3] ,
    \dc_we[35][2] ,
    \dc_we[35][1] ,
    \dc_we[35][0] }),
    .cb_north_in({\dc_ns[37][4] ,
    \dc_ns[37][3] ,
    \dc_ns[37][2] ,
    \dc_ns[37][1] ,
    \dc_ns[37][0] }),
    .cb_north_out({\dc_sn[37][9] ,
    \dc_sn[37][8] ,
    \dc_sn[37][7] ,
    \dc_sn[37][6] ,
    \dc_sn[37][5] ,
    \dc_sn[37][4] ,
    \dc_sn[37][3] ,
    \dc_sn[37][2] ,
    \dc_sn[37][1] ,
    \dc_sn[37][0] }),
    .clb_south_in({\dc_sn[30][9] ,
    \dc_sn[30][8] ,
    \dc_sn[30][7] ,
    \dc_sn[30][6] ,
    \dc_sn[30][5] ,
    \dc_sn[30][4] ,
    \dc_sn[30][3] ,
    \dc_sn[30][2] ,
    \dc_sn[30][1] ,
    \dc_sn[30][0] }),
    .clb_south_out({\dc_ns[30][4] ,
    \dc_ns[30][3] ,
    \dc_ns[30][2] ,
    \dc_ns[30][1] ,
    \dc_ns[30][0] }),
    .clb_west_in({\dc_we[34][9] ,
    \dc_we[34][8] ,
    \dc_we[34][7] ,
    \dc_we[34][6] ,
    \dc_we[34][5] ,
    \dc_we[34][4] ,
    \dc_we[34][3] ,
    \dc_we[34][2] ,
    \dc_we[34][1] ,
    \dc_we[34][0] }),
    .clb_west_out({\dc_ew[34][4] ,
    \dc_ew[34][3] ,
    \dc_ew[34][2] ,
    \dc_ew[34][1] ,
    \dc_ew[34][0] }),
    .east_double({\ix_double_ew[35][7] ,
    \ix_double_ew[35][6] ,
    \ix_double_ew[35][5] ,
    \ix_double_ew[35][4] ,
    \ix_double_ew[35][3] ,
    \ix_double_ew[35][2] ,
    \ix_double_ew[35][1] ,
    \ix_double_ew[35][0] }),
    .east_single({\ix_single_ew[35][3] ,
    \ix_single_ew[35][2] ,
    \ix_single_ew[35][1] ,
    \ix_single_ew[35][0] }),
    .north_double({\ix_double_ns[37][7] ,
    \ix_double_ns[37][6] ,
    \ix_double_ns[37][5] ,
    \ix_double_ns[37][4] ,
    \ix_double_ns[37][3] ,
    \ix_double_ns[37][2] ,
    \ix_double_ns[37][1] ,
    \ix_double_ns[37][0] }),
    .north_single({\ix_single_ns[37][3] ,
    \ix_single_ns[37][2] ,
    \ix_single_ns[37][1] ,
    \ix_single_ns[37][0] }),
    .south_double({\ix_double_ns[30][7] ,
    \ix_double_ns[30][6] ,
    \ix_double_ns[30][5] ,
    \ix_double_ns[30][4] ,
    \ix_double_ns[30][3] ,
    \ix_double_ns[30][2] ,
    \ix_double_ns[30][1] ,
    \ix_double_ns[30][0] }),
    .south_single({\ix_single_ns[30][3] ,
    \ix_single_ns[30][2] ,
    \ix_single_ns[30][1] ,
    \ix_single_ns[30][0] }),
    .west_double({\ix_double_ew[34][7] ,
    \ix_double_ew[34][6] ,
    \ix_double_ew[34][5] ,
    \ix_double_ew[34][4] ,
    \ix_double_ew[34][3] ,
    \ix_double_ew[34][2] ,
    \ix_double_ew[34][1] ,
    \ix_double_ew[34][0] }),
    .west_single({\ix_single_ew[34][3] ,
    \ix_single_ew[34][2] ,
    \ix_single_ew[34][1] ,
    \ix_single_ew[34][0] }));
 clb_tile \X[2].Y[5].clb  (.carry_in(\carry[5][2] ),
    .carry_out(\carry[6][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][2] ),
    .set_out_hard(\col_set[6][2] ),
    .shift_in_hard(\col_shift[5][2] ),
    .shift_out_hard(\col_shift[6][2] ),
    .cb_east_in({\dc_ew[43][4] ,
    \dc_ew[43][3] ,
    \dc_ew[43][2] ,
    \dc_ew[43][1] ,
    \dc_ew[43][0] }),
    .cb_east_out({\dc_we[43][9] ,
    \dc_we[43][8] ,
    \dc_we[43][7] ,
    \dc_we[43][6] ,
    \dc_we[43][5] ,
    \dc_we[43][4] ,
    \dc_we[43][3] ,
    \dc_we[43][2] ,
    \dc_we[43][1] ,
    \dc_we[43][0] }),
    .cb_north_in({\dc_ns[44][4] ,
    \dc_ns[44][3] ,
    \dc_ns[44][2] ,
    \dc_ns[44][1] ,
    \dc_ns[44][0] }),
    .cb_north_out({\dc_sn[44][9] ,
    \dc_sn[44][8] ,
    \dc_sn[44][7] ,
    \dc_sn[44][6] ,
    \dc_sn[44][5] ,
    \dc_sn[44][4] ,
    \dc_sn[44][3] ,
    \dc_sn[44][2] ,
    \dc_sn[44][1] ,
    \dc_sn[44][0] }),
    .clb_south_in({\dc_sn[37][9] ,
    \dc_sn[37][8] ,
    \dc_sn[37][7] ,
    \dc_sn[37][6] ,
    \dc_sn[37][5] ,
    \dc_sn[37][4] ,
    \dc_sn[37][3] ,
    \dc_sn[37][2] ,
    \dc_sn[37][1] ,
    \dc_sn[37][0] }),
    .clb_south_out({\dc_ns[37][4] ,
    \dc_ns[37][3] ,
    \dc_ns[37][2] ,
    \dc_ns[37][1] ,
    \dc_ns[37][0] }),
    .clb_west_in({\dc_we[42][9] ,
    \dc_we[42][8] ,
    \dc_we[42][7] ,
    \dc_we[42][6] ,
    \dc_we[42][5] ,
    \dc_we[42][4] ,
    \dc_we[42][3] ,
    \dc_we[42][2] ,
    \dc_we[42][1] ,
    \dc_we[42][0] }),
    .clb_west_out({\dc_ew[42][4] ,
    \dc_ew[42][3] ,
    \dc_ew[42][2] ,
    \dc_ew[42][1] ,
    \dc_ew[42][0] }),
    .east_double({\ix_double_ew[43][7] ,
    \ix_double_ew[43][6] ,
    \ix_double_ew[43][5] ,
    \ix_double_ew[43][4] ,
    \ix_double_ew[43][3] ,
    \ix_double_ew[43][2] ,
    \ix_double_ew[43][1] ,
    \ix_double_ew[43][0] }),
    .east_single({\ix_single_ew[43][3] ,
    \ix_single_ew[43][2] ,
    \ix_single_ew[43][1] ,
    \ix_single_ew[43][0] }),
    .north_double({\ix_double_ns[44][7] ,
    \ix_double_ns[44][6] ,
    \ix_double_ns[44][5] ,
    \ix_double_ns[44][4] ,
    \ix_double_ns[44][3] ,
    \ix_double_ns[44][2] ,
    \ix_double_ns[44][1] ,
    \ix_double_ns[44][0] }),
    .north_single({\ix_single_ns[44][3] ,
    \ix_single_ns[44][2] ,
    \ix_single_ns[44][1] ,
    \ix_single_ns[44][0] }),
    .south_double({\ix_double_ns[37][7] ,
    \ix_double_ns[37][6] ,
    \ix_double_ns[37][5] ,
    \ix_double_ns[37][4] ,
    \ix_double_ns[37][3] ,
    \ix_double_ns[37][2] ,
    \ix_double_ns[37][1] ,
    \ix_double_ns[37][0] }),
    .south_single({\ix_single_ns[37][3] ,
    \ix_single_ns[37][2] ,
    \ix_single_ns[37][1] ,
    \ix_single_ns[37][0] }),
    .west_double({\ix_double_ew[42][7] ,
    \ix_double_ew[42][6] ,
    \ix_double_ew[42][5] ,
    \ix_double_ew[42][4] ,
    \ix_double_ew[42][3] ,
    \ix_double_ew[42][2] ,
    \ix_double_ew[42][1] ,
    \ix_double_ew[42][0] }),
    .west_single({\ix_single_ew[42][3] ,
    \ix_single_ew[42][2] ,
    \ix_single_ew[42][1] ,
    \ix_single_ew[42][0] }));
 clb_tile \X[2].Y[6].clb  (.carry_in(\carry[6][2] ),
    .carry_out(\carry[7][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][2] ),
    .set_out_hard(\col_set[7][2] ),
    .shift_in_hard(\col_shift[6][2] ),
    .shift_out_hard(\col_shift[7][2] ),
    .cb_east_in({\dc_ew[51][4] ,
    \dc_ew[51][3] ,
    \dc_ew[51][2] ,
    \dc_ew[51][1] ,
    \dc_ew[51][0] }),
    .cb_east_out({\dc_we[51][9] ,
    \dc_we[51][8] ,
    \dc_we[51][7] ,
    \dc_we[51][6] ,
    \dc_we[51][5] ,
    \dc_we[51][4] ,
    \dc_we[51][3] ,
    \dc_we[51][2] ,
    \dc_we[51][1] ,
    \dc_we[51][0] }),
    .cb_north_in({\dc_ns[51][4] ,
    \dc_ns[51][3] ,
    \dc_ns[51][2] ,
    \dc_ns[51][1] ,
    \dc_ns[51][0] }),
    .cb_north_out({\dc_sn[51][9] ,
    \dc_sn[51][8] ,
    \dc_sn[51][7] ,
    \dc_sn[51][6] ,
    \dc_sn[51][5] ,
    \dc_sn[51][4] ,
    \dc_sn[51][3] ,
    \dc_sn[51][2] ,
    \dc_sn[51][1] ,
    \dc_sn[51][0] }),
    .clb_south_in({\dc_sn[44][9] ,
    \dc_sn[44][8] ,
    \dc_sn[44][7] ,
    \dc_sn[44][6] ,
    \dc_sn[44][5] ,
    \dc_sn[44][4] ,
    \dc_sn[44][3] ,
    \dc_sn[44][2] ,
    \dc_sn[44][1] ,
    \dc_sn[44][0] }),
    .clb_south_out({\dc_ns[44][4] ,
    \dc_ns[44][3] ,
    \dc_ns[44][2] ,
    \dc_ns[44][1] ,
    \dc_ns[44][0] }),
    .clb_west_in({\dc_we[50][9] ,
    \dc_we[50][8] ,
    \dc_we[50][7] ,
    \dc_we[50][6] ,
    \dc_we[50][5] ,
    \dc_we[50][4] ,
    \dc_we[50][3] ,
    \dc_we[50][2] ,
    \dc_we[50][1] ,
    \dc_we[50][0] }),
    .clb_west_out({\dc_ew[50][4] ,
    \dc_ew[50][3] ,
    \dc_ew[50][2] ,
    \dc_ew[50][1] ,
    \dc_ew[50][0] }),
    .east_double({\ix_double_ew[51][7] ,
    \ix_double_ew[51][6] ,
    \ix_double_ew[51][5] ,
    \ix_double_ew[51][4] ,
    \ix_double_ew[51][3] ,
    \ix_double_ew[51][2] ,
    \ix_double_ew[51][1] ,
    \ix_double_ew[51][0] }),
    .east_single({\ix_single_ew[51][3] ,
    \ix_single_ew[51][2] ,
    \ix_single_ew[51][1] ,
    \ix_single_ew[51][0] }),
    .north_double({\ix_double_ns[51][7] ,
    \ix_double_ns[51][6] ,
    \ix_double_ns[51][5] ,
    \ix_double_ns[51][4] ,
    \ix_double_ns[51][3] ,
    \ix_double_ns[51][2] ,
    \ix_double_ns[51][1] ,
    \ix_double_ns[51][0] }),
    .north_single({\ix_single_ns[51][3] ,
    \ix_single_ns[51][2] ,
    \ix_single_ns[51][1] ,
    \ix_single_ns[51][0] }),
    .south_double({\ix_double_ns[44][7] ,
    \ix_double_ns[44][6] ,
    \ix_double_ns[44][5] ,
    \ix_double_ns[44][4] ,
    \ix_double_ns[44][3] ,
    \ix_double_ns[44][2] ,
    \ix_double_ns[44][1] ,
    \ix_double_ns[44][0] }),
    .south_single({\ix_single_ns[44][3] ,
    \ix_single_ns[44][2] ,
    \ix_single_ns[44][1] ,
    \ix_single_ns[44][0] }),
    .west_double({\ix_double_ew[50][7] ,
    \ix_double_ew[50][6] ,
    \ix_double_ew[50][5] ,
    \ix_double_ew[50][4] ,
    \ix_double_ew[50][3] ,
    \ix_double_ew[50][2] ,
    \ix_double_ew[50][1] ,
    \ix_double_ew[50][0] }),
    .west_single({\ix_single_ew[50][3] ,
    \ix_single_ew[50][2] ,
    \ix_single_ew[50][1] ,
    \ix_single_ew[50][0] }));
 clb_tile \X[2].Y[7].clb  (.carry_in(\carry[7][2] ),
    .carry_out(\carry[8][2] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][2] ),
    .set_out_hard(\col_set[8][2] ),
    .shift_in_hard(\col_shift[7][2] ),
    .shift_out_hard(\col_shift[8][2] ),
    .cb_east_in({\dc_ew[59][4] ,
    \dc_ew[59][3] ,
    \dc_ew[59][2] ,
    \dc_ew[59][1] ,
    \dc_ew[59][0] }),
    .cb_east_out({\dc_we[59][9] ,
    \dc_we[59][8] ,
    \dc_we[59][7] ,
    \dc_we[59][6] ,
    \dc_we[59][5] ,
    \dc_we[59][4] ,
    \dc_we[59][3] ,
    \dc_we[59][2] ,
    \dc_we[59][1] ,
    \dc_we[59][0] }),
    .cb_north_in({_127_,
    _126_,
    _125_,
    _124_,
    _123_}),
    .cb_north_out({\dc_sn[58][9] ,
    \dc_sn[58][8] ,
    \dc_sn[58][7] ,
    \dc_sn[58][6] ,
    \dc_sn[58][5] ,
    \dc_sn[58][4] ,
    \dc_sn[58][3] ,
    \dc_sn[58][2] ,
    \dc_sn[58][1] ,
    \dc_sn[58][0] }),
    .clb_south_in({\dc_sn[51][9] ,
    \dc_sn[51][8] ,
    \dc_sn[51][7] ,
    \dc_sn[51][6] ,
    \dc_sn[51][5] ,
    \dc_sn[51][4] ,
    \dc_sn[51][3] ,
    \dc_sn[51][2] ,
    \dc_sn[51][1] ,
    \dc_sn[51][0] }),
    .clb_south_out({\dc_ns[51][4] ,
    \dc_ns[51][3] ,
    \dc_ns[51][2] ,
    \dc_ns[51][1] ,
    \dc_ns[51][0] }),
    .clb_west_in({\dc_we[58][9] ,
    \dc_we[58][8] ,
    \dc_we[58][7] ,
    \dc_we[58][6] ,
    \dc_we[58][5] ,
    \dc_we[58][4] ,
    \dc_we[58][3] ,
    \dc_we[58][2] ,
    \dc_we[58][1] ,
    \dc_we[58][0] }),
    .clb_west_out({\dc_ew[58][4] ,
    \dc_ew[58][3] ,
    \dc_ew[58][2] ,
    \dc_ew[58][1] ,
    \dc_ew[58][0] }),
    .east_double({\ix_double_ew[59][7] ,
    \ix_double_ew[59][6] ,
    \ix_double_ew[59][5] ,
    \ix_double_ew[59][4] ,
    \ix_double_ew[59][3] ,
    \ix_double_ew[59][2] ,
    \ix_double_ew[59][1] ,
    \ix_double_ew[59][0] }),
    .east_single({\ix_single_ew[59][3] ,
    \ix_single_ew[59][2] ,
    \ix_single_ew[59][1] ,
    \ix_single_ew[59][0] }),
    .north_double({\ix_double_ns[58][7] ,
    \ix_double_ns[58][6] ,
    \ix_double_ns[58][5] ,
    \ix_double_ns[58][4] ,
    \ix_double_ns[58][3] ,
    \ix_double_ns[58][2] ,
    \ix_double_ns[58][1] ,
    \ix_double_ns[58][0] }),
    .north_single({\ix_single_ns[58][3] ,
    \ix_single_ns[58][2] ,
    \ix_single_ns[58][1] ,
    gpio_north[2]}),
    .south_double({\ix_double_ns[51][7] ,
    \ix_double_ns[51][6] ,
    \ix_double_ns[51][5] ,
    \ix_double_ns[51][4] ,
    \ix_double_ns[51][3] ,
    \ix_double_ns[51][2] ,
    \ix_double_ns[51][1] ,
    \ix_double_ns[51][0] }),
    .south_single({\ix_single_ns[51][3] ,
    \ix_single_ns[51][2] ,
    \ix_single_ns[51][1] ,
    \ix_single_ns[51][0] }),
    .west_double({\ix_double_ew[58][7] ,
    \ix_double_ew[58][6] ,
    \ix_double_ew[58][5] ,
    \ix_double_ew[58][4] ,
    \ix_double_ew[58][3] ,
    \ix_double_ew[58][2] ,
    \ix_double_ew[58][1] ,
    \ix_double_ew[58][0] }),
    .west_single({\ix_single_ew[58][3] ,
    \ix_single_ew[58][2] ,
    \ix_single_ew[58][1] ,
    \ix_single_ew[58][0] }));
 clb_tile \X[3].Y[0].clb  (.carry_in(_128_),
    .carry_out(\carry[1][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[0][3] ),
    .set_out_hard(\col_set[1][3] ),
    .shift_in_hard(\wb_shift_out[0][3] ),
    .shift_out_hard(\col_shift[1][3] ),
    .cb_east_in({\dc_ew[4][4] ,
    \dc_ew[4][3] ,
    \dc_ew[4][2] ,
    \dc_ew[4][1] ,
    \dc_ew[4][0] }),
    .cb_east_out({\dc_we[4][9] ,
    \dc_we[4][8] ,
    \dc_we[4][7] ,
    \dc_we[4][6] ,
    \dc_we[4][5] ,
    \dc_we[4][4] ,
    \dc_we[4][3] ,
    \dc_we[4][2] ,
    \dc_we[4][1] ,
    \dc_we[4][0] }),
    .cb_north_in({\dc_ns[10][4] ,
    \dc_ns[10][3] ,
    \dc_ns[10][2] ,
    \dc_ns[10][1] ,
    \dc_ns[10][0] }),
    .cb_north_out({\dc_sn[10][9] ,
    \dc_sn[10][8] ,
    \dc_sn[10][7] ,
    \dc_sn[10][6] ,
    \dc_sn[10][5] ,
    \dc_sn[10][4] ,
    \dc_sn[10][3] ,
    \dc_sn[10][2] ,
    \dc_sn[10][1] ,
    \dc_sn[10][0] }),
    .clb_south_in({_138_,
    _137_,
    _136_,
    _135_,
    _134_,
    _133_,
    _132_,
    _131_,
    _130_,
    _129_}),
    .clb_south_out({\dc_ns[3][4] ,
    \dc_ns[3][3] ,
    \dc_ns[3][2] ,
    \dc_ns[3][1] ,
    \dc_ns[3][0] }),
    .clb_west_in({\dc_we[3][9] ,
    \dc_we[3][8] ,
    \dc_we[3][7] ,
    \dc_we[3][6] ,
    \dc_we[3][5] ,
    \dc_we[3][4] ,
    \dc_we[3][3] ,
    \dc_we[3][2] ,
    \dc_we[3][1] ,
    \dc_we[3][0] }),
    .clb_west_out({\dc_ew[3][4] ,
    \dc_ew[3][3] ,
    \dc_ew[3][2] ,
    \dc_ew[3][1] ,
    \dc_ew[3][0] }),
    .east_double({\ix_double_ew[4][7] ,
    \ix_double_ew[4][6] ,
    \ix_double_ew[4][5] ,
    \ix_double_ew[4][4] ,
    \ix_double_ew[4][3] ,
    \ix_double_ew[4][2] ,
    \ix_double_ew[4][1] ,
    \ix_double_ew[4][0] }),
    .east_single({\ix_single_ew[4][3] ,
    \ix_single_ew[4][2] ,
    \ix_single_ew[4][1] ,
    \ix_single_ew[4][0] }),
    .north_double({\ix_double_ns[10][7] ,
    \ix_double_ns[10][6] ,
    \ix_double_ns[10][5] ,
    \ix_double_ns[10][4] ,
    \ix_double_ns[10][3] ,
    \ix_double_ns[10][2] ,
    \ix_double_ns[10][1] ,
    \ix_double_ns[10][0] }),
    .north_single({\ix_single_ns[10][3] ,
    \ix_single_ns[10][2] ,
    \ix_single_ns[10][1] ,
    \ix_single_ns[10][0] }),
    .south_double({\ix_double_ns[3][7] ,
    \ix_double_ns[3][6] ,
    \ix_double_ns[3][5] ,
    \ix_double_ns[3][4] ,
    \ix_double_ns[3][3] ,
    \ix_double_ns[3][2] ,
    \ix_double_ns[3][1] ,
    \ix_double_ns[3][0] }),
    .south_single({\ix_single_ns[3][3] ,
    \ix_single_ns[3][2] ,
    \ix_single_ns[3][1] ,
    gpio_south[3]}),
    .west_double({\ix_double_ew[3][7] ,
    \ix_double_ew[3][6] ,
    \ix_double_ew[3][5] ,
    \ix_double_ew[3][4] ,
    \ix_double_ew[3][3] ,
    \ix_double_ew[3][2] ,
    \ix_double_ew[3][1] ,
    \ix_double_ew[3][0] }),
    .west_single({\ix_single_ew[3][3] ,
    \ix_single_ew[3][2] ,
    \ix_single_ew[3][1] ,
    \ix_single_ew[3][0] }));
 clb_tile \X[3].Y[1].clb  (.carry_in(\carry[1][3] ),
    .carry_out(\carry[2][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][3] ),
    .set_out_hard(\col_set[2][3] ),
    .shift_in_hard(\col_shift[1][3] ),
    .shift_out_hard(\col_shift[2][3] ),
    .cb_east_in({\dc_ew[12][4] ,
    \dc_ew[12][3] ,
    \dc_ew[12][2] ,
    \dc_ew[12][1] ,
    \dc_ew[12][0] }),
    .cb_east_out({\dc_we[12][9] ,
    \dc_we[12][8] ,
    \dc_we[12][7] ,
    \dc_we[12][6] ,
    \dc_we[12][5] ,
    \dc_we[12][4] ,
    \dc_we[12][3] ,
    \dc_we[12][2] ,
    \dc_we[12][1] ,
    \dc_we[12][0] }),
    .cb_north_in({\dc_ns[17][4] ,
    \dc_ns[17][3] ,
    \dc_ns[17][2] ,
    \dc_ns[17][1] ,
    \dc_ns[17][0] }),
    .cb_north_out({\dc_sn[17][9] ,
    \dc_sn[17][8] ,
    \dc_sn[17][7] ,
    \dc_sn[17][6] ,
    \dc_sn[17][5] ,
    \dc_sn[17][4] ,
    \dc_sn[17][3] ,
    \dc_sn[17][2] ,
    \dc_sn[17][1] ,
    \dc_sn[17][0] }),
    .clb_south_in({\dc_sn[10][9] ,
    \dc_sn[10][8] ,
    \dc_sn[10][7] ,
    \dc_sn[10][6] ,
    \dc_sn[10][5] ,
    \dc_sn[10][4] ,
    \dc_sn[10][3] ,
    \dc_sn[10][2] ,
    \dc_sn[10][1] ,
    \dc_sn[10][0] }),
    .clb_south_out({\dc_ns[10][4] ,
    \dc_ns[10][3] ,
    \dc_ns[10][2] ,
    \dc_ns[10][1] ,
    \dc_ns[10][0] }),
    .clb_west_in({\dc_we[11][9] ,
    \dc_we[11][8] ,
    \dc_we[11][7] ,
    \dc_we[11][6] ,
    \dc_we[11][5] ,
    \dc_we[11][4] ,
    \dc_we[11][3] ,
    \dc_we[11][2] ,
    \dc_we[11][1] ,
    \dc_we[11][0] }),
    .clb_west_out({\dc_ew[11][4] ,
    \dc_ew[11][3] ,
    \dc_ew[11][2] ,
    \dc_ew[11][1] ,
    \dc_ew[11][0] }),
    .east_double({\ix_double_ew[12][7] ,
    \ix_double_ew[12][6] ,
    \ix_double_ew[12][5] ,
    \ix_double_ew[12][4] ,
    \ix_double_ew[12][3] ,
    \ix_double_ew[12][2] ,
    \ix_double_ew[12][1] ,
    \ix_double_ew[12][0] }),
    .east_single({\ix_single_ew[12][3] ,
    \ix_single_ew[12][2] ,
    \ix_single_ew[12][1] ,
    \ix_single_ew[12][0] }),
    .north_double({\ix_double_ns[17][7] ,
    \ix_double_ns[17][6] ,
    \ix_double_ns[17][5] ,
    \ix_double_ns[17][4] ,
    \ix_double_ns[17][3] ,
    \ix_double_ns[17][2] ,
    \ix_double_ns[17][1] ,
    \ix_double_ns[17][0] }),
    .north_single({\ix_single_ns[17][3] ,
    \ix_single_ns[17][2] ,
    \ix_single_ns[17][1] ,
    \ix_single_ns[17][0] }),
    .south_double({\ix_double_ns[10][7] ,
    \ix_double_ns[10][6] ,
    \ix_double_ns[10][5] ,
    \ix_double_ns[10][4] ,
    \ix_double_ns[10][3] ,
    \ix_double_ns[10][2] ,
    \ix_double_ns[10][1] ,
    \ix_double_ns[10][0] }),
    .south_single({\ix_single_ns[10][3] ,
    \ix_single_ns[10][2] ,
    \ix_single_ns[10][1] ,
    \ix_single_ns[10][0] }),
    .west_double({\ix_double_ew[11][7] ,
    \ix_double_ew[11][6] ,
    \ix_double_ew[11][5] ,
    \ix_double_ew[11][4] ,
    \ix_double_ew[11][3] ,
    \ix_double_ew[11][2] ,
    \ix_double_ew[11][1] ,
    \ix_double_ew[11][0] }),
    .west_single({\ix_single_ew[11][3] ,
    \ix_single_ew[11][2] ,
    \ix_single_ew[11][1] ,
    \ix_single_ew[11][0] }));
 clb_tile \X[3].Y[2].clb  (.carry_in(\carry[2][3] ),
    .carry_out(\carry[3][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][3] ),
    .set_out_hard(\col_set[3][3] ),
    .shift_in_hard(\col_shift[2][3] ),
    .shift_out_hard(\col_shift[3][3] ),
    .cb_east_in({\dc_ew[20][4] ,
    \dc_ew[20][3] ,
    \dc_ew[20][2] ,
    \dc_ew[20][1] ,
    \dc_ew[20][0] }),
    .cb_east_out({\dc_we[20][9] ,
    \dc_we[20][8] ,
    \dc_we[20][7] ,
    \dc_we[20][6] ,
    \dc_we[20][5] ,
    \dc_we[20][4] ,
    \dc_we[20][3] ,
    \dc_we[20][2] ,
    \dc_we[20][1] ,
    \dc_we[20][0] }),
    .cb_north_in({\dc_ns[24][4] ,
    \dc_ns[24][3] ,
    \dc_ns[24][2] ,
    \dc_ns[24][1] ,
    \dc_ns[24][0] }),
    .cb_north_out({\dc_sn[24][9] ,
    \dc_sn[24][8] ,
    \dc_sn[24][7] ,
    \dc_sn[24][6] ,
    \dc_sn[24][5] ,
    \dc_sn[24][4] ,
    \dc_sn[24][3] ,
    \dc_sn[24][2] ,
    \dc_sn[24][1] ,
    \dc_sn[24][0] }),
    .clb_south_in({\dc_sn[17][9] ,
    \dc_sn[17][8] ,
    \dc_sn[17][7] ,
    \dc_sn[17][6] ,
    \dc_sn[17][5] ,
    \dc_sn[17][4] ,
    \dc_sn[17][3] ,
    \dc_sn[17][2] ,
    \dc_sn[17][1] ,
    \dc_sn[17][0] }),
    .clb_south_out({\dc_ns[17][4] ,
    \dc_ns[17][3] ,
    \dc_ns[17][2] ,
    \dc_ns[17][1] ,
    \dc_ns[17][0] }),
    .clb_west_in({\dc_we[19][9] ,
    \dc_we[19][8] ,
    \dc_we[19][7] ,
    \dc_we[19][6] ,
    \dc_we[19][5] ,
    \dc_we[19][4] ,
    \dc_we[19][3] ,
    \dc_we[19][2] ,
    \dc_we[19][1] ,
    \dc_we[19][0] }),
    .clb_west_out({\dc_ew[19][4] ,
    \dc_ew[19][3] ,
    \dc_ew[19][2] ,
    \dc_ew[19][1] ,
    \dc_ew[19][0] }),
    .east_double({\ix_double_ew[20][7] ,
    \ix_double_ew[20][6] ,
    \ix_double_ew[20][5] ,
    \ix_double_ew[20][4] ,
    \ix_double_ew[20][3] ,
    \ix_double_ew[20][2] ,
    \ix_double_ew[20][1] ,
    \ix_double_ew[20][0] }),
    .east_single({\ix_single_ew[20][3] ,
    \ix_single_ew[20][2] ,
    \ix_single_ew[20][1] ,
    \ix_single_ew[20][0] }),
    .north_double({\ix_double_ns[24][7] ,
    \ix_double_ns[24][6] ,
    \ix_double_ns[24][5] ,
    \ix_double_ns[24][4] ,
    \ix_double_ns[24][3] ,
    \ix_double_ns[24][2] ,
    \ix_double_ns[24][1] ,
    \ix_double_ns[24][0] }),
    .north_single({\ix_single_ns[24][3] ,
    \ix_single_ns[24][2] ,
    \ix_single_ns[24][1] ,
    \ix_single_ns[24][0] }),
    .south_double({\ix_double_ns[17][7] ,
    \ix_double_ns[17][6] ,
    \ix_double_ns[17][5] ,
    \ix_double_ns[17][4] ,
    \ix_double_ns[17][3] ,
    \ix_double_ns[17][2] ,
    \ix_double_ns[17][1] ,
    \ix_double_ns[17][0] }),
    .south_single({\ix_single_ns[17][3] ,
    \ix_single_ns[17][2] ,
    \ix_single_ns[17][1] ,
    \ix_single_ns[17][0] }),
    .west_double({\ix_double_ew[19][7] ,
    \ix_double_ew[19][6] ,
    \ix_double_ew[19][5] ,
    \ix_double_ew[19][4] ,
    \ix_double_ew[19][3] ,
    \ix_double_ew[19][2] ,
    \ix_double_ew[19][1] ,
    \ix_double_ew[19][0] }),
    .west_single({\ix_single_ew[19][3] ,
    \ix_single_ew[19][2] ,
    \ix_single_ew[19][1] ,
    \ix_single_ew[19][0] }));
 clb_tile \X[3].Y[3].clb  (.carry_in(\carry[3][3] ),
    .carry_out(\carry[4][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][3] ),
    .set_out_hard(\col_set[4][3] ),
    .shift_in_hard(\col_shift[3][3] ),
    .shift_out_hard(\col_shift[4][3] ),
    .cb_east_in({\dc_ew[28][4] ,
    \dc_ew[28][3] ,
    \dc_ew[28][2] ,
    \dc_ew[28][1] ,
    \dc_ew[28][0] }),
    .cb_east_out({\dc_we[28][9] ,
    \dc_we[28][8] ,
    \dc_we[28][7] ,
    \dc_we[28][6] ,
    \dc_we[28][5] ,
    \dc_we[28][4] ,
    \dc_we[28][3] ,
    \dc_we[28][2] ,
    \dc_we[28][1] ,
    \dc_we[28][0] }),
    .cb_north_in({\dc_ns[31][4] ,
    \dc_ns[31][3] ,
    \dc_ns[31][2] ,
    \dc_ns[31][1] ,
    \dc_ns[31][0] }),
    .cb_north_out({\dc_sn[31][9] ,
    \dc_sn[31][8] ,
    \dc_sn[31][7] ,
    \dc_sn[31][6] ,
    \dc_sn[31][5] ,
    \dc_sn[31][4] ,
    \dc_sn[31][3] ,
    \dc_sn[31][2] ,
    \dc_sn[31][1] ,
    \dc_sn[31][0] }),
    .clb_south_in({\dc_sn[24][9] ,
    \dc_sn[24][8] ,
    \dc_sn[24][7] ,
    \dc_sn[24][6] ,
    \dc_sn[24][5] ,
    \dc_sn[24][4] ,
    \dc_sn[24][3] ,
    \dc_sn[24][2] ,
    \dc_sn[24][1] ,
    \dc_sn[24][0] }),
    .clb_south_out({\dc_ns[24][4] ,
    \dc_ns[24][3] ,
    \dc_ns[24][2] ,
    \dc_ns[24][1] ,
    \dc_ns[24][0] }),
    .clb_west_in({\dc_we[27][9] ,
    \dc_we[27][8] ,
    \dc_we[27][7] ,
    \dc_we[27][6] ,
    \dc_we[27][5] ,
    \dc_we[27][4] ,
    \dc_we[27][3] ,
    \dc_we[27][2] ,
    \dc_we[27][1] ,
    \dc_we[27][0] }),
    .clb_west_out({\dc_ew[27][4] ,
    \dc_ew[27][3] ,
    \dc_ew[27][2] ,
    \dc_ew[27][1] ,
    \dc_ew[27][0] }),
    .east_double({\ix_double_ew[28][7] ,
    \ix_double_ew[28][6] ,
    \ix_double_ew[28][5] ,
    \ix_double_ew[28][4] ,
    \ix_double_ew[28][3] ,
    \ix_double_ew[28][2] ,
    \ix_double_ew[28][1] ,
    \ix_double_ew[28][0] }),
    .east_single({\ix_single_ew[28][3] ,
    \ix_single_ew[28][2] ,
    \ix_single_ew[28][1] ,
    \ix_single_ew[28][0] }),
    .north_double({\ix_double_ns[31][7] ,
    \ix_double_ns[31][6] ,
    \ix_double_ns[31][5] ,
    \ix_double_ns[31][4] ,
    \ix_double_ns[31][3] ,
    \ix_double_ns[31][2] ,
    \ix_double_ns[31][1] ,
    \ix_double_ns[31][0] }),
    .north_single({\ix_single_ns[31][3] ,
    \ix_single_ns[31][2] ,
    \ix_single_ns[31][1] ,
    \ix_single_ns[31][0] }),
    .south_double({\ix_double_ns[24][7] ,
    \ix_double_ns[24][6] ,
    \ix_double_ns[24][5] ,
    \ix_double_ns[24][4] ,
    \ix_double_ns[24][3] ,
    \ix_double_ns[24][2] ,
    \ix_double_ns[24][1] ,
    \ix_double_ns[24][0] }),
    .south_single({\ix_single_ns[24][3] ,
    \ix_single_ns[24][2] ,
    \ix_single_ns[24][1] ,
    \ix_single_ns[24][0] }),
    .west_double({\ix_double_ew[27][7] ,
    \ix_double_ew[27][6] ,
    \ix_double_ew[27][5] ,
    \ix_double_ew[27][4] ,
    \ix_double_ew[27][3] ,
    \ix_double_ew[27][2] ,
    \ix_double_ew[27][1] ,
    \ix_double_ew[27][0] }),
    .west_single({\ix_single_ew[27][3] ,
    \ix_single_ew[27][2] ,
    \ix_single_ew[27][1] ,
    \ix_single_ew[27][0] }));
 clb_tile \X[3].Y[4].clb  (.carry_in(\carry[4][3] ),
    .carry_out(\carry[5][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][3] ),
    .set_out_hard(\col_set[5][3] ),
    .shift_in_hard(\col_shift[4][3] ),
    .shift_out_hard(\col_shift[5][3] ),
    .cb_east_in({\dc_ew[36][4] ,
    \dc_ew[36][3] ,
    \dc_ew[36][2] ,
    \dc_ew[36][1] ,
    \dc_ew[36][0] }),
    .cb_east_out({\dc_we[36][9] ,
    \dc_we[36][8] ,
    \dc_we[36][7] ,
    \dc_we[36][6] ,
    \dc_we[36][5] ,
    \dc_we[36][4] ,
    \dc_we[36][3] ,
    \dc_we[36][2] ,
    \dc_we[36][1] ,
    \dc_we[36][0] }),
    .cb_north_in({\dc_ns[38][4] ,
    \dc_ns[38][3] ,
    \dc_ns[38][2] ,
    \dc_ns[38][1] ,
    \dc_ns[38][0] }),
    .cb_north_out({\dc_sn[38][9] ,
    \dc_sn[38][8] ,
    \dc_sn[38][7] ,
    \dc_sn[38][6] ,
    \dc_sn[38][5] ,
    \dc_sn[38][4] ,
    \dc_sn[38][3] ,
    \dc_sn[38][2] ,
    \dc_sn[38][1] ,
    \dc_sn[38][0] }),
    .clb_south_in({\dc_sn[31][9] ,
    \dc_sn[31][8] ,
    \dc_sn[31][7] ,
    \dc_sn[31][6] ,
    \dc_sn[31][5] ,
    \dc_sn[31][4] ,
    \dc_sn[31][3] ,
    \dc_sn[31][2] ,
    \dc_sn[31][1] ,
    \dc_sn[31][0] }),
    .clb_south_out({\dc_ns[31][4] ,
    \dc_ns[31][3] ,
    \dc_ns[31][2] ,
    \dc_ns[31][1] ,
    \dc_ns[31][0] }),
    .clb_west_in({\dc_we[35][9] ,
    \dc_we[35][8] ,
    \dc_we[35][7] ,
    \dc_we[35][6] ,
    \dc_we[35][5] ,
    \dc_we[35][4] ,
    \dc_we[35][3] ,
    \dc_we[35][2] ,
    \dc_we[35][1] ,
    \dc_we[35][0] }),
    .clb_west_out({\dc_ew[35][4] ,
    \dc_ew[35][3] ,
    \dc_ew[35][2] ,
    \dc_ew[35][1] ,
    \dc_ew[35][0] }),
    .east_double({\ix_double_ew[36][7] ,
    \ix_double_ew[36][6] ,
    \ix_double_ew[36][5] ,
    \ix_double_ew[36][4] ,
    \ix_double_ew[36][3] ,
    \ix_double_ew[36][2] ,
    \ix_double_ew[36][1] ,
    \ix_double_ew[36][0] }),
    .east_single({\ix_single_ew[36][3] ,
    \ix_single_ew[36][2] ,
    \ix_single_ew[36][1] ,
    \ix_single_ew[36][0] }),
    .north_double({\ix_double_ns[38][7] ,
    \ix_double_ns[38][6] ,
    \ix_double_ns[38][5] ,
    \ix_double_ns[38][4] ,
    \ix_double_ns[38][3] ,
    \ix_double_ns[38][2] ,
    \ix_double_ns[38][1] ,
    \ix_double_ns[38][0] }),
    .north_single({\ix_single_ns[38][3] ,
    \ix_single_ns[38][2] ,
    \ix_single_ns[38][1] ,
    \ix_single_ns[38][0] }),
    .south_double({\ix_double_ns[31][7] ,
    \ix_double_ns[31][6] ,
    \ix_double_ns[31][5] ,
    \ix_double_ns[31][4] ,
    \ix_double_ns[31][3] ,
    \ix_double_ns[31][2] ,
    \ix_double_ns[31][1] ,
    \ix_double_ns[31][0] }),
    .south_single({\ix_single_ns[31][3] ,
    \ix_single_ns[31][2] ,
    \ix_single_ns[31][1] ,
    \ix_single_ns[31][0] }),
    .west_double({\ix_double_ew[35][7] ,
    \ix_double_ew[35][6] ,
    \ix_double_ew[35][5] ,
    \ix_double_ew[35][4] ,
    \ix_double_ew[35][3] ,
    \ix_double_ew[35][2] ,
    \ix_double_ew[35][1] ,
    \ix_double_ew[35][0] }),
    .west_single({\ix_single_ew[35][3] ,
    \ix_single_ew[35][2] ,
    \ix_single_ew[35][1] ,
    \ix_single_ew[35][0] }));
 clb_tile \X[3].Y[5].clb  (.carry_in(\carry[5][3] ),
    .carry_out(\carry[6][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][3] ),
    .set_out_hard(\col_set[6][3] ),
    .shift_in_hard(\col_shift[5][3] ),
    .shift_out_hard(\col_shift[6][3] ),
    .cb_east_in({\dc_ew[44][4] ,
    \dc_ew[44][3] ,
    \dc_ew[44][2] ,
    \dc_ew[44][1] ,
    \dc_ew[44][0] }),
    .cb_east_out({\dc_we[44][9] ,
    \dc_we[44][8] ,
    \dc_we[44][7] ,
    \dc_we[44][6] ,
    \dc_we[44][5] ,
    \dc_we[44][4] ,
    \dc_we[44][3] ,
    \dc_we[44][2] ,
    \dc_we[44][1] ,
    \dc_we[44][0] }),
    .cb_north_in({\dc_ns[45][4] ,
    \dc_ns[45][3] ,
    \dc_ns[45][2] ,
    \dc_ns[45][1] ,
    \dc_ns[45][0] }),
    .cb_north_out({\dc_sn[45][9] ,
    \dc_sn[45][8] ,
    \dc_sn[45][7] ,
    \dc_sn[45][6] ,
    \dc_sn[45][5] ,
    \dc_sn[45][4] ,
    \dc_sn[45][3] ,
    \dc_sn[45][2] ,
    \dc_sn[45][1] ,
    \dc_sn[45][0] }),
    .clb_south_in({\dc_sn[38][9] ,
    \dc_sn[38][8] ,
    \dc_sn[38][7] ,
    \dc_sn[38][6] ,
    \dc_sn[38][5] ,
    \dc_sn[38][4] ,
    \dc_sn[38][3] ,
    \dc_sn[38][2] ,
    \dc_sn[38][1] ,
    \dc_sn[38][0] }),
    .clb_south_out({\dc_ns[38][4] ,
    \dc_ns[38][3] ,
    \dc_ns[38][2] ,
    \dc_ns[38][1] ,
    \dc_ns[38][0] }),
    .clb_west_in({\dc_we[43][9] ,
    \dc_we[43][8] ,
    \dc_we[43][7] ,
    \dc_we[43][6] ,
    \dc_we[43][5] ,
    \dc_we[43][4] ,
    \dc_we[43][3] ,
    \dc_we[43][2] ,
    \dc_we[43][1] ,
    \dc_we[43][0] }),
    .clb_west_out({\dc_ew[43][4] ,
    \dc_ew[43][3] ,
    \dc_ew[43][2] ,
    \dc_ew[43][1] ,
    \dc_ew[43][0] }),
    .east_double({\ix_double_ew[44][7] ,
    \ix_double_ew[44][6] ,
    \ix_double_ew[44][5] ,
    \ix_double_ew[44][4] ,
    \ix_double_ew[44][3] ,
    \ix_double_ew[44][2] ,
    \ix_double_ew[44][1] ,
    \ix_double_ew[44][0] }),
    .east_single({\ix_single_ew[44][3] ,
    \ix_single_ew[44][2] ,
    \ix_single_ew[44][1] ,
    \ix_single_ew[44][0] }),
    .north_double({\ix_double_ns[45][7] ,
    \ix_double_ns[45][6] ,
    \ix_double_ns[45][5] ,
    \ix_double_ns[45][4] ,
    \ix_double_ns[45][3] ,
    \ix_double_ns[45][2] ,
    \ix_double_ns[45][1] ,
    \ix_double_ns[45][0] }),
    .north_single({\ix_single_ns[45][3] ,
    \ix_single_ns[45][2] ,
    \ix_single_ns[45][1] ,
    \ix_single_ns[45][0] }),
    .south_double({\ix_double_ns[38][7] ,
    \ix_double_ns[38][6] ,
    \ix_double_ns[38][5] ,
    \ix_double_ns[38][4] ,
    \ix_double_ns[38][3] ,
    \ix_double_ns[38][2] ,
    \ix_double_ns[38][1] ,
    \ix_double_ns[38][0] }),
    .south_single({\ix_single_ns[38][3] ,
    \ix_single_ns[38][2] ,
    \ix_single_ns[38][1] ,
    \ix_single_ns[38][0] }),
    .west_double({\ix_double_ew[43][7] ,
    \ix_double_ew[43][6] ,
    \ix_double_ew[43][5] ,
    \ix_double_ew[43][4] ,
    \ix_double_ew[43][3] ,
    \ix_double_ew[43][2] ,
    \ix_double_ew[43][1] ,
    \ix_double_ew[43][0] }),
    .west_single({\ix_single_ew[43][3] ,
    \ix_single_ew[43][2] ,
    \ix_single_ew[43][1] ,
    \ix_single_ew[43][0] }));
 clb_tile \X[3].Y[6].clb  (.carry_in(\carry[6][3] ),
    .carry_out(\carry[7][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][3] ),
    .set_out_hard(\col_set[7][3] ),
    .shift_in_hard(\col_shift[6][3] ),
    .shift_out_hard(\col_shift[7][3] ),
    .cb_east_in({\dc_ew[52][4] ,
    \dc_ew[52][3] ,
    \dc_ew[52][2] ,
    \dc_ew[52][1] ,
    \dc_ew[52][0] }),
    .cb_east_out({\dc_we[52][9] ,
    \dc_we[52][8] ,
    \dc_we[52][7] ,
    \dc_we[52][6] ,
    \dc_we[52][5] ,
    \dc_we[52][4] ,
    \dc_we[52][3] ,
    \dc_we[52][2] ,
    \dc_we[52][1] ,
    \dc_we[52][0] }),
    .cb_north_in({\dc_ns[52][4] ,
    \dc_ns[52][3] ,
    \dc_ns[52][2] ,
    \dc_ns[52][1] ,
    \dc_ns[52][0] }),
    .cb_north_out({\dc_sn[52][9] ,
    \dc_sn[52][8] ,
    \dc_sn[52][7] ,
    \dc_sn[52][6] ,
    \dc_sn[52][5] ,
    \dc_sn[52][4] ,
    \dc_sn[52][3] ,
    \dc_sn[52][2] ,
    \dc_sn[52][1] ,
    \dc_sn[52][0] }),
    .clb_south_in({\dc_sn[45][9] ,
    \dc_sn[45][8] ,
    \dc_sn[45][7] ,
    \dc_sn[45][6] ,
    \dc_sn[45][5] ,
    \dc_sn[45][4] ,
    \dc_sn[45][3] ,
    \dc_sn[45][2] ,
    \dc_sn[45][1] ,
    \dc_sn[45][0] }),
    .clb_south_out({\dc_ns[45][4] ,
    \dc_ns[45][3] ,
    \dc_ns[45][2] ,
    \dc_ns[45][1] ,
    \dc_ns[45][0] }),
    .clb_west_in({\dc_we[51][9] ,
    \dc_we[51][8] ,
    \dc_we[51][7] ,
    \dc_we[51][6] ,
    \dc_we[51][5] ,
    \dc_we[51][4] ,
    \dc_we[51][3] ,
    \dc_we[51][2] ,
    \dc_we[51][1] ,
    \dc_we[51][0] }),
    .clb_west_out({\dc_ew[51][4] ,
    \dc_ew[51][3] ,
    \dc_ew[51][2] ,
    \dc_ew[51][1] ,
    \dc_ew[51][0] }),
    .east_double({\ix_double_ew[52][7] ,
    \ix_double_ew[52][6] ,
    \ix_double_ew[52][5] ,
    \ix_double_ew[52][4] ,
    \ix_double_ew[52][3] ,
    \ix_double_ew[52][2] ,
    \ix_double_ew[52][1] ,
    \ix_double_ew[52][0] }),
    .east_single({\ix_single_ew[52][3] ,
    \ix_single_ew[52][2] ,
    \ix_single_ew[52][1] ,
    \ix_single_ew[52][0] }),
    .north_double({\ix_double_ns[52][7] ,
    \ix_double_ns[52][6] ,
    \ix_double_ns[52][5] ,
    \ix_double_ns[52][4] ,
    \ix_double_ns[52][3] ,
    \ix_double_ns[52][2] ,
    \ix_double_ns[52][1] ,
    \ix_double_ns[52][0] }),
    .north_single({\ix_single_ns[52][3] ,
    \ix_single_ns[52][2] ,
    \ix_single_ns[52][1] ,
    \ix_single_ns[52][0] }),
    .south_double({\ix_double_ns[45][7] ,
    \ix_double_ns[45][6] ,
    \ix_double_ns[45][5] ,
    \ix_double_ns[45][4] ,
    \ix_double_ns[45][3] ,
    \ix_double_ns[45][2] ,
    \ix_double_ns[45][1] ,
    \ix_double_ns[45][0] }),
    .south_single({\ix_single_ns[45][3] ,
    \ix_single_ns[45][2] ,
    \ix_single_ns[45][1] ,
    \ix_single_ns[45][0] }),
    .west_double({\ix_double_ew[51][7] ,
    \ix_double_ew[51][6] ,
    \ix_double_ew[51][5] ,
    \ix_double_ew[51][4] ,
    \ix_double_ew[51][3] ,
    \ix_double_ew[51][2] ,
    \ix_double_ew[51][1] ,
    \ix_double_ew[51][0] }),
    .west_single({\ix_single_ew[51][3] ,
    \ix_single_ew[51][2] ,
    \ix_single_ew[51][1] ,
    \ix_single_ew[51][0] }));
 clb_tile \X[3].Y[7].clb  (.carry_in(\carry[7][3] ),
    .carry_out(\carry[8][3] ),
    .cen(\wb_cen_out[0] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][3] ),
    .set_out_hard(\col_set[8][3] ),
    .shift_in_hard(\col_shift[7][3] ),
    .shift_out_hard(\col_shift[8][3] ),
    .cb_east_in({\dc_ew[60][4] ,
    \dc_ew[60][3] ,
    \dc_ew[60][2] ,
    \dc_ew[60][1] ,
    \dc_ew[60][0] }),
    .cb_east_out({\dc_we[60][9] ,
    \dc_we[60][8] ,
    \dc_we[60][7] ,
    \dc_we[60][6] ,
    \dc_we[60][5] ,
    \dc_we[60][4] ,
    \dc_we[60][3] ,
    \dc_we[60][2] ,
    \dc_we[60][1] ,
    \dc_we[60][0] }),
    .cb_north_in({_143_,
    _142_,
    _141_,
    _140_,
    _139_}),
    .cb_north_out({\dc_sn[59][9] ,
    \dc_sn[59][8] ,
    \dc_sn[59][7] ,
    \dc_sn[59][6] ,
    \dc_sn[59][5] ,
    \dc_sn[59][4] ,
    \dc_sn[59][3] ,
    \dc_sn[59][2] ,
    \dc_sn[59][1] ,
    \dc_sn[59][0] }),
    .clb_south_in({\dc_sn[52][9] ,
    \dc_sn[52][8] ,
    \dc_sn[52][7] ,
    \dc_sn[52][6] ,
    \dc_sn[52][5] ,
    \dc_sn[52][4] ,
    \dc_sn[52][3] ,
    \dc_sn[52][2] ,
    \dc_sn[52][1] ,
    \dc_sn[52][0] }),
    .clb_south_out({\dc_ns[52][4] ,
    \dc_ns[52][3] ,
    \dc_ns[52][2] ,
    \dc_ns[52][1] ,
    \dc_ns[52][0] }),
    .clb_west_in({\dc_we[59][9] ,
    \dc_we[59][8] ,
    \dc_we[59][7] ,
    \dc_we[59][6] ,
    \dc_we[59][5] ,
    \dc_we[59][4] ,
    \dc_we[59][3] ,
    \dc_we[59][2] ,
    \dc_we[59][1] ,
    \dc_we[59][0] }),
    .clb_west_out({\dc_ew[59][4] ,
    \dc_ew[59][3] ,
    \dc_ew[59][2] ,
    \dc_ew[59][1] ,
    \dc_ew[59][0] }),
    .east_double({\ix_double_ew[60][7] ,
    \ix_double_ew[60][6] ,
    \ix_double_ew[60][5] ,
    \ix_double_ew[60][4] ,
    \ix_double_ew[60][3] ,
    \ix_double_ew[60][2] ,
    \ix_double_ew[60][1] ,
    \ix_double_ew[60][0] }),
    .east_single({\ix_single_ew[60][3] ,
    \ix_single_ew[60][2] ,
    \ix_single_ew[60][1] ,
    \ix_single_ew[60][0] }),
    .north_double({\ix_double_ns[59][7] ,
    \ix_double_ns[59][6] ,
    \ix_double_ns[59][5] ,
    \ix_double_ns[59][4] ,
    \ix_double_ns[59][3] ,
    \ix_double_ns[59][2] ,
    \ix_double_ns[59][1] ,
    \ix_double_ns[59][0] }),
    .north_single({\ix_single_ns[59][3] ,
    \ix_single_ns[59][2] ,
    \ix_single_ns[59][1] ,
    gpio_north[3]}),
    .south_double({\ix_double_ns[52][7] ,
    \ix_double_ns[52][6] ,
    \ix_double_ns[52][5] ,
    \ix_double_ns[52][4] ,
    \ix_double_ns[52][3] ,
    \ix_double_ns[52][2] ,
    \ix_double_ns[52][1] ,
    \ix_double_ns[52][0] }),
    .south_single({\ix_single_ns[52][3] ,
    \ix_single_ns[52][2] ,
    \ix_single_ns[52][1] ,
    \ix_single_ns[52][0] }),
    .west_double({\ix_double_ew[59][7] ,
    \ix_double_ew[59][6] ,
    \ix_double_ew[59][5] ,
    \ix_double_ew[59][4] ,
    \ix_double_ew[59][3] ,
    \ix_double_ew[59][2] ,
    \ix_double_ew[59][1] ,
    \ix_double_ew[59][0] }),
    .west_single({\ix_single_ew[59][3] ,
    \ix_single_ew[59][2] ,
    \ix_single_ew[59][1] ,
    \ix_single_ew[59][0] }));
 clb_tile \X[4].Y[0].clb  (.carry_in(_144_),
    .carry_out(\carry[1][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[1][0] ),
    .set_out_hard(\col_set[1][4] ),
    .shift_in_hard(\wb_shift_out[1][0] ),
    .shift_out_hard(\col_shift[1][4] ),
    .cb_east_in({\dc_ew[5][4] ,
    \dc_ew[5][3] ,
    \dc_ew[5][2] ,
    \dc_ew[5][1] ,
    \dc_ew[5][0] }),
    .cb_east_out({\dc_we[5][9] ,
    \dc_we[5][8] ,
    \dc_we[5][7] ,
    \dc_we[5][6] ,
    \dc_we[5][5] ,
    \dc_we[5][4] ,
    \dc_we[5][3] ,
    \dc_we[5][2] ,
    \dc_we[5][1] ,
    \dc_we[5][0] }),
    .cb_north_in({\dc_ns[11][4] ,
    \dc_ns[11][3] ,
    \dc_ns[11][2] ,
    \dc_ns[11][1] ,
    \dc_ns[11][0] }),
    .cb_north_out({\dc_sn[11][9] ,
    \dc_sn[11][8] ,
    \dc_sn[11][7] ,
    \dc_sn[11][6] ,
    \dc_sn[11][5] ,
    \dc_sn[11][4] ,
    \dc_sn[11][3] ,
    \dc_sn[11][2] ,
    \dc_sn[11][1] ,
    \dc_sn[11][0] }),
    .clb_south_in({_154_,
    _153_,
    _152_,
    _151_,
    _150_,
    _149_,
    _148_,
    _147_,
    _146_,
    _145_}),
    .clb_south_out({\dc_ns[4][4] ,
    \dc_ns[4][3] ,
    \dc_ns[4][2] ,
    \dc_ns[4][1] ,
    \dc_ns[4][0] }),
    .clb_west_in({\dc_we[4][9] ,
    \dc_we[4][8] ,
    \dc_we[4][7] ,
    \dc_we[4][6] ,
    \dc_we[4][5] ,
    \dc_we[4][4] ,
    \dc_we[4][3] ,
    \dc_we[4][2] ,
    \dc_we[4][1] ,
    \dc_we[4][0] }),
    .clb_west_out({\dc_ew[4][4] ,
    \dc_ew[4][3] ,
    \dc_ew[4][2] ,
    \dc_ew[4][1] ,
    \dc_ew[4][0] }),
    .east_double({\ix_double_ew[5][7] ,
    \ix_double_ew[5][6] ,
    \ix_double_ew[5][5] ,
    \ix_double_ew[5][4] ,
    \ix_double_ew[5][3] ,
    \ix_double_ew[5][2] ,
    \ix_double_ew[5][1] ,
    \ix_double_ew[5][0] }),
    .east_single({\ix_single_ew[5][3] ,
    \ix_single_ew[5][2] ,
    \ix_single_ew[5][1] ,
    \ix_single_ew[5][0] }),
    .north_double({\ix_double_ns[11][7] ,
    \ix_double_ns[11][6] ,
    \ix_double_ns[11][5] ,
    \ix_double_ns[11][4] ,
    \ix_double_ns[11][3] ,
    \ix_double_ns[11][2] ,
    \ix_double_ns[11][1] ,
    \ix_double_ns[11][0] }),
    .north_single({\ix_single_ns[11][3] ,
    \ix_single_ns[11][2] ,
    \ix_single_ns[11][1] ,
    \ix_single_ns[11][0] }),
    .south_double({\ix_double_ns[4][7] ,
    \ix_double_ns[4][6] ,
    \ix_double_ns[4][5] ,
    \ix_double_ns[4][4] ,
    \ix_double_ns[4][3] ,
    \ix_double_ns[4][2] ,
    \ix_double_ns[4][1] ,
    \ix_double_ns[4][0] }),
    .south_single({\ix_single_ns[4][3] ,
    \ix_single_ns[4][2] ,
    \ix_single_ns[4][1] ,
    gpio_south[4]}),
    .west_double({\ix_double_ew[4][7] ,
    \ix_double_ew[4][6] ,
    \ix_double_ew[4][5] ,
    \ix_double_ew[4][4] ,
    \ix_double_ew[4][3] ,
    \ix_double_ew[4][2] ,
    \ix_double_ew[4][1] ,
    \ix_double_ew[4][0] }),
    .west_single({\ix_single_ew[4][3] ,
    \ix_single_ew[4][2] ,
    \ix_single_ew[4][1] ,
    \ix_single_ew[4][0] }));
 clb_tile \X[4].Y[1].clb  (.carry_in(\carry[1][4] ),
    .carry_out(\carry[2][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][4] ),
    .set_out_hard(\col_set[2][4] ),
    .shift_in_hard(\col_shift[1][4] ),
    .shift_out_hard(\col_shift[2][4] ),
    .cb_east_in({\dc_ew[13][4] ,
    \dc_ew[13][3] ,
    \dc_ew[13][2] ,
    \dc_ew[13][1] ,
    \dc_ew[13][0] }),
    .cb_east_out({\dc_we[13][9] ,
    \dc_we[13][8] ,
    \dc_we[13][7] ,
    \dc_we[13][6] ,
    \dc_we[13][5] ,
    \dc_we[13][4] ,
    \dc_we[13][3] ,
    \dc_we[13][2] ,
    \dc_we[13][1] ,
    \dc_we[13][0] }),
    .cb_north_in({\dc_ns[18][4] ,
    \dc_ns[18][3] ,
    \dc_ns[18][2] ,
    \dc_ns[18][1] ,
    \dc_ns[18][0] }),
    .cb_north_out({\dc_sn[18][9] ,
    \dc_sn[18][8] ,
    \dc_sn[18][7] ,
    \dc_sn[18][6] ,
    \dc_sn[18][5] ,
    \dc_sn[18][4] ,
    \dc_sn[18][3] ,
    \dc_sn[18][2] ,
    \dc_sn[18][1] ,
    \dc_sn[18][0] }),
    .clb_south_in({\dc_sn[11][9] ,
    \dc_sn[11][8] ,
    \dc_sn[11][7] ,
    \dc_sn[11][6] ,
    \dc_sn[11][5] ,
    \dc_sn[11][4] ,
    \dc_sn[11][3] ,
    \dc_sn[11][2] ,
    \dc_sn[11][1] ,
    \dc_sn[11][0] }),
    .clb_south_out({\dc_ns[11][4] ,
    \dc_ns[11][3] ,
    \dc_ns[11][2] ,
    \dc_ns[11][1] ,
    \dc_ns[11][0] }),
    .clb_west_in({\dc_we[12][9] ,
    \dc_we[12][8] ,
    \dc_we[12][7] ,
    \dc_we[12][6] ,
    \dc_we[12][5] ,
    \dc_we[12][4] ,
    \dc_we[12][3] ,
    \dc_we[12][2] ,
    \dc_we[12][1] ,
    \dc_we[12][0] }),
    .clb_west_out({\dc_ew[12][4] ,
    \dc_ew[12][3] ,
    \dc_ew[12][2] ,
    \dc_ew[12][1] ,
    \dc_ew[12][0] }),
    .east_double({\ix_double_ew[13][7] ,
    \ix_double_ew[13][6] ,
    \ix_double_ew[13][5] ,
    \ix_double_ew[13][4] ,
    \ix_double_ew[13][3] ,
    \ix_double_ew[13][2] ,
    \ix_double_ew[13][1] ,
    \ix_double_ew[13][0] }),
    .east_single({\ix_single_ew[13][3] ,
    \ix_single_ew[13][2] ,
    \ix_single_ew[13][1] ,
    \ix_single_ew[13][0] }),
    .north_double({\ix_double_ns[18][7] ,
    \ix_double_ns[18][6] ,
    \ix_double_ns[18][5] ,
    \ix_double_ns[18][4] ,
    \ix_double_ns[18][3] ,
    \ix_double_ns[18][2] ,
    \ix_double_ns[18][1] ,
    \ix_double_ns[18][0] }),
    .north_single({\ix_single_ns[18][3] ,
    \ix_single_ns[18][2] ,
    \ix_single_ns[18][1] ,
    \ix_single_ns[18][0] }),
    .south_double({\ix_double_ns[11][7] ,
    \ix_double_ns[11][6] ,
    \ix_double_ns[11][5] ,
    \ix_double_ns[11][4] ,
    \ix_double_ns[11][3] ,
    \ix_double_ns[11][2] ,
    \ix_double_ns[11][1] ,
    \ix_double_ns[11][0] }),
    .south_single({\ix_single_ns[11][3] ,
    \ix_single_ns[11][2] ,
    \ix_single_ns[11][1] ,
    \ix_single_ns[11][0] }),
    .west_double({\ix_double_ew[12][7] ,
    \ix_double_ew[12][6] ,
    \ix_double_ew[12][5] ,
    \ix_double_ew[12][4] ,
    \ix_double_ew[12][3] ,
    \ix_double_ew[12][2] ,
    \ix_double_ew[12][1] ,
    \ix_double_ew[12][0] }),
    .west_single({\ix_single_ew[12][3] ,
    \ix_single_ew[12][2] ,
    \ix_single_ew[12][1] ,
    \ix_single_ew[12][0] }));
 clb_tile \X[4].Y[2].clb  (.carry_in(\carry[2][4] ),
    .carry_out(\carry[3][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][4] ),
    .set_out_hard(\col_set[3][4] ),
    .shift_in_hard(\col_shift[2][4] ),
    .shift_out_hard(\col_shift[3][4] ),
    .cb_east_in({\dc_ew[21][4] ,
    \dc_ew[21][3] ,
    \dc_ew[21][2] ,
    \dc_ew[21][1] ,
    \dc_ew[21][0] }),
    .cb_east_out({\dc_we[21][9] ,
    \dc_we[21][8] ,
    \dc_we[21][7] ,
    \dc_we[21][6] ,
    \dc_we[21][5] ,
    \dc_we[21][4] ,
    \dc_we[21][3] ,
    \dc_we[21][2] ,
    \dc_we[21][1] ,
    \dc_we[21][0] }),
    .cb_north_in({\dc_ns[25][4] ,
    \dc_ns[25][3] ,
    \dc_ns[25][2] ,
    \dc_ns[25][1] ,
    \dc_ns[25][0] }),
    .cb_north_out({\dc_sn[25][9] ,
    \dc_sn[25][8] ,
    \dc_sn[25][7] ,
    \dc_sn[25][6] ,
    \dc_sn[25][5] ,
    \dc_sn[25][4] ,
    \dc_sn[25][3] ,
    \dc_sn[25][2] ,
    \dc_sn[25][1] ,
    \dc_sn[25][0] }),
    .clb_south_in({\dc_sn[18][9] ,
    \dc_sn[18][8] ,
    \dc_sn[18][7] ,
    \dc_sn[18][6] ,
    \dc_sn[18][5] ,
    \dc_sn[18][4] ,
    \dc_sn[18][3] ,
    \dc_sn[18][2] ,
    \dc_sn[18][1] ,
    \dc_sn[18][0] }),
    .clb_south_out({\dc_ns[18][4] ,
    \dc_ns[18][3] ,
    \dc_ns[18][2] ,
    \dc_ns[18][1] ,
    \dc_ns[18][0] }),
    .clb_west_in({\dc_we[20][9] ,
    \dc_we[20][8] ,
    \dc_we[20][7] ,
    \dc_we[20][6] ,
    \dc_we[20][5] ,
    \dc_we[20][4] ,
    \dc_we[20][3] ,
    \dc_we[20][2] ,
    \dc_we[20][1] ,
    \dc_we[20][0] }),
    .clb_west_out({\dc_ew[20][4] ,
    \dc_ew[20][3] ,
    \dc_ew[20][2] ,
    \dc_ew[20][1] ,
    \dc_ew[20][0] }),
    .east_double({\ix_double_ew[21][7] ,
    \ix_double_ew[21][6] ,
    \ix_double_ew[21][5] ,
    \ix_double_ew[21][4] ,
    \ix_double_ew[21][3] ,
    \ix_double_ew[21][2] ,
    \ix_double_ew[21][1] ,
    \ix_double_ew[21][0] }),
    .east_single({\ix_single_ew[21][3] ,
    \ix_single_ew[21][2] ,
    \ix_single_ew[21][1] ,
    \ix_single_ew[21][0] }),
    .north_double({\ix_double_ns[25][7] ,
    \ix_double_ns[25][6] ,
    \ix_double_ns[25][5] ,
    \ix_double_ns[25][4] ,
    \ix_double_ns[25][3] ,
    \ix_double_ns[25][2] ,
    \ix_double_ns[25][1] ,
    \ix_double_ns[25][0] }),
    .north_single({\ix_single_ns[25][3] ,
    \ix_single_ns[25][2] ,
    \ix_single_ns[25][1] ,
    \ix_single_ns[25][0] }),
    .south_double({\ix_double_ns[18][7] ,
    \ix_double_ns[18][6] ,
    \ix_double_ns[18][5] ,
    \ix_double_ns[18][4] ,
    \ix_double_ns[18][3] ,
    \ix_double_ns[18][2] ,
    \ix_double_ns[18][1] ,
    \ix_double_ns[18][0] }),
    .south_single({\ix_single_ns[18][3] ,
    \ix_single_ns[18][2] ,
    \ix_single_ns[18][1] ,
    \ix_single_ns[18][0] }),
    .west_double({\ix_double_ew[20][7] ,
    \ix_double_ew[20][6] ,
    \ix_double_ew[20][5] ,
    \ix_double_ew[20][4] ,
    \ix_double_ew[20][3] ,
    \ix_double_ew[20][2] ,
    \ix_double_ew[20][1] ,
    \ix_double_ew[20][0] }),
    .west_single({\ix_single_ew[20][3] ,
    \ix_single_ew[20][2] ,
    \ix_single_ew[20][1] ,
    \ix_single_ew[20][0] }));
 clb_tile \X[4].Y[3].clb  (.carry_in(\carry[3][4] ),
    .carry_out(\carry[4][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][4] ),
    .set_out_hard(\col_set[4][4] ),
    .shift_in_hard(\col_shift[3][4] ),
    .shift_out_hard(\col_shift[4][4] ),
    .cb_east_in({\dc_ew[29][4] ,
    \dc_ew[29][3] ,
    \dc_ew[29][2] ,
    \dc_ew[29][1] ,
    \dc_ew[29][0] }),
    .cb_east_out({\dc_we[29][9] ,
    \dc_we[29][8] ,
    \dc_we[29][7] ,
    \dc_we[29][6] ,
    \dc_we[29][5] ,
    \dc_we[29][4] ,
    \dc_we[29][3] ,
    \dc_we[29][2] ,
    \dc_we[29][1] ,
    \dc_we[29][0] }),
    .cb_north_in({\dc_ns[32][4] ,
    \dc_ns[32][3] ,
    \dc_ns[32][2] ,
    \dc_ns[32][1] ,
    \dc_ns[32][0] }),
    .cb_north_out({\dc_sn[32][9] ,
    \dc_sn[32][8] ,
    \dc_sn[32][7] ,
    \dc_sn[32][6] ,
    \dc_sn[32][5] ,
    \dc_sn[32][4] ,
    \dc_sn[32][3] ,
    \dc_sn[32][2] ,
    \dc_sn[32][1] ,
    \dc_sn[32][0] }),
    .clb_south_in({\dc_sn[25][9] ,
    \dc_sn[25][8] ,
    \dc_sn[25][7] ,
    \dc_sn[25][6] ,
    \dc_sn[25][5] ,
    \dc_sn[25][4] ,
    \dc_sn[25][3] ,
    \dc_sn[25][2] ,
    \dc_sn[25][1] ,
    \dc_sn[25][0] }),
    .clb_south_out({\dc_ns[25][4] ,
    \dc_ns[25][3] ,
    \dc_ns[25][2] ,
    \dc_ns[25][1] ,
    \dc_ns[25][0] }),
    .clb_west_in({\dc_we[28][9] ,
    \dc_we[28][8] ,
    \dc_we[28][7] ,
    \dc_we[28][6] ,
    \dc_we[28][5] ,
    \dc_we[28][4] ,
    \dc_we[28][3] ,
    \dc_we[28][2] ,
    \dc_we[28][1] ,
    \dc_we[28][0] }),
    .clb_west_out({\dc_ew[28][4] ,
    \dc_ew[28][3] ,
    \dc_ew[28][2] ,
    \dc_ew[28][1] ,
    \dc_ew[28][0] }),
    .east_double({\ix_double_ew[29][7] ,
    \ix_double_ew[29][6] ,
    \ix_double_ew[29][5] ,
    \ix_double_ew[29][4] ,
    \ix_double_ew[29][3] ,
    \ix_double_ew[29][2] ,
    \ix_double_ew[29][1] ,
    \ix_double_ew[29][0] }),
    .east_single({\ix_single_ew[29][3] ,
    \ix_single_ew[29][2] ,
    \ix_single_ew[29][1] ,
    \ix_single_ew[29][0] }),
    .north_double({\ix_double_ns[32][7] ,
    \ix_double_ns[32][6] ,
    \ix_double_ns[32][5] ,
    \ix_double_ns[32][4] ,
    \ix_double_ns[32][3] ,
    \ix_double_ns[32][2] ,
    \ix_double_ns[32][1] ,
    \ix_double_ns[32][0] }),
    .north_single({\ix_single_ns[32][3] ,
    \ix_single_ns[32][2] ,
    \ix_single_ns[32][1] ,
    \ix_single_ns[32][0] }),
    .south_double({\ix_double_ns[25][7] ,
    \ix_double_ns[25][6] ,
    \ix_double_ns[25][5] ,
    \ix_double_ns[25][4] ,
    \ix_double_ns[25][3] ,
    \ix_double_ns[25][2] ,
    \ix_double_ns[25][1] ,
    \ix_double_ns[25][0] }),
    .south_single({\ix_single_ns[25][3] ,
    \ix_single_ns[25][2] ,
    \ix_single_ns[25][1] ,
    \ix_single_ns[25][0] }),
    .west_double({\ix_double_ew[28][7] ,
    \ix_double_ew[28][6] ,
    \ix_double_ew[28][5] ,
    \ix_double_ew[28][4] ,
    \ix_double_ew[28][3] ,
    \ix_double_ew[28][2] ,
    \ix_double_ew[28][1] ,
    \ix_double_ew[28][0] }),
    .west_single({\ix_single_ew[28][3] ,
    \ix_single_ew[28][2] ,
    \ix_single_ew[28][1] ,
    \ix_single_ew[28][0] }));
 clb_tile \X[4].Y[4].clb  (.carry_in(\carry[4][4] ),
    .carry_out(\carry[5][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][4] ),
    .set_out_hard(\col_set[5][4] ),
    .shift_in_hard(\col_shift[4][4] ),
    .shift_out_hard(\col_shift[5][4] ),
    .cb_east_in({\dc_ew[37][4] ,
    \dc_ew[37][3] ,
    \dc_ew[37][2] ,
    \dc_ew[37][1] ,
    \dc_ew[37][0] }),
    .cb_east_out({\dc_we[37][9] ,
    \dc_we[37][8] ,
    \dc_we[37][7] ,
    \dc_we[37][6] ,
    \dc_we[37][5] ,
    \dc_we[37][4] ,
    \dc_we[37][3] ,
    \dc_we[37][2] ,
    \dc_we[37][1] ,
    \dc_we[37][0] }),
    .cb_north_in({\dc_ns[39][4] ,
    \dc_ns[39][3] ,
    \dc_ns[39][2] ,
    \dc_ns[39][1] ,
    \dc_ns[39][0] }),
    .cb_north_out({\dc_sn[39][9] ,
    \dc_sn[39][8] ,
    \dc_sn[39][7] ,
    \dc_sn[39][6] ,
    \dc_sn[39][5] ,
    \dc_sn[39][4] ,
    \dc_sn[39][3] ,
    \dc_sn[39][2] ,
    \dc_sn[39][1] ,
    \dc_sn[39][0] }),
    .clb_south_in({\dc_sn[32][9] ,
    \dc_sn[32][8] ,
    \dc_sn[32][7] ,
    \dc_sn[32][6] ,
    \dc_sn[32][5] ,
    \dc_sn[32][4] ,
    \dc_sn[32][3] ,
    \dc_sn[32][2] ,
    \dc_sn[32][1] ,
    \dc_sn[32][0] }),
    .clb_south_out({\dc_ns[32][4] ,
    \dc_ns[32][3] ,
    \dc_ns[32][2] ,
    \dc_ns[32][1] ,
    \dc_ns[32][0] }),
    .clb_west_in({\dc_we[36][9] ,
    \dc_we[36][8] ,
    \dc_we[36][7] ,
    \dc_we[36][6] ,
    \dc_we[36][5] ,
    \dc_we[36][4] ,
    \dc_we[36][3] ,
    \dc_we[36][2] ,
    \dc_we[36][1] ,
    \dc_we[36][0] }),
    .clb_west_out({\dc_ew[36][4] ,
    \dc_ew[36][3] ,
    \dc_ew[36][2] ,
    \dc_ew[36][1] ,
    \dc_ew[36][0] }),
    .east_double({\ix_double_ew[37][7] ,
    \ix_double_ew[37][6] ,
    \ix_double_ew[37][5] ,
    \ix_double_ew[37][4] ,
    \ix_double_ew[37][3] ,
    \ix_double_ew[37][2] ,
    \ix_double_ew[37][1] ,
    \ix_double_ew[37][0] }),
    .east_single({\ix_single_ew[37][3] ,
    \ix_single_ew[37][2] ,
    \ix_single_ew[37][1] ,
    \ix_single_ew[37][0] }),
    .north_double({\ix_double_ns[39][7] ,
    \ix_double_ns[39][6] ,
    \ix_double_ns[39][5] ,
    \ix_double_ns[39][4] ,
    \ix_double_ns[39][3] ,
    \ix_double_ns[39][2] ,
    \ix_double_ns[39][1] ,
    \ix_double_ns[39][0] }),
    .north_single({\ix_single_ns[39][3] ,
    \ix_single_ns[39][2] ,
    \ix_single_ns[39][1] ,
    \ix_single_ns[39][0] }),
    .south_double({\ix_double_ns[32][7] ,
    \ix_double_ns[32][6] ,
    \ix_double_ns[32][5] ,
    \ix_double_ns[32][4] ,
    \ix_double_ns[32][3] ,
    \ix_double_ns[32][2] ,
    \ix_double_ns[32][1] ,
    \ix_double_ns[32][0] }),
    .south_single({\ix_single_ns[32][3] ,
    \ix_single_ns[32][2] ,
    \ix_single_ns[32][1] ,
    \ix_single_ns[32][0] }),
    .west_double({\ix_double_ew[36][7] ,
    \ix_double_ew[36][6] ,
    \ix_double_ew[36][5] ,
    \ix_double_ew[36][4] ,
    \ix_double_ew[36][3] ,
    \ix_double_ew[36][2] ,
    \ix_double_ew[36][1] ,
    \ix_double_ew[36][0] }),
    .west_single({\ix_single_ew[36][3] ,
    \ix_single_ew[36][2] ,
    \ix_single_ew[36][1] ,
    \ix_single_ew[36][0] }));
 clb_tile \X[4].Y[5].clb  (.carry_in(\carry[5][4] ),
    .carry_out(\carry[6][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][4] ),
    .set_out_hard(\col_set[6][4] ),
    .shift_in_hard(\col_shift[5][4] ),
    .shift_out_hard(\col_shift[6][4] ),
    .cb_east_in({\dc_ew[45][4] ,
    \dc_ew[45][3] ,
    \dc_ew[45][2] ,
    \dc_ew[45][1] ,
    \dc_ew[45][0] }),
    .cb_east_out({\dc_we[45][9] ,
    \dc_we[45][8] ,
    \dc_we[45][7] ,
    \dc_we[45][6] ,
    \dc_we[45][5] ,
    \dc_we[45][4] ,
    \dc_we[45][3] ,
    \dc_we[45][2] ,
    \dc_we[45][1] ,
    \dc_we[45][0] }),
    .cb_north_in({\dc_ns[46][4] ,
    \dc_ns[46][3] ,
    \dc_ns[46][2] ,
    \dc_ns[46][1] ,
    \dc_ns[46][0] }),
    .cb_north_out({\dc_sn[46][9] ,
    \dc_sn[46][8] ,
    \dc_sn[46][7] ,
    \dc_sn[46][6] ,
    \dc_sn[46][5] ,
    \dc_sn[46][4] ,
    \dc_sn[46][3] ,
    \dc_sn[46][2] ,
    \dc_sn[46][1] ,
    \dc_sn[46][0] }),
    .clb_south_in({\dc_sn[39][9] ,
    \dc_sn[39][8] ,
    \dc_sn[39][7] ,
    \dc_sn[39][6] ,
    \dc_sn[39][5] ,
    \dc_sn[39][4] ,
    \dc_sn[39][3] ,
    \dc_sn[39][2] ,
    \dc_sn[39][1] ,
    \dc_sn[39][0] }),
    .clb_south_out({\dc_ns[39][4] ,
    \dc_ns[39][3] ,
    \dc_ns[39][2] ,
    \dc_ns[39][1] ,
    \dc_ns[39][0] }),
    .clb_west_in({\dc_we[44][9] ,
    \dc_we[44][8] ,
    \dc_we[44][7] ,
    \dc_we[44][6] ,
    \dc_we[44][5] ,
    \dc_we[44][4] ,
    \dc_we[44][3] ,
    \dc_we[44][2] ,
    \dc_we[44][1] ,
    \dc_we[44][0] }),
    .clb_west_out({\dc_ew[44][4] ,
    \dc_ew[44][3] ,
    \dc_ew[44][2] ,
    \dc_ew[44][1] ,
    \dc_ew[44][0] }),
    .east_double({\ix_double_ew[45][7] ,
    \ix_double_ew[45][6] ,
    \ix_double_ew[45][5] ,
    \ix_double_ew[45][4] ,
    \ix_double_ew[45][3] ,
    \ix_double_ew[45][2] ,
    \ix_double_ew[45][1] ,
    \ix_double_ew[45][0] }),
    .east_single({\ix_single_ew[45][3] ,
    \ix_single_ew[45][2] ,
    \ix_single_ew[45][1] ,
    \ix_single_ew[45][0] }),
    .north_double({\ix_double_ns[46][7] ,
    \ix_double_ns[46][6] ,
    \ix_double_ns[46][5] ,
    \ix_double_ns[46][4] ,
    \ix_double_ns[46][3] ,
    \ix_double_ns[46][2] ,
    \ix_double_ns[46][1] ,
    \ix_double_ns[46][0] }),
    .north_single({\ix_single_ns[46][3] ,
    \ix_single_ns[46][2] ,
    \ix_single_ns[46][1] ,
    \ix_single_ns[46][0] }),
    .south_double({\ix_double_ns[39][7] ,
    \ix_double_ns[39][6] ,
    \ix_double_ns[39][5] ,
    \ix_double_ns[39][4] ,
    \ix_double_ns[39][3] ,
    \ix_double_ns[39][2] ,
    \ix_double_ns[39][1] ,
    \ix_double_ns[39][0] }),
    .south_single({\ix_single_ns[39][3] ,
    \ix_single_ns[39][2] ,
    \ix_single_ns[39][1] ,
    \ix_single_ns[39][0] }),
    .west_double({\ix_double_ew[44][7] ,
    \ix_double_ew[44][6] ,
    \ix_double_ew[44][5] ,
    \ix_double_ew[44][4] ,
    \ix_double_ew[44][3] ,
    \ix_double_ew[44][2] ,
    \ix_double_ew[44][1] ,
    \ix_double_ew[44][0] }),
    .west_single({\ix_single_ew[44][3] ,
    \ix_single_ew[44][2] ,
    \ix_single_ew[44][1] ,
    \ix_single_ew[44][0] }));
 clb_tile \X[4].Y[6].clb  (.carry_in(\carry[6][4] ),
    .carry_out(\carry[7][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][4] ),
    .set_out_hard(\col_set[7][4] ),
    .shift_in_hard(\col_shift[6][4] ),
    .shift_out_hard(\col_shift[7][4] ),
    .cb_east_in({\dc_ew[53][4] ,
    \dc_ew[53][3] ,
    \dc_ew[53][2] ,
    \dc_ew[53][1] ,
    \dc_ew[53][0] }),
    .cb_east_out({\dc_we[53][9] ,
    \dc_we[53][8] ,
    \dc_we[53][7] ,
    \dc_we[53][6] ,
    \dc_we[53][5] ,
    \dc_we[53][4] ,
    \dc_we[53][3] ,
    \dc_we[53][2] ,
    \dc_we[53][1] ,
    \dc_we[53][0] }),
    .cb_north_in({\dc_ns[53][4] ,
    \dc_ns[53][3] ,
    \dc_ns[53][2] ,
    \dc_ns[53][1] ,
    \dc_ns[53][0] }),
    .cb_north_out({\dc_sn[53][9] ,
    \dc_sn[53][8] ,
    \dc_sn[53][7] ,
    \dc_sn[53][6] ,
    \dc_sn[53][5] ,
    \dc_sn[53][4] ,
    \dc_sn[53][3] ,
    \dc_sn[53][2] ,
    \dc_sn[53][1] ,
    \dc_sn[53][0] }),
    .clb_south_in({\dc_sn[46][9] ,
    \dc_sn[46][8] ,
    \dc_sn[46][7] ,
    \dc_sn[46][6] ,
    \dc_sn[46][5] ,
    \dc_sn[46][4] ,
    \dc_sn[46][3] ,
    \dc_sn[46][2] ,
    \dc_sn[46][1] ,
    \dc_sn[46][0] }),
    .clb_south_out({\dc_ns[46][4] ,
    \dc_ns[46][3] ,
    \dc_ns[46][2] ,
    \dc_ns[46][1] ,
    \dc_ns[46][0] }),
    .clb_west_in({\dc_we[52][9] ,
    \dc_we[52][8] ,
    \dc_we[52][7] ,
    \dc_we[52][6] ,
    \dc_we[52][5] ,
    \dc_we[52][4] ,
    \dc_we[52][3] ,
    \dc_we[52][2] ,
    \dc_we[52][1] ,
    \dc_we[52][0] }),
    .clb_west_out({\dc_ew[52][4] ,
    \dc_ew[52][3] ,
    \dc_ew[52][2] ,
    \dc_ew[52][1] ,
    \dc_ew[52][0] }),
    .east_double({\ix_double_ew[53][7] ,
    \ix_double_ew[53][6] ,
    \ix_double_ew[53][5] ,
    \ix_double_ew[53][4] ,
    \ix_double_ew[53][3] ,
    \ix_double_ew[53][2] ,
    \ix_double_ew[53][1] ,
    \ix_double_ew[53][0] }),
    .east_single({\ix_single_ew[53][3] ,
    \ix_single_ew[53][2] ,
    \ix_single_ew[53][1] ,
    \ix_single_ew[53][0] }),
    .north_double({\ix_double_ns[53][7] ,
    \ix_double_ns[53][6] ,
    \ix_double_ns[53][5] ,
    \ix_double_ns[53][4] ,
    \ix_double_ns[53][3] ,
    \ix_double_ns[53][2] ,
    \ix_double_ns[53][1] ,
    \ix_double_ns[53][0] }),
    .north_single({\ix_single_ns[53][3] ,
    \ix_single_ns[53][2] ,
    \ix_single_ns[53][1] ,
    \ix_single_ns[53][0] }),
    .south_double({\ix_double_ns[46][7] ,
    \ix_double_ns[46][6] ,
    \ix_double_ns[46][5] ,
    \ix_double_ns[46][4] ,
    \ix_double_ns[46][3] ,
    \ix_double_ns[46][2] ,
    \ix_double_ns[46][1] ,
    \ix_double_ns[46][0] }),
    .south_single({\ix_single_ns[46][3] ,
    \ix_single_ns[46][2] ,
    \ix_single_ns[46][1] ,
    \ix_single_ns[46][0] }),
    .west_double({\ix_double_ew[52][7] ,
    \ix_double_ew[52][6] ,
    \ix_double_ew[52][5] ,
    \ix_double_ew[52][4] ,
    \ix_double_ew[52][3] ,
    \ix_double_ew[52][2] ,
    \ix_double_ew[52][1] ,
    \ix_double_ew[52][0] }),
    .west_single({\ix_single_ew[52][3] ,
    \ix_single_ew[52][2] ,
    \ix_single_ew[52][1] ,
    \ix_single_ew[52][0] }));
 clb_tile \X[4].Y[7].clb  (.carry_in(\carry[7][4] ),
    .carry_out(\carry[8][4] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][4] ),
    .set_out_hard(\col_set[8][4] ),
    .shift_in_hard(\col_shift[7][4] ),
    .shift_out_hard(\col_shift[8][4] ),
    .cb_east_in({\dc_ew[61][4] ,
    \dc_ew[61][3] ,
    \dc_ew[61][2] ,
    \dc_ew[61][1] ,
    \dc_ew[61][0] }),
    .cb_east_out({\dc_we[61][9] ,
    \dc_we[61][8] ,
    \dc_we[61][7] ,
    \dc_we[61][6] ,
    \dc_we[61][5] ,
    \dc_we[61][4] ,
    \dc_we[61][3] ,
    \dc_we[61][2] ,
    \dc_we[61][1] ,
    \dc_we[61][0] }),
    .cb_north_in({_159_,
    _158_,
    _157_,
    _156_,
    _155_}),
    .cb_north_out({\dc_sn[60][9] ,
    \dc_sn[60][8] ,
    \dc_sn[60][7] ,
    \dc_sn[60][6] ,
    \dc_sn[60][5] ,
    \dc_sn[60][4] ,
    \dc_sn[60][3] ,
    \dc_sn[60][2] ,
    \dc_sn[60][1] ,
    \dc_sn[60][0] }),
    .clb_south_in({\dc_sn[53][9] ,
    \dc_sn[53][8] ,
    \dc_sn[53][7] ,
    \dc_sn[53][6] ,
    \dc_sn[53][5] ,
    \dc_sn[53][4] ,
    \dc_sn[53][3] ,
    \dc_sn[53][2] ,
    \dc_sn[53][1] ,
    \dc_sn[53][0] }),
    .clb_south_out({\dc_ns[53][4] ,
    \dc_ns[53][3] ,
    \dc_ns[53][2] ,
    \dc_ns[53][1] ,
    \dc_ns[53][0] }),
    .clb_west_in({\dc_we[60][9] ,
    \dc_we[60][8] ,
    \dc_we[60][7] ,
    \dc_we[60][6] ,
    \dc_we[60][5] ,
    \dc_we[60][4] ,
    \dc_we[60][3] ,
    \dc_we[60][2] ,
    \dc_we[60][1] ,
    \dc_we[60][0] }),
    .clb_west_out({\dc_ew[60][4] ,
    \dc_ew[60][3] ,
    \dc_ew[60][2] ,
    \dc_ew[60][1] ,
    \dc_ew[60][0] }),
    .east_double({\ix_double_ew[61][7] ,
    \ix_double_ew[61][6] ,
    \ix_double_ew[61][5] ,
    \ix_double_ew[61][4] ,
    \ix_double_ew[61][3] ,
    \ix_double_ew[61][2] ,
    \ix_double_ew[61][1] ,
    \ix_double_ew[61][0] }),
    .east_single({\ix_single_ew[61][3] ,
    \ix_single_ew[61][2] ,
    \ix_single_ew[61][1] ,
    \ix_single_ew[61][0] }),
    .north_double({\ix_double_ns[60][7] ,
    \ix_double_ns[60][6] ,
    \ix_double_ns[60][5] ,
    \ix_double_ns[60][4] ,
    \ix_double_ns[60][3] ,
    \ix_double_ns[60][2] ,
    \ix_double_ns[60][1] ,
    \ix_double_ns[60][0] }),
    .north_single({\ix_single_ns[60][3] ,
    \ix_single_ns[60][2] ,
    \ix_single_ns[60][1] ,
    gpio_north[4]}),
    .south_double({\ix_double_ns[53][7] ,
    \ix_double_ns[53][6] ,
    \ix_double_ns[53][5] ,
    \ix_double_ns[53][4] ,
    \ix_double_ns[53][3] ,
    \ix_double_ns[53][2] ,
    \ix_double_ns[53][1] ,
    \ix_double_ns[53][0] }),
    .south_single({\ix_single_ns[53][3] ,
    \ix_single_ns[53][2] ,
    \ix_single_ns[53][1] ,
    \ix_single_ns[53][0] }),
    .west_double({\ix_double_ew[60][7] ,
    \ix_double_ew[60][6] ,
    \ix_double_ew[60][5] ,
    \ix_double_ew[60][4] ,
    \ix_double_ew[60][3] ,
    \ix_double_ew[60][2] ,
    \ix_double_ew[60][1] ,
    \ix_double_ew[60][0] }),
    .west_single({\ix_single_ew[60][3] ,
    \ix_single_ew[60][2] ,
    \ix_single_ew[60][1] ,
    \ix_single_ew[60][0] }));
 clb_tile \X[5].Y[0].clb  (.carry_in(_160_),
    .carry_out(\carry[1][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[1][1] ),
    .set_out_hard(\col_set[1][5] ),
    .shift_in_hard(\wb_shift_out[1][1] ),
    .shift_out_hard(\col_shift[1][5] ),
    .cb_east_in({\dc_ew[6][4] ,
    \dc_ew[6][3] ,
    \dc_ew[6][2] ,
    \dc_ew[6][1] ,
    \dc_ew[6][0] }),
    .cb_east_out({\dc_we[6][9] ,
    \dc_we[6][8] ,
    \dc_we[6][7] ,
    \dc_we[6][6] ,
    \dc_we[6][5] ,
    \dc_we[6][4] ,
    \dc_we[6][3] ,
    \dc_we[6][2] ,
    \dc_we[6][1] ,
    \dc_we[6][0] }),
    .cb_north_in({\dc_ns[12][4] ,
    \dc_ns[12][3] ,
    \dc_ns[12][2] ,
    \dc_ns[12][1] ,
    \dc_ns[12][0] }),
    .cb_north_out({\dc_sn[12][9] ,
    \dc_sn[12][8] ,
    \dc_sn[12][7] ,
    \dc_sn[12][6] ,
    \dc_sn[12][5] ,
    \dc_sn[12][4] ,
    \dc_sn[12][3] ,
    \dc_sn[12][2] ,
    \dc_sn[12][1] ,
    \dc_sn[12][0] }),
    .clb_south_in({_170_,
    _169_,
    _168_,
    _167_,
    _166_,
    _165_,
    _164_,
    _163_,
    _162_,
    _161_}),
    .clb_south_out({\dc_ns[5][4] ,
    \dc_ns[5][3] ,
    \dc_ns[5][2] ,
    \dc_ns[5][1] ,
    \dc_ns[5][0] }),
    .clb_west_in({\dc_we[5][9] ,
    \dc_we[5][8] ,
    \dc_we[5][7] ,
    \dc_we[5][6] ,
    \dc_we[5][5] ,
    \dc_we[5][4] ,
    \dc_we[5][3] ,
    \dc_we[5][2] ,
    \dc_we[5][1] ,
    \dc_we[5][0] }),
    .clb_west_out({\dc_ew[5][4] ,
    \dc_ew[5][3] ,
    \dc_ew[5][2] ,
    \dc_ew[5][1] ,
    \dc_ew[5][0] }),
    .east_double({\ix_double_ew[6][7] ,
    \ix_double_ew[6][6] ,
    \ix_double_ew[6][5] ,
    \ix_double_ew[6][4] ,
    \ix_double_ew[6][3] ,
    \ix_double_ew[6][2] ,
    \ix_double_ew[6][1] ,
    \ix_double_ew[6][0] }),
    .east_single({\ix_single_ew[6][3] ,
    \ix_single_ew[6][2] ,
    \ix_single_ew[6][1] ,
    \ix_single_ew[6][0] }),
    .north_double({\ix_double_ns[12][7] ,
    \ix_double_ns[12][6] ,
    \ix_double_ns[12][5] ,
    \ix_double_ns[12][4] ,
    \ix_double_ns[12][3] ,
    \ix_double_ns[12][2] ,
    \ix_double_ns[12][1] ,
    \ix_double_ns[12][0] }),
    .north_single({\ix_single_ns[12][3] ,
    \ix_single_ns[12][2] ,
    \ix_single_ns[12][1] ,
    \ix_single_ns[12][0] }),
    .south_double({\ix_double_ns[5][7] ,
    \ix_double_ns[5][6] ,
    \ix_double_ns[5][5] ,
    \ix_double_ns[5][4] ,
    \ix_double_ns[5][3] ,
    \ix_double_ns[5][2] ,
    \ix_double_ns[5][1] ,
    \ix_double_ns[5][0] }),
    .south_single({\ix_single_ns[5][3] ,
    \ix_single_ns[5][2] ,
    \ix_single_ns[5][1] ,
    gpio_south[5]}),
    .west_double({\ix_double_ew[5][7] ,
    \ix_double_ew[5][6] ,
    \ix_double_ew[5][5] ,
    \ix_double_ew[5][4] ,
    \ix_double_ew[5][3] ,
    \ix_double_ew[5][2] ,
    \ix_double_ew[5][1] ,
    \ix_double_ew[5][0] }),
    .west_single({\ix_single_ew[5][3] ,
    \ix_single_ew[5][2] ,
    \ix_single_ew[5][1] ,
    \ix_single_ew[5][0] }));
 clb_tile \X[5].Y[1].clb  (.carry_in(\carry[1][5] ),
    .carry_out(\carry[2][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][5] ),
    .set_out_hard(\col_set[2][5] ),
    .shift_in_hard(\col_shift[1][5] ),
    .shift_out_hard(\col_shift[2][5] ),
    .cb_east_in({\dc_ew[14][4] ,
    \dc_ew[14][3] ,
    \dc_ew[14][2] ,
    \dc_ew[14][1] ,
    \dc_ew[14][0] }),
    .cb_east_out({\dc_we[14][9] ,
    \dc_we[14][8] ,
    \dc_we[14][7] ,
    \dc_we[14][6] ,
    \dc_we[14][5] ,
    \dc_we[14][4] ,
    \dc_we[14][3] ,
    \dc_we[14][2] ,
    \dc_we[14][1] ,
    \dc_we[14][0] }),
    .cb_north_in({\dc_ns[19][4] ,
    \dc_ns[19][3] ,
    \dc_ns[19][2] ,
    \dc_ns[19][1] ,
    \dc_ns[19][0] }),
    .cb_north_out({\dc_sn[19][9] ,
    \dc_sn[19][8] ,
    \dc_sn[19][7] ,
    \dc_sn[19][6] ,
    \dc_sn[19][5] ,
    \dc_sn[19][4] ,
    \dc_sn[19][3] ,
    \dc_sn[19][2] ,
    \dc_sn[19][1] ,
    \dc_sn[19][0] }),
    .clb_south_in({\dc_sn[12][9] ,
    \dc_sn[12][8] ,
    \dc_sn[12][7] ,
    \dc_sn[12][6] ,
    \dc_sn[12][5] ,
    \dc_sn[12][4] ,
    \dc_sn[12][3] ,
    \dc_sn[12][2] ,
    \dc_sn[12][1] ,
    \dc_sn[12][0] }),
    .clb_south_out({\dc_ns[12][4] ,
    \dc_ns[12][3] ,
    \dc_ns[12][2] ,
    \dc_ns[12][1] ,
    \dc_ns[12][0] }),
    .clb_west_in({\dc_we[13][9] ,
    \dc_we[13][8] ,
    \dc_we[13][7] ,
    \dc_we[13][6] ,
    \dc_we[13][5] ,
    \dc_we[13][4] ,
    \dc_we[13][3] ,
    \dc_we[13][2] ,
    \dc_we[13][1] ,
    \dc_we[13][0] }),
    .clb_west_out({\dc_ew[13][4] ,
    \dc_ew[13][3] ,
    \dc_ew[13][2] ,
    \dc_ew[13][1] ,
    \dc_ew[13][0] }),
    .east_double({\ix_double_ew[14][7] ,
    \ix_double_ew[14][6] ,
    \ix_double_ew[14][5] ,
    \ix_double_ew[14][4] ,
    \ix_double_ew[14][3] ,
    \ix_double_ew[14][2] ,
    \ix_double_ew[14][1] ,
    \ix_double_ew[14][0] }),
    .east_single({\ix_single_ew[14][3] ,
    \ix_single_ew[14][2] ,
    \ix_single_ew[14][1] ,
    \ix_single_ew[14][0] }),
    .north_double({\ix_double_ns[19][7] ,
    \ix_double_ns[19][6] ,
    \ix_double_ns[19][5] ,
    \ix_double_ns[19][4] ,
    \ix_double_ns[19][3] ,
    \ix_double_ns[19][2] ,
    \ix_double_ns[19][1] ,
    \ix_double_ns[19][0] }),
    .north_single({\ix_single_ns[19][3] ,
    \ix_single_ns[19][2] ,
    \ix_single_ns[19][1] ,
    \ix_single_ns[19][0] }),
    .south_double({\ix_double_ns[12][7] ,
    \ix_double_ns[12][6] ,
    \ix_double_ns[12][5] ,
    \ix_double_ns[12][4] ,
    \ix_double_ns[12][3] ,
    \ix_double_ns[12][2] ,
    \ix_double_ns[12][1] ,
    \ix_double_ns[12][0] }),
    .south_single({\ix_single_ns[12][3] ,
    \ix_single_ns[12][2] ,
    \ix_single_ns[12][1] ,
    \ix_single_ns[12][0] }),
    .west_double({\ix_double_ew[13][7] ,
    \ix_double_ew[13][6] ,
    \ix_double_ew[13][5] ,
    \ix_double_ew[13][4] ,
    \ix_double_ew[13][3] ,
    \ix_double_ew[13][2] ,
    \ix_double_ew[13][1] ,
    \ix_double_ew[13][0] }),
    .west_single({\ix_single_ew[13][3] ,
    \ix_single_ew[13][2] ,
    \ix_single_ew[13][1] ,
    \ix_single_ew[13][0] }));
 clb_tile \X[5].Y[2].clb  (.carry_in(\carry[2][5] ),
    .carry_out(\carry[3][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][5] ),
    .set_out_hard(\col_set[3][5] ),
    .shift_in_hard(\col_shift[2][5] ),
    .shift_out_hard(\col_shift[3][5] ),
    .cb_east_in({\dc_ew[22][4] ,
    \dc_ew[22][3] ,
    \dc_ew[22][2] ,
    \dc_ew[22][1] ,
    \dc_ew[22][0] }),
    .cb_east_out({\dc_we[22][9] ,
    \dc_we[22][8] ,
    \dc_we[22][7] ,
    \dc_we[22][6] ,
    \dc_we[22][5] ,
    \dc_we[22][4] ,
    \dc_we[22][3] ,
    \dc_we[22][2] ,
    \dc_we[22][1] ,
    \dc_we[22][0] }),
    .cb_north_in({\dc_ns[26][4] ,
    \dc_ns[26][3] ,
    \dc_ns[26][2] ,
    \dc_ns[26][1] ,
    \dc_ns[26][0] }),
    .cb_north_out({\dc_sn[26][9] ,
    \dc_sn[26][8] ,
    \dc_sn[26][7] ,
    \dc_sn[26][6] ,
    \dc_sn[26][5] ,
    \dc_sn[26][4] ,
    \dc_sn[26][3] ,
    \dc_sn[26][2] ,
    \dc_sn[26][1] ,
    \dc_sn[26][0] }),
    .clb_south_in({\dc_sn[19][9] ,
    \dc_sn[19][8] ,
    \dc_sn[19][7] ,
    \dc_sn[19][6] ,
    \dc_sn[19][5] ,
    \dc_sn[19][4] ,
    \dc_sn[19][3] ,
    \dc_sn[19][2] ,
    \dc_sn[19][1] ,
    \dc_sn[19][0] }),
    .clb_south_out({\dc_ns[19][4] ,
    \dc_ns[19][3] ,
    \dc_ns[19][2] ,
    \dc_ns[19][1] ,
    \dc_ns[19][0] }),
    .clb_west_in({\dc_we[21][9] ,
    \dc_we[21][8] ,
    \dc_we[21][7] ,
    \dc_we[21][6] ,
    \dc_we[21][5] ,
    \dc_we[21][4] ,
    \dc_we[21][3] ,
    \dc_we[21][2] ,
    \dc_we[21][1] ,
    \dc_we[21][0] }),
    .clb_west_out({\dc_ew[21][4] ,
    \dc_ew[21][3] ,
    \dc_ew[21][2] ,
    \dc_ew[21][1] ,
    \dc_ew[21][0] }),
    .east_double({\ix_double_ew[22][7] ,
    \ix_double_ew[22][6] ,
    \ix_double_ew[22][5] ,
    \ix_double_ew[22][4] ,
    \ix_double_ew[22][3] ,
    \ix_double_ew[22][2] ,
    \ix_double_ew[22][1] ,
    \ix_double_ew[22][0] }),
    .east_single({\ix_single_ew[22][3] ,
    \ix_single_ew[22][2] ,
    \ix_single_ew[22][1] ,
    \ix_single_ew[22][0] }),
    .north_double({\ix_double_ns[26][7] ,
    \ix_double_ns[26][6] ,
    \ix_double_ns[26][5] ,
    \ix_double_ns[26][4] ,
    \ix_double_ns[26][3] ,
    \ix_double_ns[26][2] ,
    \ix_double_ns[26][1] ,
    \ix_double_ns[26][0] }),
    .north_single({\ix_single_ns[26][3] ,
    \ix_single_ns[26][2] ,
    \ix_single_ns[26][1] ,
    \ix_single_ns[26][0] }),
    .south_double({\ix_double_ns[19][7] ,
    \ix_double_ns[19][6] ,
    \ix_double_ns[19][5] ,
    \ix_double_ns[19][4] ,
    \ix_double_ns[19][3] ,
    \ix_double_ns[19][2] ,
    \ix_double_ns[19][1] ,
    \ix_double_ns[19][0] }),
    .south_single({\ix_single_ns[19][3] ,
    \ix_single_ns[19][2] ,
    \ix_single_ns[19][1] ,
    \ix_single_ns[19][0] }),
    .west_double({\ix_double_ew[21][7] ,
    \ix_double_ew[21][6] ,
    \ix_double_ew[21][5] ,
    \ix_double_ew[21][4] ,
    \ix_double_ew[21][3] ,
    \ix_double_ew[21][2] ,
    \ix_double_ew[21][1] ,
    \ix_double_ew[21][0] }),
    .west_single({\ix_single_ew[21][3] ,
    \ix_single_ew[21][2] ,
    \ix_single_ew[21][1] ,
    \ix_single_ew[21][0] }));
 clb_tile \X[5].Y[3].clb  (.carry_in(\carry[3][5] ),
    .carry_out(\carry[4][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][5] ),
    .set_out_hard(\col_set[4][5] ),
    .shift_in_hard(\col_shift[3][5] ),
    .shift_out_hard(\col_shift[4][5] ),
    .cb_east_in({\dc_ew[30][4] ,
    \dc_ew[30][3] ,
    \dc_ew[30][2] ,
    \dc_ew[30][1] ,
    \dc_ew[30][0] }),
    .cb_east_out({\dc_we[30][9] ,
    \dc_we[30][8] ,
    \dc_we[30][7] ,
    \dc_we[30][6] ,
    \dc_we[30][5] ,
    \dc_we[30][4] ,
    \dc_we[30][3] ,
    \dc_we[30][2] ,
    \dc_we[30][1] ,
    \dc_we[30][0] }),
    .cb_north_in({\dc_ns[33][4] ,
    \dc_ns[33][3] ,
    \dc_ns[33][2] ,
    \dc_ns[33][1] ,
    \dc_ns[33][0] }),
    .cb_north_out({\dc_sn[33][9] ,
    \dc_sn[33][8] ,
    \dc_sn[33][7] ,
    \dc_sn[33][6] ,
    \dc_sn[33][5] ,
    \dc_sn[33][4] ,
    \dc_sn[33][3] ,
    \dc_sn[33][2] ,
    \dc_sn[33][1] ,
    \dc_sn[33][0] }),
    .clb_south_in({\dc_sn[26][9] ,
    \dc_sn[26][8] ,
    \dc_sn[26][7] ,
    \dc_sn[26][6] ,
    \dc_sn[26][5] ,
    \dc_sn[26][4] ,
    \dc_sn[26][3] ,
    \dc_sn[26][2] ,
    \dc_sn[26][1] ,
    \dc_sn[26][0] }),
    .clb_south_out({\dc_ns[26][4] ,
    \dc_ns[26][3] ,
    \dc_ns[26][2] ,
    \dc_ns[26][1] ,
    \dc_ns[26][0] }),
    .clb_west_in({\dc_we[29][9] ,
    \dc_we[29][8] ,
    \dc_we[29][7] ,
    \dc_we[29][6] ,
    \dc_we[29][5] ,
    \dc_we[29][4] ,
    \dc_we[29][3] ,
    \dc_we[29][2] ,
    \dc_we[29][1] ,
    \dc_we[29][0] }),
    .clb_west_out({\dc_ew[29][4] ,
    \dc_ew[29][3] ,
    \dc_ew[29][2] ,
    \dc_ew[29][1] ,
    \dc_ew[29][0] }),
    .east_double({\ix_double_ew[30][7] ,
    \ix_double_ew[30][6] ,
    \ix_double_ew[30][5] ,
    \ix_double_ew[30][4] ,
    \ix_double_ew[30][3] ,
    \ix_double_ew[30][2] ,
    \ix_double_ew[30][1] ,
    \ix_double_ew[30][0] }),
    .east_single({\ix_single_ew[30][3] ,
    \ix_single_ew[30][2] ,
    \ix_single_ew[30][1] ,
    \ix_single_ew[30][0] }),
    .north_double({\ix_double_ns[33][7] ,
    \ix_double_ns[33][6] ,
    \ix_double_ns[33][5] ,
    \ix_double_ns[33][4] ,
    \ix_double_ns[33][3] ,
    \ix_double_ns[33][2] ,
    \ix_double_ns[33][1] ,
    \ix_double_ns[33][0] }),
    .north_single({\ix_single_ns[33][3] ,
    \ix_single_ns[33][2] ,
    \ix_single_ns[33][1] ,
    \ix_single_ns[33][0] }),
    .south_double({\ix_double_ns[26][7] ,
    \ix_double_ns[26][6] ,
    \ix_double_ns[26][5] ,
    \ix_double_ns[26][4] ,
    \ix_double_ns[26][3] ,
    \ix_double_ns[26][2] ,
    \ix_double_ns[26][1] ,
    \ix_double_ns[26][0] }),
    .south_single({\ix_single_ns[26][3] ,
    \ix_single_ns[26][2] ,
    \ix_single_ns[26][1] ,
    \ix_single_ns[26][0] }),
    .west_double({\ix_double_ew[29][7] ,
    \ix_double_ew[29][6] ,
    \ix_double_ew[29][5] ,
    \ix_double_ew[29][4] ,
    \ix_double_ew[29][3] ,
    \ix_double_ew[29][2] ,
    \ix_double_ew[29][1] ,
    \ix_double_ew[29][0] }),
    .west_single({\ix_single_ew[29][3] ,
    \ix_single_ew[29][2] ,
    \ix_single_ew[29][1] ,
    \ix_single_ew[29][0] }));
 clb_tile \X[5].Y[4].clb  (.carry_in(\carry[4][5] ),
    .carry_out(\carry[5][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][5] ),
    .set_out_hard(\col_set[5][5] ),
    .shift_in_hard(\col_shift[4][5] ),
    .shift_out_hard(\col_shift[5][5] ),
    .cb_east_in({\dc_ew[38][4] ,
    \dc_ew[38][3] ,
    \dc_ew[38][2] ,
    \dc_ew[38][1] ,
    \dc_ew[38][0] }),
    .cb_east_out({\dc_we[38][9] ,
    \dc_we[38][8] ,
    \dc_we[38][7] ,
    \dc_we[38][6] ,
    \dc_we[38][5] ,
    \dc_we[38][4] ,
    \dc_we[38][3] ,
    \dc_we[38][2] ,
    \dc_we[38][1] ,
    \dc_we[38][0] }),
    .cb_north_in({\dc_ns[40][4] ,
    \dc_ns[40][3] ,
    \dc_ns[40][2] ,
    \dc_ns[40][1] ,
    \dc_ns[40][0] }),
    .cb_north_out({\dc_sn[40][9] ,
    \dc_sn[40][8] ,
    \dc_sn[40][7] ,
    \dc_sn[40][6] ,
    \dc_sn[40][5] ,
    \dc_sn[40][4] ,
    \dc_sn[40][3] ,
    \dc_sn[40][2] ,
    \dc_sn[40][1] ,
    \dc_sn[40][0] }),
    .clb_south_in({\dc_sn[33][9] ,
    \dc_sn[33][8] ,
    \dc_sn[33][7] ,
    \dc_sn[33][6] ,
    \dc_sn[33][5] ,
    \dc_sn[33][4] ,
    \dc_sn[33][3] ,
    \dc_sn[33][2] ,
    \dc_sn[33][1] ,
    \dc_sn[33][0] }),
    .clb_south_out({\dc_ns[33][4] ,
    \dc_ns[33][3] ,
    \dc_ns[33][2] ,
    \dc_ns[33][1] ,
    \dc_ns[33][0] }),
    .clb_west_in({\dc_we[37][9] ,
    \dc_we[37][8] ,
    \dc_we[37][7] ,
    \dc_we[37][6] ,
    \dc_we[37][5] ,
    \dc_we[37][4] ,
    \dc_we[37][3] ,
    \dc_we[37][2] ,
    \dc_we[37][1] ,
    \dc_we[37][0] }),
    .clb_west_out({\dc_ew[37][4] ,
    \dc_ew[37][3] ,
    \dc_ew[37][2] ,
    \dc_ew[37][1] ,
    \dc_ew[37][0] }),
    .east_double({\ix_double_ew[38][7] ,
    \ix_double_ew[38][6] ,
    \ix_double_ew[38][5] ,
    \ix_double_ew[38][4] ,
    \ix_double_ew[38][3] ,
    \ix_double_ew[38][2] ,
    \ix_double_ew[38][1] ,
    \ix_double_ew[38][0] }),
    .east_single({\ix_single_ew[38][3] ,
    \ix_single_ew[38][2] ,
    \ix_single_ew[38][1] ,
    \ix_single_ew[38][0] }),
    .north_double({\ix_double_ns[40][7] ,
    \ix_double_ns[40][6] ,
    \ix_double_ns[40][5] ,
    \ix_double_ns[40][4] ,
    \ix_double_ns[40][3] ,
    \ix_double_ns[40][2] ,
    \ix_double_ns[40][1] ,
    \ix_double_ns[40][0] }),
    .north_single({\ix_single_ns[40][3] ,
    \ix_single_ns[40][2] ,
    \ix_single_ns[40][1] ,
    \ix_single_ns[40][0] }),
    .south_double({\ix_double_ns[33][7] ,
    \ix_double_ns[33][6] ,
    \ix_double_ns[33][5] ,
    \ix_double_ns[33][4] ,
    \ix_double_ns[33][3] ,
    \ix_double_ns[33][2] ,
    \ix_double_ns[33][1] ,
    \ix_double_ns[33][0] }),
    .south_single({\ix_single_ns[33][3] ,
    \ix_single_ns[33][2] ,
    \ix_single_ns[33][1] ,
    \ix_single_ns[33][0] }),
    .west_double({\ix_double_ew[37][7] ,
    \ix_double_ew[37][6] ,
    \ix_double_ew[37][5] ,
    \ix_double_ew[37][4] ,
    \ix_double_ew[37][3] ,
    \ix_double_ew[37][2] ,
    \ix_double_ew[37][1] ,
    \ix_double_ew[37][0] }),
    .west_single({\ix_single_ew[37][3] ,
    \ix_single_ew[37][2] ,
    \ix_single_ew[37][1] ,
    \ix_single_ew[37][0] }));
 clb_tile \X[5].Y[5].clb  (.carry_in(\carry[5][5] ),
    .carry_out(\carry[6][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][5] ),
    .set_out_hard(\col_set[6][5] ),
    .shift_in_hard(\col_shift[5][5] ),
    .shift_out_hard(\col_shift[6][5] ),
    .cb_east_in({\dc_ew[46][4] ,
    \dc_ew[46][3] ,
    \dc_ew[46][2] ,
    \dc_ew[46][1] ,
    \dc_ew[46][0] }),
    .cb_east_out({\dc_we[46][9] ,
    \dc_we[46][8] ,
    \dc_we[46][7] ,
    \dc_we[46][6] ,
    \dc_we[46][5] ,
    \dc_we[46][4] ,
    \dc_we[46][3] ,
    \dc_we[46][2] ,
    \dc_we[46][1] ,
    \dc_we[46][0] }),
    .cb_north_in({\dc_ns[47][4] ,
    \dc_ns[47][3] ,
    \dc_ns[47][2] ,
    \dc_ns[47][1] ,
    \dc_ns[47][0] }),
    .cb_north_out({\dc_sn[47][9] ,
    \dc_sn[47][8] ,
    \dc_sn[47][7] ,
    \dc_sn[47][6] ,
    \dc_sn[47][5] ,
    \dc_sn[47][4] ,
    \dc_sn[47][3] ,
    \dc_sn[47][2] ,
    \dc_sn[47][1] ,
    \dc_sn[47][0] }),
    .clb_south_in({\dc_sn[40][9] ,
    \dc_sn[40][8] ,
    \dc_sn[40][7] ,
    \dc_sn[40][6] ,
    \dc_sn[40][5] ,
    \dc_sn[40][4] ,
    \dc_sn[40][3] ,
    \dc_sn[40][2] ,
    \dc_sn[40][1] ,
    \dc_sn[40][0] }),
    .clb_south_out({\dc_ns[40][4] ,
    \dc_ns[40][3] ,
    \dc_ns[40][2] ,
    \dc_ns[40][1] ,
    \dc_ns[40][0] }),
    .clb_west_in({\dc_we[45][9] ,
    \dc_we[45][8] ,
    \dc_we[45][7] ,
    \dc_we[45][6] ,
    \dc_we[45][5] ,
    \dc_we[45][4] ,
    \dc_we[45][3] ,
    \dc_we[45][2] ,
    \dc_we[45][1] ,
    \dc_we[45][0] }),
    .clb_west_out({\dc_ew[45][4] ,
    \dc_ew[45][3] ,
    \dc_ew[45][2] ,
    \dc_ew[45][1] ,
    \dc_ew[45][0] }),
    .east_double({\ix_double_ew[46][7] ,
    \ix_double_ew[46][6] ,
    \ix_double_ew[46][5] ,
    \ix_double_ew[46][4] ,
    \ix_double_ew[46][3] ,
    \ix_double_ew[46][2] ,
    \ix_double_ew[46][1] ,
    \ix_double_ew[46][0] }),
    .east_single({\ix_single_ew[46][3] ,
    \ix_single_ew[46][2] ,
    \ix_single_ew[46][1] ,
    \ix_single_ew[46][0] }),
    .north_double({\ix_double_ns[47][7] ,
    \ix_double_ns[47][6] ,
    \ix_double_ns[47][5] ,
    \ix_double_ns[47][4] ,
    \ix_double_ns[47][3] ,
    \ix_double_ns[47][2] ,
    \ix_double_ns[47][1] ,
    \ix_double_ns[47][0] }),
    .north_single({\ix_single_ns[47][3] ,
    \ix_single_ns[47][2] ,
    \ix_single_ns[47][1] ,
    \ix_single_ns[47][0] }),
    .south_double({\ix_double_ns[40][7] ,
    \ix_double_ns[40][6] ,
    \ix_double_ns[40][5] ,
    \ix_double_ns[40][4] ,
    \ix_double_ns[40][3] ,
    \ix_double_ns[40][2] ,
    \ix_double_ns[40][1] ,
    \ix_double_ns[40][0] }),
    .south_single({\ix_single_ns[40][3] ,
    \ix_single_ns[40][2] ,
    \ix_single_ns[40][1] ,
    \ix_single_ns[40][0] }),
    .west_double({\ix_double_ew[45][7] ,
    \ix_double_ew[45][6] ,
    \ix_double_ew[45][5] ,
    \ix_double_ew[45][4] ,
    \ix_double_ew[45][3] ,
    \ix_double_ew[45][2] ,
    \ix_double_ew[45][1] ,
    \ix_double_ew[45][0] }),
    .west_single({\ix_single_ew[45][3] ,
    \ix_single_ew[45][2] ,
    \ix_single_ew[45][1] ,
    \ix_single_ew[45][0] }));
 clb_tile \X[5].Y[6].clb  (.carry_in(\carry[6][5] ),
    .carry_out(\carry[7][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][5] ),
    .set_out_hard(\col_set[7][5] ),
    .shift_in_hard(\col_shift[6][5] ),
    .shift_out_hard(\col_shift[7][5] ),
    .cb_east_in({\dc_ew[54][4] ,
    \dc_ew[54][3] ,
    \dc_ew[54][2] ,
    \dc_ew[54][1] ,
    \dc_ew[54][0] }),
    .cb_east_out({\dc_we[54][9] ,
    \dc_we[54][8] ,
    \dc_we[54][7] ,
    \dc_we[54][6] ,
    \dc_we[54][5] ,
    \dc_we[54][4] ,
    \dc_we[54][3] ,
    \dc_we[54][2] ,
    \dc_we[54][1] ,
    \dc_we[54][0] }),
    .cb_north_in({\dc_ns[54][4] ,
    \dc_ns[54][3] ,
    \dc_ns[54][2] ,
    \dc_ns[54][1] ,
    \dc_ns[54][0] }),
    .cb_north_out({\dc_sn[54][9] ,
    \dc_sn[54][8] ,
    \dc_sn[54][7] ,
    \dc_sn[54][6] ,
    \dc_sn[54][5] ,
    \dc_sn[54][4] ,
    \dc_sn[54][3] ,
    \dc_sn[54][2] ,
    \dc_sn[54][1] ,
    \dc_sn[54][0] }),
    .clb_south_in({\dc_sn[47][9] ,
    \dc_sn[47][8] ,
    \dc_sn[47][7] ,
    \dc_sn[47][6] ,
    \dc_sn[47][5] ,
    \dc_sn[47][4] ,
    \dc_sn[47][3] ,
    \dc_sn[47][2] ,
    \dc_sn[47][1] ,
    \dc_sn[47][0] }),
    .clb_south_out({\dc_ns[47][4] ,
    \dc_ns[47][3] ,
    \dc_ns[47][2] ,
    \dc_ns[47][1] ,
    \dc_ns[47][0] }),
    .clb_west_in({\dc_we[53][9] ,
    \dc_we[53][8] ,
    \dc_we[53][7] ,
    \dc_we[53][6] ,
    \dc_we[53][5] ,
    \dc_we[53][4] ,
    \dc_we[53][3] ,
    \dc_we[53][2] ,
    \dc_we[53][1] ,
    \dc_we[53][0] }),
    .clb_west_out({\dc_ew[53][4] ,
    \dc_ew[53][3] ,
    \dc_ew[53][2] ,
    \dc_ew[53][1] ,
    \dc_ew[53][0] }),
    .east_double({\ix_double_ew[54][7] ,
    \ix_double_ew[54][6] ,
    \ix_double_ew[54][5] ,
    \ix_double_ew[54][4] ,
    \ix_double_ew[54][3] ,
    \ix_double_ew[54][2] ,
    \ix_double_ew[54][1] ,
    \ix_double_ew[54][0] }),
    .east_single({\ix_single_ew[54][3] ,
    \ix_single_ew[54][2] ,
    \ix_single_ew[54][1] ,
    \ix_single_ew[54][0] }),
    .north_double({\ix_double_ns[54][7] ,
    \ix_double_ns[54][6] ,
    \ix_double_ns[54][5] ,
    \ix_double_ns[54][4] ,
    \ix_double_ns[54][3] ,
    \ix_double_ns[54][2] ,
    \ix_double_ns[54][1] ,
    \ix_double_ns[54][0] }),
    .north_single({\ix_single_ns[54][3] ,
    \ix_single_ns[54][2] ,
    \ix_single_ns[54][1] ,
    \ix_single_ns[54][0] }),
    .south_double({\ix_double_ns[47][7] ,
    \ix_double_ns[47][6] ,
    \ix_double_ns[47][5] ,
    \ix_double_ns[47][4] ,
    \ix_double_ns[47][3] ,
    \ix_double_ns[47][2] ,
    \ix_double_ns[47][1] ,
    \ix_double_ns[47][0] }),
    .south_single({\ix_single_ns[47][3] ,
    \ix_single_ns[47][2] ,
    \ix_single_ns[47][1] ,
    \ix_single_ns[47][0] }),
    .west_double({\ix_double_ew[53][7] ,
    \ix_double_ew[53][6] ,
    \ix_double_ew[53][5] ,
    \ix_double_ew[53][4] ,
    \ix_double_ew[53][3] ,
    \ix_double_ew[53][2] ,
    \ix_double_ew[53][1] ,
    \ix_double_ew[53][0] }),
    .west_single({\ix_single_ew[53][3] ,
    \ix_single_ew[53][2] ,
    \ix_single_ew[53][1] ,
    \ix_single_ew[53][0] }));
 clb_tile \X[5].Y[7].clb  (.carry_in(\carry[7][5] ),
    .carry_out(\carry[8][5] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][5] ),
    .set_out_hard(\col_set[8][5] ),
    .shift_in_hard(\col_shift[7][5] ),
    .shift_out_hard(\col_shift[8][5] ),
    .cb_east_in({\dc_ew[62][4] ,
    \dc_ew[62][3] ,
    \dc_ew[62][2] ,
    \dc_ew[62][1] ,
    \dc_ew[62][0] }),
    .cb_east_out({\dc_we[62][9] ,
    \dc_we[62][8] ,
    \dc_we[62][7] ,
    \dc_we[62][6] ,
    \dc_we[62][5] ,
    \dc_we[62][4] ,
    \dc_we[62][3] ,
    \dc_we[62][2] ,
    \dc_we[62][1] ,
    \dc_we[62][0] }),
    .cb_north_in({_175_,
    _174_,
    _173_,
    _172_,
    _171_}),
    .cb_north_out({\dc_sn[61][9] ,
    \dc_sn[61][8] ,
    \dc_sn[61][7] ,
    \dc_sn[61][6] ,
    \dc_sn[61][5] ,
    \dc_sn[61][4] ,
    \dc_sn[61][3] ,
    \dc_sn[61][2] ,
    \dc_sn[61][1] ,
    \dc_sn[61][0] }),
    .clb_south_in({\dc_sn[54][9] ,
    \dc_sn[54][8] ,
    \dc_sn[54][7] ,
    \dc_sn[54][6] ,
    \dc_sn[54][5] ,
    \dc_sn[54][4] ,
    \dc_sn[54][3] ,
    \dc_sn[54][2] ,
    \dc_sn[54][1] ,
    \dc_sn[54][0] }),
    .clb_south_out({\dc_ns[54][4] ,
    \dc_ns[54][3] ,
    \dc_ns[54][2] ,
    \dc_ns[54][1] ,
    \dc_ns[54][0] }),
    .clb_west_in({\dc_we[61][9] ,
    \dc_we[61][8] ,
    \dc_we[61][7] ,
    \dc_we[61][6] ,
    \dc_we[61][5] ,
    \dc_we[61][4] ,
    \dc_we[61][3] ,
    \dc_we[61][2] ,
    \dc_we[61][1] ,
    \dc_we[61][0] }),
    .clb_west_out({\dc_ew[61][4] ,
    \dc_ew[61][3] ,
    \dc_ew[61][2] ,
    \dc_ew[61][1] ,
    \dc_ew[61][0] }),
    .east_double({\ix_double_ew[62][7] ,
    \ix_double_ew[62][6] ,
    \ix_double_ew[62][5] ,
    \ix_double_ew[62][4] ,
    \ix_double_ew[62][3] ,
    \ix_double_ew[62][2] ,
    \ix_double_ew[62][1] ,
    \ix_double_ew[62][0] }),
    .east_single({\ix_single_ew[62][3] ,
    \ix_single_ew[62][2] ,
    \ix_single_ew[62][1] ,
    \ix_single_ew[62][0] }),
    .north_double({\ix_double_ns[61][7] ,
    \ix_double_ns[61][6] ,
    \ix_double_ns[61][5] ,
    \ix_double_ns[61][4] ,
    \ix_double_ns[61][3] ,
    \ix_double_ns[61][2] ,
    \ix_double_ns[61][1] ,
    \ix_double_ns[61][0] }),
    .north_single({\ix_single_ns[61][3] ,
    \ix_single_ns[61][2] ,
    \ix_single_ns[61][1] ,
    gpio_north[5]}),
    .south_double({\ix_double_ns[54][7] ,
    \ix_double_ns[54][6] ,
    \ix_double_ns[54][5] ,
    \ix_double_ns[54][4] ,
    \ix_double_ns[54][3] ,
    \ix_double_ns[54][2] ,
    \ix_double_ns[54][1] ,
    \ix_double_ns[54][0] }),
    .south_single({\ix_single_ns[54][3] ,
    \ix_single_ns[54][2] ,
    \ix_single_ns[54][1] ,
    \ix_single_ns[54][0] }),
    .west_double({\ix_double_ew[61][7] ,
    \ix_double_ew[61][6] ,
    \ix_double_ew[61][5] ,
    \ix_double_ew[61][4] ,
    \ix_double_ew[61][3] ,
    \ix_double_ew[61][2] ,
    \ix_double_ew[61][1] ,
    \ix_double_ew[61][0] }),
    .west_single({\ix_single_ew[61][3] ,
    \ix_single_ew[61][2] ,
    \ix_single_ew[61][1] ,
    \ix_single_ew[61][0] }));
 clb_tile \X[6].Y[0].clb  (.carry_in(_176_),
    .carry_out(\carry[1][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\wb_set_out[1][2] ),
    .set_out_hard(\col_set[1][6] ),
    .shift_in_hard(\wb_shift_out[1][2] ),
    .shift_out_hard(\col_shift[1][6] ),
    .cb_east_in({_181_,
    _180_,
    _179_,
    _178_,
    _177_}),
    .cb_east_out({\dc_we[7][9] ,
    \dc_we[7][8] ,
    \dc_we[7][7] ,
    \dc_we[7][6] ,
    \dc_we[7][5] ,
    \dc_we[7][4] ,
    \dc_we[7][3] ,
    \dc_we[7][2] ,
    \dc_we[7][1] ,
    \dc_we[7][0] }),
    .cb_north_in({\dc_ns[13][4] ,
    \dc_ns[13][3] ,
    \dc_ns[13][2] ,
    \dc_ns[13][1] ,
    \dc_ns[13][0] }),
    .cb_north_out({\dc_sn[13][9] ,
    \dc_sn[13][8] ,
    \dc_sn[13][7] ,
    \dc_sn[13][6] ,
    \dc_sn[13][5] ,
    \dc_sn[13][4] ,
    \dc_sn[13][3] ,
    \dc_sn[13][2] ,
    \dc_sn[13][1] ,
    \dc_sn[13][0] }),
    .clb_south_in({_191_,
    _190_,
    _189_,
    _188_,
    _187_,
    _186_,
    _185_,
    _184_,
    _183_,
    _182_}),
    .clb_south_out({\dc_ns[6][4] ,
    \dc_ns[6][3] ,
    \dc_ns[6][2] ,
    \dc_ns[6][1] ,
    \dc_ns[6][0] }),
    .clb_west_in({\dc_we[6][9] ,
    \dc_we[6][8] ,
    \dc_we[6][7] ,
    \dc_we[6][6] ,
    \dc_we[6][5] ,
    \dc_we[6][4] ,
    \dc_we[6][3] ,
    \dc_we[6][2] ,
    \dc_we[6][1] ,
    \dc_we[6][0] }),
    .clb_west_out({\dc_ew[6][4] ,
    \dc_ew[6][3] ,
    \dc_ew[6][2] ,
    \dc_ew[6][1] ,
    \dc_ew[6][0] }),
    .east_double({\ix_double_ew[7][7] ,
    \ix_double_ew[7][6] ,
    \ix_double_ew[7][5] ,
    \ix_double_ew[7][4] ,
    \ix_double_ew[7][3] ,
    \ix_double_ew[7][2] ,
    \ix_double_ew[7][1] ,
    \ix_double_ew[7][0] }),
    .east_single({\ix_single_ew[7][3] ,
    \ix_single_ew[7][2] ,
    \ix_single_ew[7][1] ,
    gpio_east[0]}),
    .north_double({\ix_double_ns[13][7] ,
    \ix_double_ns[13][6] ,
    \ix_double_ns[13][5] ,
    \ix_double_ns[13][4] ,
    \ix_double_ns[13][3] ,
    \ix_double_ns[13][2] ,
    \ix_double_ns[13][1] ,
    \ix_double_ns[13][0] }),
    .north_single({\ix_single_ns[13][3] ,
    \ix_single_ns[13][2] ,
    \ix_single_ns[13][1] ,
    \ix_single_ns[13][0] }),
    .south_double({\ix_double_ns[6][7] ,
    \ix_double_ns[6][6] ,
    \ix_double_ns[6][5] ,
    \ix_double_ns[6][4] ,
    \ix_double_ns[6][3] ,
    \ix_double_ns[6][2] ,
    \ix_double_ns[6][1] ,
    \ix_double_ns[6][0] }),
    .south_single({\ix_single_ns[6][3] ,
    \ix_single_ns[6][2] ,
    \ix_single_ns[6][1] ,
    gpio_south[6]}),
    .west_double({\ix_double_ew[6][7] ,
    \ix_double_ew[6][6] ,
    \ix_double_ew[6][5] ,
    \ix_double_ew[6][4] ,
    \ix_double_ew[6][3] ,
    \ix_double_ew[6][2] ,
    \ix_double_ew[6][1] ,
    \ix_double_ew[6][0] }),
    .west_single({\ix_single_ew[6][3] ,
    \ix_single_ew[6][2] ,
    \ix_single_ew[6][1] ,
    \ix_single_ew[6][0] }));
 clb_tile \X[6].Y[1].clb  (.carry_in(\carry[1][6] ),
    .carry_out(\carry[2][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[1][6] ),
    .set_out_hard(\col_set[2][6] ),
    .shift_in_hard(\col_shift[1][6] ),
    .shift_out_hard(\col_shift[2][6] ),
    .cb_east_in({_196_,
    _195_,
    _194_,
    _193_,
    _192_}),
    .cb_east_out({\dc_we[15][9] ,
    \dc_we[15][8] ,
    \dc_we[15][7] ,
    \dc_we[15][6] ,
    \dc_we[15][5] ,
    \dc_we[15][4] ,
    \dc_we[15][3] ,
    \dc_we[15][2] ,
    \dc_we[15][1] ,
    \dc_we[15][0] }),
    .cb_north_in({\dc_ns[20][4] ,
    \dc_ns[20][3] ,
    \dc_ns[20][2] ,
    \dc_ns[20][1] ,
    \dc_ns[20][0] }),
    .cb_north_out({\dc_sn[20][9] ,
    \dc_sn[20][8] ,
    \dc_sn[20][7] ,
    \dc_sn[20][6] ,
    \dc_sn[20][5] ,
    \dc_sn[20][4] ,
    \dc_sn[20][3] ,
    \dc_sn[20][2] ,
    \dc_sn[20][1] ,
    \dc_sn[20][0] }),
    .clb_south_in({\dc_sn[13][9] ,
    \dc_sn[13][8] ,
    \dc_sn[13][7] ,
    \dc_sn[13][6] ,
    \dc_sn[13][5] ,
    \dc_sn[13][4] ,
    \dc_sn[13][3] ,
    \dc_sn[13][2] ,
    \dc_sn[13][1] ,
    \dc_sn[13][0] }),
    .clb_south_out({\dc_ns[13][4] ,
    \dc_ns[13][3] ,
    \dc_ns[13][2] ,
    \dc_ns[13][1] ,
    \dc_ns[13][0] }),
    .clb_west_in({\dc_we[14][9] ,
    \dc_we[14][8] ,
    \dc_we[14][7] ,
    \dc_we[14][6] ,
    \dc_we[14][5] ,
    \dc_we[14][4] ,
    \dc_we[14][3] ,
    \dc_we[14][2] ,
    \dc_we[14][1] ,
    \dc_we[14][0] }),
    .clb_west_out({\dc_ew[14][4] ,
    \dc_ew[14][3] ,
    \dc_ew[14][2] ,
    \dc_ew[14][1] ,
    \dc_ew[14][0] }),
    .east_double({\ix_double_ew[15][7] ,
    \ix_double_ew[15][6] ,
    \ix_double_ew[15][5] ,
    \ix_double_ew[15][4] ,
    \ix_double_ew[15][3] ,
    \ix_double_ew[15][2] ,
    \ix_double_ew[15][1] ,
    \ix_double_ew[15][0] }),
    .east_single({\ix_single_ew[15][3] ,
    \ix_single_ew[15][2] ,
    \ix_single_ew[15][1] ,
    gpio_east[1]}),
    .north_double({\ix_double_ns[20][7] ,
    \ix_double_ns[20][6] ,
    \ix_double_ns[20][5] ,
    \ix_double_ns[20][4] ,
    \ix_double_ns[20][3] ,
    \ix_double_ns[20][2] ,
    \ix_double_ns[20][1] ,
    \ix_double_ns[20][0] }),
    .north_single({\ix_single_ns[20][3] ,
    \ix_single_ns[20][2] ,
    \ix_single_ns[20][1] ,
    \ix_single_ns[20][0] }),
    .south_double({\ix_double_ns[13][7] ,
    \ix_double_ns[13][6] ,
    \ix_double_ns[13][5] ,
    \ix_double_ns[13][4] ,
    \ix_double_ns[13][3] ,
    \ix_double_ns[13][2] ,
    \ix_double_ns[13][1] ,
    \ix_double_ns[13][0] }),
    .south_single({\ix_single_ns[13][3] ,
    \ix_single_ns[13][2] ,
    \ix_single_ns[13][1] ,
    \ix_single_ns[13][0] }),
    .west_double({\ix_double_ew[14][7] ,
    \ix_double_ew[14][6] ,
    \ix_double_ew[14][5] ,
    \ix_double_ew[14][4] ,
    \ix_double_ew[14][3] ,
    \ix_double_ew[14][2] ,
    \ix_double_ew[14][1] ,
    \ix_double_ew[14][0] }),
    .west_single({\ix_single_ew[14][3] ,
    \ix_single_ew[14][2] ,
    \ix_single_ew[14][1] ,
    \ix_single_ew[14][0] }));
 clb_tile \X[6].Y[2].clb  (.carry_in(\carry[2][6] ),
    .carry_out(\carry[3][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[2][6] ),
    .set_out_hard(\col_set[3][6] ),
    .shift_in_hard(\col_shift[2][6] ),
    .shift_out_hard(\col_shift[3][6] ),
    .cb_east_in({_201_,
    _200_,
    _199_,
    _198_,
    _197_}),
    .cb_east_out({\dc_we[23][9] ,
    \dc_we[23][8] ,
    \dc_we[23][7] ,
    \dc_we[23][6] ,
    \dc_we[23][5] ,
    \dc_we[23][4] ,
    \dc_we[23][3] ,
    \dc_we[23][2] ,
    \dc_we[23][1] ,
    \dc_we[23][0] }),
    .cb_north_in({\dc_ns[27][4] ,
    \dc_ns[27][3] ,
    \dc_ns[27][2] ,
    \dc_ns[27][1] ,
    \dc_ns[27][0] }),
    .cb_north_out({\dc_sn[27][9] ,
    \dc_sn[27][8] ,
    \dc_sn[27][7] ,
    \dc_sn[27][6] ,
    \dc_sn[27][5] ,
    \dc_sn[27][4] ,
    \dc_sn[27][3] ,
    \dc_sn[27][2] ,
    \dc_sn[27][1] ,
    \dc_sn[27][0] }),
    .clb_south_in({\dc_sn[20][9] ,
    \dc_sn[20][8] ,
    \dc_sn[20][7] ,
    \dc_sn[20][6] ,
    \dc_sn[20][5] ,
    \dc_sn[20][4] ,
    \dc_sn[20][3] ,
    \dc_sn[20][2] ,
    \dc_sn[20][1] ,
    \dc_sn[20][0] }),
    .clb_south_out({\dc_ns[20][4] ,
    \dc_ns[20][3] ,
    \dc_ns[20][2] ,
    \dc_ns[20][1] ,
    \dc_ns[20][0] }),
    .clb_west_in({\dc_we[22][9] ,
    \dc_we[22][8] ,
    \dc_we[22][7] ,
    \dc_we[22][6] ,
    \dc_we[22][5] ,
    \dc_we[22][4] ,
    \dc_we[22][3] ,
    \dc_we[22][2] ,
    \dc_we[22][1] ,
    \dc_we[22][0] }),
    .clb_west_out({\dc_ew[22][4] ,
    \dc_ew[22][3] ,
    \dc_ew[22][2] ,
    \dc_ew[22][1] ,
    \dc_ew[22][0] }),
    .east_double({\ix_double_ew[23][7] ,
    \ix_double_ew[23][6] ,
    \ix_double_ew[23][5] ,
    \ix_double_ew[23][4] ,
    \ix_double_ew[23][3] ,
    \ix_double_ew[23][2] ,
    \ix_double_ew[23][1] ,
    \ix_double_ew[23][0] }),
    .east_single({\ix_single_ew[23][3] ,
    \ix_single_ew[23][2] ,
    \ix_single_ew[23][1] ,
    gpio_east[2]}),
    .north_double({\ix_double_ns[27][7] ,
    \ix_double_ns[27][6] ,
    \ix_double_ns[27][5] ,
    \ix_double_ns[27][4] ,
    \ix_double_ns[27][3] ,
    \ix_double_ns[27][2] ,
    \ix_double_ns[27][1] ,
    \ix_double_ns[27][0] }),
    .north_single({\ix_single_ns[27][3] ,
    \ix_single_ns[27][2] ,
    \ix_single_ns[27][1] ,
    \ix_single_ns[27][0] }),
    .south_double({\ix_double_ns[20][7] ,
    \ix_double_ns[20][6] ,
    \ix_double_ns[20][5] ,
    \ix_double_ns[20][4] ,
    \ix_double_ns[20][3] ,
    \ix_double_ns[20][2] ,
    \ix_double_ns[20][1] ,
    \ix_double_ns[20][0] }),
    .south_single({\ix_single_ns[20][3] ,
    \ix_single_ns[20][2] ,
    \ix_single_ns[20][1] ,
    \ix_single_ns[20][0] }),
    .west_double({\ix_double_ew[22][7] ,
    \ix_double_ew[22][6] ,
    \ix_double_ew[22][5] ,
    \ix_double_ew[22][4] ,
    \ix_double_ew[22][3] ,
    \ix_double_ew[22][2] ,
    \ix_double_ew[22][1] ,
    \ix_double_ew[22][0] }),
    .west_single({\ix_single_ew[22][3] ,
    \ix_single_ew[22][2] ,
    \ix_single_ew[22][1] ,
    \ix_single_ew[22][0] }));
 clb_tile \X[6].Y[3].clb  (.carry_in(\carry[3][6] ),
    .carry_out(\carry[4][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[3][6] ),
    .set_out_hard(\col_set[4][6] ),
    .shift_in_hard(\col_shift[3][6] ),
    .shift_out_hard(\col_shift[4][6] ),
    .cb_east_in({_206_,
    _205_,
    _204_,
    _203_,
    _202_}),
    .cb_east_out({\dc_we[31][9] ,
    \dc_we[31][8] ,
    \dc_we[31][7] ,
    \dc_we[31][6] ,
    \dc_we[31][5] ,
    \dc_we[31][4] ,
    \dc_we[31][3] ,
    \dc_we[31][2] ,
    \dc_we[31][1] ,
    \dc_we[31][0] }),
    .cb_north_in({\dc_ns[34][4] ,
    \dc_ns[34][3] ,
    \dc_ns[34][2] ,
    \dc_ns[34][1] ,
    \dc_ns[34][0] }),
    .cb_north_out({\dc_sn[34][9] ,
    \dc_sn[34][8] ,
    \dc_sn[34][7] ,
    \dc_sn[34][6] ,
    \dc_sn[34][5] ,
    \dc_sn[34][4] ,
    \dc_sn[34][3] ,
    \dc_sn[34][2] ,
    \dc_sn[34][1] ,
    \dc_sn[34][0] }),
    .clb_south_in({\dc_sn[27][9] ,
    \dc_sn[27][8] ,
    \dc_sn[27][7] ,
    \dc_sn[27][6] ,
    \dc_sn[27][5] ,
    \dc_sn[27][4] ,
    \dc_sn[27][3] ,
    \dc_sn[27][2] ,
    \dc_sn[27][1] ,
    \dc_sn[27][0] }),
    .clb_south_out({\dc_ns[27][4] ,
    \dc_ns[27][3] ,
    \dc_ns[27][2] ,
    \dc_ns[27][1] ,
    \dc_ns[27][0] }),
    .clb_west_in({\dc_we[30][9] ,
    \dc_we[30][8] ,
    \dc_we[30][7] ,
    \dc_we[30][6] ,
    \dc_we[30][5] ,
    \dc_we[30][4] ,
    \dc_we[30][3] ,
    \dc_we[30][2] ,
    \dc_we[30][1] ,
    \dc_we[30][0] }),
    .clb_west_out({\dc_ew[30][4] ,
    \dc_ew[30][3] ,
    \dc_ew[30][2] ,
    \dc_ew[30][1] ,
    \dc_ew[30][0] }),
    .east_double({\ix_double_ew[31][7] ,
    \ix_double_ew[31][6] ,
    \ix_double_ew[31][5] ,
    \ix_double_ew[31][4] ,
    \ix_double_ew[31][3] ,
    \ix_double_ew[31][2] ,
    \ix_double_ew[31][1] ,
    \ix_double_ew[31][0] }),
    .east_single({\ix_single_ew[31][3] ,
    \ix_single_ew[31][2] ,
    \ix_single_ew[31][1] ,
    gpio_east[3]}),
    .north_double({\ix_double_ns[34][7] ,
    \ix_double_ns[34][6] ,
    \ix_double_ns[34][5] ,
    \ix_double_ns[34][4] ,
    \ix_double_ns[34][3] ,
    \ix_double_ns[34][2] ,
    \ix_double_ns[34][1] ,
    \ix_double_ns[34][0] }),
    .north_single({\ix_single_ns[34][3] ,
    \ix_single_ns[34][2] ,
    \ix_single_ns[34][1] ,
    \ix_single_ns[34][0] }),
    .south_double({\ix_double_ns[27][7] ,
    \ix_double_ns[27][6] ,
    \ix_double_ns[27][5] ,
    \ix_double_ns[27][4] ,
    \ix_double_ns[27][3] ,
    \ix_double_ns[27][2] ,
    \ix_double_ns[27][1] ,
    \ix_double_ns[27][0] }),
    .south_single({\ix_single_ns[27][3] ,
    \ix_single_ns[27][2] ,
    \ix_single_ns[27][1] ,
    \ix_single_ns[27][0] }),
    .west_double({\ix_double_ew[30][7] ,
    \ix_double_ew[30][6] ,
    \ix_double_ew[30][5] ,
    \ix_double_ew[30][4] ,
    \ix_double_ew[30][3] ,
    \ix_double_ew[30][2] ,
    \ix_double_ew[30][1] ,
    \ix_double_ew[30][0] }),
    .west_single({\ix_single_ew[30][3] ,
    \ix_single_ew[30][2] ,
    \ix_single_ew[30][1] ,
    \ix_single_ew[30][0] }));
 clb_tile \X[6].Y[4].clb  (.carry_in(\carry[4][6] ),
    .carry_out(\carry[5][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[4][6] ),
    .set_out_hard(\col_set[5][6] ),
    .shift_in_hard(\col_shift[4][6] ),
    .shift_out_hard(\col_shift[5][6] ),
    .cb_east_in({_211_,
    _210_,
    _209_,
    _208_,
    _207_}),
    .cb_east_out({\dc_we[39][9] ,
    \dc_we[39][8] ,
    \dc_we[39][7] ,
    \dc_we[39][6] ,
    \dc_we[39][5] ,
    \dc_we[39][4] ,
    \dc_we[39][3] ,
    \dc_we[39][2] ,
    \dc_we[39][1] ,
    \dc_we[39][0] }),
    .cb_north_in({\dc_ns[41][4] ,
    \dc_ns[41][3] ,
    \dc_ns[41][2] ,
    \dc_ns[41][1] ,
    \dc_ns[41][0] }),
    .cb_north_out({\dc_sn[41][9] ,
    \dc_sn[41][8] ,
    \dc_sn[41][7] ,
    \dc_sn[41][6] ,
    \dc_sn[41][5] ,
    \dc_sn[41][4] ,
    \dc_sn[41][3] ,
    \dc_sn[41][2] ,
    \dc_sn[41][1] ,
    \dc_sn[41][0] }),
    .clb_south_in({\dc_sn[34][9] ,
    \dc_sn[34][8] ,
    \dc_sn[34][7] ,
    \dc_sn[34][6] ,
    \dc_sn[34][5] ,
    \dc_sn[34][4] ,
    \dc_sn[34][3] ,
    \dc_sn[34][2] ,
    \dc_sn[34][1] ,
    \dc_sn[34][0] }),
    .clb_south_out({\dc_ns[34][4] ,
    \dc_ns[34][3] ,
    \dc_ns[34][2] ,
    \dc_ns[34][1] ,
    \dc_ns[34][0] }),
    .clb_west_in({\dc_we[38][9] ,
    \dc_we[38][8] ,
    \dc_we[38][7] ,
    \dc_we[38][6] ,
    \dc_we[38][5] ,
    \dc_we[38][4] ,
    \dc_we[38][3] ,
    \dc_we[38][2] ,
    \dc_we[38][1] ,
    \dc_we[38][0] }),
    .clb_west_out({\dc_ew[38][4] ,
    \dc_ew[38][3] ,
    \dc_ew[38][2] ,
    \dc_ew[38][1] ,
    \dc_ew[38][0] }),
    .east_double({\ix_double_ew[39][7] ,
    \ix_double_ew[39][6] ,
    \ix_double_ew[39][5] ,
    \ix_double_ew[39][4] ,
    \ix_double_ew[39][3] ,
    \ix_double_ew[39][2] ,
    \ix_double_ew[39][1] ,
    \ix_double_ew[39][0] }),
    .east_single({\ix_single_ew[39][3] ,
    \ix_single_ew[39][2] ,
    \ix_single_ew[39][1] ,
    gpio_east[4]}),
    .north_double({\ix_double_ns[41][7] ,
    \ix_double_ns[41][6] ,
    \ix_double_ns[41][5] ,
    \ix_double_ns[41][4] ,
    \ix_double_ns[41][3] ,
    \ix_double_ns[41][2] ,
    \ix_double_ns[41][1] ,
    \ix_double_ns[41][0] }),
    .north_single({\ix_single_ns[41][3] ,
    \ix_single_ns[41][2] ,
    \ix_single_ns[41][1] ,
    \ix_single_ns[41][0] }),
    .south_double({\ix_double_ns[34][7] ,
    \ix_double_ns[34][6] ,
    \ix_double_ns[34][5] ,
    \ix_double_ns[34][4] ,
    \ix_double_ns[34][3] ,
    \ix_double_ns[34][2] ,
    \ix_double_ns[34][1] ,
    \ix_double_ns[34][0] }),
    .south_single({\ix_single_ns[34][3] ,
    \ix_single_ns[34][2] ,
    \ix_single_ns[34][1] ,
    \ix_single_ns[34][0] }),
    .west_double({\ix_double_ew[38][7] ,
    \ix_double_ew[38][6] ,
    \ix_double_ew[38][5] ,
    \ix_double_ew[38][4] ,
    \ix_double_ew[38][3] ,
    \ix_double_ew[38][2] ,
    \ix_double_ew[38][1] ,
    \ix_double_ew[38][0] }),
    .west_single({\ix_single_ew[38][3] ,
    \ix_single_ew[38][2] ,
    \ix_single_ew[38][1] ,
    \ix_single_ew[38][0] }));
 clb_tile \X[6].Y[5].clb  (.carry_in(\carry[5][6] ),
    .carry_out(\carry[6][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[5][6] ),
    .set_out_hard(\col_set[6][6] ),
    .shift_in_hard(\col_shift[5][6] ),
    .shift_out_hard(\col_shift[6][6] ),
    .cb_east_in({_216_,
    _215_,
    _214_,
    _213_,
    _212_}),
    .cb_east_out({\dc_we[47][9] ,
    \dc_we[47][8] ,
    \dc_we[47][7] ,
    \dc_we[47][6] ,
    \dc_we[47][5] ,
    \dc_we[47][4] ,
    \dc_we[47][3] ,
    \dc_we[47][2] ,
    \dc_we[47][1] ,
    \dc_we[47][0] }),
    .cb_north_in({\dc_ns[48][4] ,
    \dc_ns[48][3] ,
    \dc_ns[48][2] ,
    \dc_ns[48][1] ,
    \dc_ns[48][0] }),
    .cb_north_out({\dc_sn[48][9] ,
    \dc_sn[48][8] ,
    \dc_sn[48][7] ,
    \dc_sn[48][6] ,
    \dc_sn[48][5] ,
    \dc_sn[48][4] ,
    \dc_sn[48][3] ,
    \dc_sn[48][2] ,
    \dc_sn[48][1] ,
    \dc_sn[48][0] }),
    .clb_south_in({\dc_sn[41][9] ,
    \dc_sn[41][8] ,
    \dc_sn[41][7] ,
    \dc_sn[41][6] ,
    \dc_sn[41][5] ,
    \dc_sn[41][4] ,
    \dc_sn[41][3] ,
    \dc_sn[41][2] ,
    \dc_sn[41][1] ,
    \dc_sn[41][0] }),
    .clb_south_out({\dc_ns[41][4] ,
    \dc_ns[41][3] ,
    \dc_ns[41][2] ,
    \dc_ns[41][1] ,
    \dc_ns[41][0] }),
    .clb_west_in({\dc_we[46][9] ,
    \dc_we[46][8] ,
    \dc_we[46][7] ,
    \dc_we[46][6] ,
    \dc_we[46][5] ,
    \dc_we[46][4] ,
    \dc_we[46][3] ,
    \dc_we[46][2] ,
    \dc_we[46][1] ,
    \dc_we[46][0] }),
    .clb_west_out({\dc_ew[46][4] ,
    \dc_ew[46][3] ,
    \dc_ew[46][2] ,
    \dc_ew[46][1] ,
    \dc_ew[46][0] }),
    .east_double({\ix_double_ew[47][7] ,
    \ix_double_ew[47][6] ,
    \ix_double_ew[47][5] ,
    \ix_double_ew[47][4] ,
    \ix_double_ew[47][3] ,
    \ix_double_ew[47][2] ,
    \ix_double_ew[47][1] ,
    \ix_double_ew[47][0] }),
    .east_single({\ix_single_ew[47][3] ,
    \ix_single_ew[47][2] ,
    \ix_single_ew[47][1] ,
    gpio_east[5]}),
    .north_double({\ix_double_ns[48][7] ,
    \ix_double_ns[48][6] ,
    \ix_double_ns[48][5] ,
    \ix_double_ns[48][4] ,
    \ix_double_ns[48][3] ,
    \ix_double_ns[48][2] ,
    \ix_double_ns[48][1] ,
    \ix_double_ns[48][0] }),
    .north_single({\ix_single_ns[48][3] ,
    \ix_single_ns[48][2] ,
    \ix_single_ns[48][1] ,
    \ix_single_ns[48][0] }),
    .south_double({\ix_double_ns[41][7] ,
    \ix_double_ns[41][6] ,
    \ix_double_ns[41][5] ,
    \ix_double_ns[41][4] ,
    \ix_double_ns[41][3] ,
    \ix_double_ns[41][2] ,
    \ix_double_ns[41][1] ,
    \ix_double_ns[41][0] }),
    .south_single({\ix_single_ns[41][3] ,
    \ix_single_ns[41][2] ,
    \ix_single_ns[41][1] ,
    \ix_single_ns[41][0] }),
    .west_double({\ix_double_ew[46][7] ,
    \ix_double_ew[46][6] ,
    \ix_double_ew[46][5] ,
    \ix_double_ew[46][4] ,
    \ix_double_ew[46][3] ,
    \ix_double_ew[46][2] ,
    \ix_double_ew[46][1] ,
    \ix_double_ew[46][0] }),
    .west_single({\ix_single_ew[46][3] ,
    \ix_single_ew[46][2] ,
    \ix_single_ew[46][1] ,
    \ix_single_ew[46][0] }));
 clb_tile \X[6].Y[6].clb  (.carry_in(\carry[6][6] ),
    .carry_out(\carry[7][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[6][6] ),
    .set_out_hard(\col_set[7][6] ),
    .shift_in_hard(\col_shift[6][6] ),
    .shift_out_hard(\col_shift[7][6] ),
    .cb_east_in({_221_,
    _220_,
    _219_,
    _218_,
    _217_}),
    .cb_east_out({\dc_we[55][9] ,
    \dc_we[55][8] ,
    \dc_we[55][7] ,
    \dc_we[55][6] ,
    \dc_we[55][5] ,
    \dc_we[55][4] ,
    \dc_we[55][3] ,
    \dc_we[55][2] ,
    \dc_we[55][1] ,
    \dc_we[55][0] }),
    .cb_north_in({\dc_ns[55][4] ,
    \dc_ns[55][3] ,
    \dc_ns[55][2] ,
    \dc_ns[55][1] ,
    \dc_ns[55][0] }),
    .cb_north_out({\dc_sn[55][9] ,
    \dc_sn[55][8] ,
    \dc_sn[55][7] ,
    \dc_sn[55][6] ,
    \dc_sn[55][5] ,
    \dc_sn[55][4] ,
    \dc_sn[55][3] ,
    \dc_sn[55][2] ,
    \dc_sn[55][1] ,
    \dc_sn[55][0] }),
    .clb_south_in({\dc_sn[48][9] ,
    \dc_sn[48][8] ,
    \dc_sn[48][7] ,
    \dc_sn[48][6] ,
    \dc_sn[48][5] ,
    \dc_sn[48][4] ,
    \dc_sn[48][3] ,
    \dc_sn[48][2] ,
    \dc_sn[48][1] ,
    \dc_sn[48][0] }),
    .clb_south_out({\dc_ns[48][4] ,
    \dc_ns[48][3] ,
    \dc_ns[48][2] ,
    \dc_ns[48][1] ,
    \dc_ns[48][0] }),
    .clb_west_in({\dc_we[54][9] ,
    \dc_we[54][8] ,
    \dc_we[54][7] ,
    \dc_we[54][6] ,
    \dc_we[54][5] ,
    \dc_we[54][4] ,
    \dc_we[54][3] ,
    \dc_we[54][2] ,
    \dc_we[54][1] ,
    \dc_we[54][0] }),
    .clb_west_out({\dc_ew[54][4] ,
    \dc_ew[54][3] ,
    \dc_ew[54][2] ,
    \dc_ew[54][1] ,
    \dc_ew[54][0] }),
    .east_double({\ix_double_ew[55][7] ,
    \ix_double_ew[55][6] ,
    \ix_double_ew[55][5] ,
    \ix_double_ew[55][4] ,
    \ix_double_ew[55][3] ,
    \ix_double_ew[55][2] ,
    \ix_double_ew[55][1] ,
    \ix_double_ew[55][0] }),
    .east_single({\ix_single_ew[55][3] ,
    \ix_single_ew[55][2] ,
    \ix_single_ew[55][1] ,
    gpio_east[6]}),
    .north_double({\ix_double_ns[55][7] ,
    \ix_double_ns[55][6] ,
    \ix_double_ns[55][5] ,
    \ix_double_ns[55][4] ,
    \ix_double_ns[55][3] ,
    \ix_double_ns[55][2] ,
    \ix_double_ns[55][1] ,
    \ix_double_ns[55][0] }),
    .north_single({\ix_single_ns[55][3] ,
    \ix_single_ns[55][2] ,
    \ix_single_ns[55][1] ,
    \ix_single_ns[55][0] }),
    .south_double({\ix_double_ns[48][7] ,
    \ix_double_ns[48][6] ,
    \ix_double_ns[48][5] ,
    \ix_double_ns[48][4] ,
    \ix_double_ns[48][3] ,
    \ix_double_ns[48][2] ,
    \ix_double_ns[48][1] ,
    \ix_double_ns[48][0] }),
    .south_single({\ix_single_ns[48][3] ,
    \ix_single_ns[48][2] ,
    \ix_single_ns[48][1] ,
    \ix_single_ns[48][0] }),
    .west_double({\ix_double_ew[54][7] ,
    \ix_double_ew[54][6] ,
    \ix_double_ew[54][5] ,
    \ix_double_ew[54][4] ,
    \ix_double_ew[54][3] ,
    \ix_double_ew[54][2] ,
    \ix_double_ew[54][1] ,
    \ix_double_ew[54][0] }),
    .west_single({\ix_single_ew[54][3] ,
    \ix_single_ew[54][2] ,
    \ix_single_ew[54][1] ,
    \ix_single_ew[54][0] }));
 clb_tile \X[6].Y[7].clb  (.carry_in(\carry[7][6] ),
    .carry_out(\carry[8][6] ),
    .cen(\wb_cen_out[1] ),
    .clk(wb_clk_i),
    .rst(gpio_north[9]),
    .set_in_hard(\col_set[7][6] ),
    .set_out_hard(\col_set[8][6] ),
    .shift_in_hard(\col_shift[7][6] ),
    .shift_out_hard(\col_shift[8][6] ),
    .cb_east_in({_226_,
    _225_,
    _224_,
    _223_,
    _222_}),
    .cb_east_out({\dc_we[63][9] ,
    \dc_we[63][8] ,
    \dc_we[63][7] ,
    \dc_we[63][6] ,
    \dc_we[63][5] ,
    \dc_we[63][4] ,
    \dc_we[63][3] ,
    \dc_we[63][2] ,
    \dc_we[63][1] ,
    \dc_we[63][0] }),
    .cb_north_in({_231_,
    _230_,
    _229_,
    _228_,
    _227_}),
    .cb_north_out({\dc_sn[62][9] ,
    \dc_sn[62][8] ,
    \dc_sn[62][7] ,
    \dc_sn[62][6] ,
    \dc_sn[62][5] ,
    \dc_sn[62][4] ,
    \dc_sn[62][3] ,
    \dc_sn[62][2] ,
    \dc_sn[62][1] ,
    \dc_sn[62][0] }),
    .clb_south_in({\dc_sn[55][9] ,
    \dc_sn[55][8] ,
    \dc_sn[55][7] ,
    \dc_sn[55][6] ,
    \dc_sn[55][5] ,
    \dc_sn[55][4] ,
    \dc_sn[55][3] ,
    \dc_sn[55][2] ,
    \dc_sn[55][1] ,
    \dc_sn[55][0] }),
    .clb_south_out({\dc_ns[55][4] ,
    \dc_ns[55][3] ,
    \dc_ns[55][2] ,
    \dc_ns[55][1] ,
    \dc_ns[55][0] }),
    .clb_west_in({\dc_we[62][9] ,
    \dc_we[62][8] ,
    \dc_we[62][7] ,
    \dc_we[62][6] ,
    \dc_we[62][5] ,
    \dc_we[62][4] ,
    \dc_we[62][3] ,
    \dc_we[62][2] ,
    \dc_we[62][1] ,
    \dc_we[62][0] }),
    .clb_west_out({\dc_ew[62][4] ,
    \dc_ew[62][3] ,
    \dc_ew[62][2] ,
    \dc_ew[62][1] ,
    \dc_ew[62][0] }),
    .east_double({\ix_double_ew[63][7] ,
    \ix_double_ew[63][6] ,
    \ix_double_ew[63][5] ,
    \ix_double_ew[63][4] ,
    \ix_double_ew[63][3] ,
    \ix_double_ew[63][2] ,
    \ix_double_ew[63][1] ,
    \ix_double_ew[63][0] }),
    .east_single({\ix_single_ew[63][3] ,
    \ix_single_ew[63][2] ,
    \ix_single_ew[63][1] ,
    gpio_east[7]}),
    .north_double({\ix_double_ns[62][7] ,
    \ix_double_ns[62][6] ,
    \ix_double_ns[62][5] ,
    \ix_double_ns[62][4] ,
    \ix_double_ns[62][3] ,
    \ix_double_ns[62][2] ,
    \ix_double_ns[62][1] ,
    \ix_double_ns[62][0] }),
    .north_single({\ix_single_ns[62][3] ,
    \ix_single_ns[62][2] ,
    \ix_single_ns[62][1] ,
    gpio_north[6]}),
    .south_double({\ix_double_ns[55][7] ,
    \ix_double_ns[55][6] ,
    \ix_double_ns[55][5] ,
    \ix_double_ns[55][4] ,
    \ix_double_ns[55][3] ,
    \ix_double_ns[55][2] ,
    \ix_double_ns[55][1] ,
    \ix_double_ns[55][0] }),
    .south_single({\ix_single_ns[55][3] ,
    \ix_single_ns[55][2] ,
    \ix_single_ns[55][1] ,
    \ix_single_ns[55][0] }),
    .west_double({\ix_double_ew[62][7] ,
    \ix_double_ew[62][6] ,
    \ix_double_ew[62][5] ,
    \ix_double_ew[62][4] ,
    \ix_double_ew[62][3] ,
    \ix_double_ew[62][2] ,
    \ix_double_ew[62][1] ,
    \ix_double_ew[62][0] }),
    .west_single({\ix_single_ew[62][3] ,
    \ix_single_ew[62][2] ,
    \ix_single_ew[62][1] ,
    \ix_single_ew[62][0] }));
 sky130_fd_sc_hd__or2_4 _232_ (.A(\wbs_data_o_internal[1][0] ),
    .B(\wbs_data_o_internal[0][0] ),
    .X(wbs_data_o[0]));
 sky130_fd_sc_hd__or2_4 _233_ (.A(\wbs_data_o_internal[1][1] ),
    .B(\wbs_data_o_internal[0][1] ),
    .X(wbs_data_o[1]));
 sky130_fd_sc_hd__or2_4 _234_ (.A(\wbs_data_o_internal[1][2] ),
    .B(\wbs_data_o_internal[0][2] ),
    .X(wbs_data_o[2]));
 sky130_fd_sc_hd__or2_4 _235_ (.A(\wbs_data_o_internal[1][3] ),
    .B(\wbs_data_o_internal[0][3] ),
    .X(wbs_data_o[3]));
 sky130_fd_sc_hd__or2_4 _236_ (.A(\wbs_data_o_internal[1][4] ),
    .B(\wbs_data_o_internal[0][4] ),
    .X(wbs_data_o[4]));
 sky130_fd_sc_hd__or2_4 _237_ (.A(\wbs_data_o_internal[1][5] ),
    .B(\wbs_data_o_internal[0][5] ),
    .X(wbs_data_o[5]));
 sky130_fd_sc_hd__or2_4 _238_ (.A(\wbs_data_o_internal[1][6] ),
    .B(\wbs_data_o_internal[0][6] ),
    .X(wbs_data_o[6]));
 sky130_fd_sc_hd__or2_4 _239_ (.A(\wbs_data_o_internal[1][7] ),
    .B(\wbs_data_o_internal[0][7] ),
    .X(wbs_data_o[7]));
 sky130_fd_sc_hd__or2_4 _240_ (.A(\wbs_data_o_internal[1][8] ),
    .B(\wbs_data_o_internal[0][8] ),
    .X(wbs_data_o[8]));
 sky130_fd_sc_hd__or2_4 _241_ (.A(\wbs_data_o_internal[1][9] ),
    .B(\wbs_data_o_internal[0][9] ),
    .X(wbs_data_o[9]));
 sky130_fd_sc_hd__or2_4 _242_ (.A(\wbs_data_o_internal[1][10] ),
    .B(\wbs_data_o_internal[0][10] ),
    .X(wbs_data_o[10]));
 sky130_fd_sc_hd__or2_4 _243_ (.A(\wbs_data_o_internal[1][11] ),
    .B(\wbs_data_o_internal[0][11] ),
    .X(wbs_data_o[11]));
 sky130_fd_sc_hd__or2_4 _244_ (.A(\wbs_data_o_internal[1][12] ),
    .B(\wbs_data_o_internal[0][12] ),
    .X(wbs_data_o[12]));
 sky130_fd_sc_hd__or2_4 _245_ (.A(\wbs_data_o_internal[1][13] ),
    .B(\wbs_data_o_internal[0][13] ),
    .X(wbs_data_o[13]));
 sky130_fd_sc_hd__or2_4 _246_ (.A(\wbs_data_o_internal[1][14] ),
    .B(\wbs_data_o_internal[0][14] ),
    .X(wbs_data_o[14]));
 sky130_fd_sc_hd__or2_4 _247_ (.A(\wbs_data_o_internal[1][15] ),
    .B(\wbs_data_o_internal[0][15] ),
    .X(wbs_data_o[15]));
 sky130_fd_sc_hd__or2_4 _248_ (.A(\wbs_data_o_internal[1][16] ),
    .B(\wbs_data_o_internal[0][16] ),
    .X(wbs_data_o[16]));
 sky130_fd_sc_hd__or2_4 _249_ (.A(\wbs_data_o_internal[1][17] ),
    .B(\wbs_data_o_internal[0][17] ),
    .X(wbs_data_o[17]));
 sky130_fd_sc_hd__or2_4 _250_ (.A(\wbs_data_o_internal[1][18] ),
    .B(\wbs_data_o_internal[0][18] ),
    .X(wbs_data_o[18]));
 sky130_fd_sc_hd__or2_4 _251_ (.A(\wbs_data_o_internal[1][19] ),
    .B(\wbs_data_o_internal[0][19] ),
    .X(wbs_data_o[19]));
 sky130_fd_sc_hd__or2_4 _252_ (.A(\wbs_data_o_internal[1][20] ),
    .B(\wbs_data_o_internal[0][20] ),
    .X(wbs_data_o[20]));
 sky130_fd_sc_hd__or2_4 _253_ (.A(\wbs_data_o_internal[1][21] ),
    .B(\wbs_data_o_internal[0][21] ),
    .X(wbs_data_o[21]));
 sky130_fd_sc_hd__or2_4 _254_ (.A(\wbs_data_o_internal[1][22] ),
    .B(\wbs_data_o_internal[0][22] ),
    .X(wbs_data_o[22]));
 sky130_fd_sc_hd__or2_4 _255_ (.A(\wbs_data_o_internal[1][23] ),
    .B(\wbs_data_o_internal[0][23] ),
    .X(wbs_data_o[23]));
 sky130_fd_sc_hd__or2_4 _256_ (.A(\wbs_data_o_internal[1][24] ),
    .B(\wbs_data_o_internal[0][24] ),
    .X(wbs_data_o[24]));
 sky130_fd_sc_hd__or2_4 _257_ (.A(\wbs_data_o_internal[1][25] ),
    .B(\wbs_data_o_internal[0][25] ),
    .X(wbs_data_o[25]));
 sky130_fd_sc_hd__or2_4 _258_ (.A(\wbs_data_o_internal[1][26] ),
    .B(\wbs_data_o_internal[0][26] ),
    .X(wbs_data_o[26]));
 sky130_fd_sc_hd__or2_4 _259_ (.A(\wbs_data_o_internal[1][27] ),
    .B(\wbs_data_o_internal[0][27] ),
    .X(wbs_data_o[27]));
 sky130_fd_sc_hd__or2_4 _260_ (.A(\wbs_data_o_internal[1][28] ),
    .B(\wbs_data_o_internal[0][28] ),
    .X(wbs_data_o[28]));
 sky130_fd_sc_hd__or2_4 _261_ (.A(\wbs_data_o_internal[1][29] ),
    .B(\wbs_data_o_internal[0][29] ),
    .X(wbs_data_o[29]));
 sky130_fd_sc_hd__or2_4 _262_ (.A(\wbs_data_o_internal[1][30] ),
    .B(\wbs_data_o_internal[0][30] ),
    .X(wbs_data_o[30]));
 sky130_fd_sc_hd__or2_4 _263_ (.A(\wbs_data_o_internal[1][31] ),
    .B(\wbs_data_o_internal[0][31] ),
    .X(wbs_data_o[31]));
 sky130_fd_sc_hd__or2_4 _264_ (.A(\wbs_ack_o_internal[1] ),
    .B(\wbs_ack_o_internal[0] ),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__conb_1 _265_ (.LO(_000_));
 sky130_fd_sc_hd__conb_1 _266_ (.LO(_001_));
 sky130_fd_sc_hd__conb_1 _267_ (.LO(_002_));
 sky130_fd_sc_hd__conb_1 _268_ (.LO(_003_));
 sky130_fd_sc_hd__conb_1 _269_ (.LO(_004_));
 sky130_fd_sc_hd__conb_1 _270_ (.LO(_005_));
 sky130_fd_sc_hd__conb_1 _271_ (.LO(_006_));
 sky130_fd_sc_hd__conb_1 _272_ (.LO(_007_));
 sky130_fd_sc_hd__conb_1 _273_ (.LO(_008_));
 sky130_fd_sc_hd__conb_1 _274_ (.LO(_009_));
 sky130_fd_sc_hd__conb_1 _275_ (.LO(_010_));
 sky130_fd_sc_hd__conb_1 _276_ (.LO(_011_));
 sky130_fd_sc_hd__conb_1 _277_ (.LO(_012_));
 sky130_fd_sc_hd__conb_1 _278_ (.LO(_013_));
 sky130_fd_sc_hd__conb_1 _279_ (.LO(_014_));
 sky130_fd_sc_hd__conb_1 _280_ (.LO(_015_));
 sky130_fd_sc_hd__conb_1 _281_ (.LO(_016_));
 sky130_fd_sc_hd__conb_1 _282_ (.LO(_017_));
 sky130_fd_sc_hd__conb_1 _283_ (.LO(_018_));
 sky130_fd_sc_hd__conb_1 _284_ (.LO(_019_));
 sky130_fd_sc_hd__conb_1 _285_ (.LO(_020_));
 sky130_fd_sc_hd__conb_1 _286_ (.LO(_021_));
 sky130_fd_sc_hd__conb_1 _287_ (.LO(_022_));
 sky130_fd_sc_hd__conb_1 _288_ (.LO(_023_));
 sky130_fd_sc_hd__conb_1 _289_ (.LO(_024_));
 sky130_fd_sc_hd__conb_1 _290_ (.LO(_025_));
 sky130_fd_sc_hd__conb_1 _291_ (.LO(_026_));
 sky130_fd_sc_hd__conb_1 _292_ (.LO(_027_));
 sky130_fd_sc_hd__conb_1 _293_ (.LO(_028_));
 sky130_fd_sc_hd__conb_1 _294_ (.LO(_029_));
 sky130_fd_sc_hd__conb_1 _295_ (.LO(_030_));
 sky130_fd_sc_hd__conb_1 _296_ (.LO(_031_));
 sky130_fd_sc_hd__conb_1 _297_ (.LO(_032_));
 sky130_fd_sc_hd__conb_1 _298_ (.LO(_033_));
 sky130_fd_sc_hd__conb_1 _299_ (.LO(_034_));
 sky130_fd_sc_hd__conb_1 _300_ (.LO(_035_));
 sky130_fd_sc_hd__conb_1 _301_ (.LO(_036_));
 sky130_fd_sc_hd__conb_1 _302_ (.LO(_037_));
 sky130_fd_sc_hd__conb_1 _303_ (.LO(_038_));
 sky130_fd_sc_hd__conb_1 _304_ (.LO(_039_));
 sky130_fd_sc_hd__conb_1 _305_ (.LO(_040_));
 sky130_fd_sc_hd__conb_1 _306_ (.LO(_041_));
 sky130_fd_sc_hd__conb_1 _307_ (.LO(_042_));
 sky130_fd_sc_hd__conb_1 _308_ (.LO(_043_));
 sky130_fd_sc_hd__conb_1 _309_ (.LO(_044_));
 sky130_fd_sc_hd__conb_1 _310_ (.LO(_045_));
 sky130_fd_sc_hd__conb_1 _311_ (.LO(_046_));
 sky130_fd_sc_hd__conb_1 _312_ (.LO(_047_));
 sky130_fd_sc_hd__conb_1 _313_ (.LO(_048_));
 sky130_fd_sc_hd__conb_1 _314_ (.LO(_049_));
 sky130_fd_sc_hd__conb_1 _315_ (.LO(_050_));
 sky130_fd_sc_hd__conb_1 _316_ (.LO(_051_));
 sky130_fd_sc_hd__conb_1 _317_ (.LO(_052_));
 sky130_fd_sc_hd__conb_1 _318_ (.LO(_053_));
 sky130_fd_sc_hd__conb_1 _319_ (.LO(_054_));
 sky130_fd_sc_hd__conb_1 _320_ (.LO(_055_));
 sky130_fd_sc_hd__conb_1 _321_ (.LO(_056_));
 sky130_fd_sc_hd__conb_1 _322_ (.LO(_057_));
 sky130_fd_sc_hd__conb_1 _323_ (.LO(_058_));
 sky130_fd_sc_hd__conb_1 _324_ (.LO(_059_));
 sky130_fd_sc_hd__conb_1 _325_ (.LO(_060_));
 sky130_fd_sc_hd__conb_1 _326_ (.LO(_061_));
 sky130_fd_sc_hd__conb_1 _327_ (.LO(_062_));
 sky130_fd_sc_hd__conb_1 _328_ (.LO(_063_));
 sky130_fd_sc_hd__conb_1 _329_ (.LO(_064_));
 sky130_fd_sc_hd__conb_1 _330_ (.LO(_065_));
 sky130_fd_sc_hd__conb_1 _331_ (.LO(_066_));
 sky130_fd_sc_hd__conb_1 _332_ (.LO(_067_));
 sky130_fd_sc_hd__conb_1 _333_ (.LO(_068_));
 sky130_fd_sc_hd__conb_1 _334_ (.LO(_069_));
 sky130_fd_sc_hd__conb_1 _335_ (.LO(_070_));
 sky130_fd_sc_hd__conb_1 _336_ (.LO(_071_));
 sky130_fd_sc_hd__conb_1 _337_ (.LO(_072_));
 sky130_fd_sc_hd__conb_1 _338_ (.LO(_073_));
 sky130_fd_sc_hd__conb_1 _339_ (.LO(_074_));
 sky130_fd_sc_hd__conb_1 _340_ (.LO(_075_));
 sky130_fd_sc_hd__conb_1 _341_ (.LO(_076_));
 sky130_fd_sc_hd__conb_1 _342_ (.LO(_077_));
 sky130_fd_sc_hd__conb_1 _343_ (.LO(_078_));
 sky130_fd_sc_hd__conb_1 _344_ (.LO(_079_));
 sky130_fd_sc_hd__conb_1 _345_ (.LO(_080_));
 sky130_fd_sc_hd__conb_1 _346_ (.LO(_081_));
 sky130_fd_sc_hd__conb_1 _347_ (.LO(_082_));
 sky130_fd_sc_hd__conb_1 _348_ (.LO(_083_));
 sky130_fd_sc_hd__conb_1 _349_ (.LO(_084_));
 sky130_fd_sc_hd__conb_1 _350_ (.LO(_085_));
 sky130_fd_sc_hd__conb_1 _351_ (.LO(_086_));
 sky130_fd_sc_hd__conb_1 _352_ (.LO(_087_));
 sky130_fd_sc_hd__conb_1 _353_ (.LO(_088_));
 sky130_fd_sc_hd__conb_1 _354_ (.LO(_089_));
 sky130_fd_sc_hd__conb_1 _355_ (.LO(_090_));
 sky130_fd_sc_hd__conb_1 _356_ (.LO(_091_));
 sky130_fd_sc_hd__conb_1 _357_ (.LO(_092_));
 sky130_fd_sc_hd__conb_1 _358_ (.LO(_093_));
 sky130_fd_sc_hd__conb_1 _359_ (.LO(_094_));
 sky130_fd_sc_hd__conb_1 _360_ (.LO(_095_));
 sky130_fd_sc_hd__conb_1 _361_ (.LO(_096_));
 sky130_fd_sc_hd__conb_1 _362_ (.LO(_097_));
 sky130_fd_sc_hd__conb_1 _363_ (.LO(_098_));
 sky130_fd_sc_hd__conb_1 _364_ (.LO(_099_));
 sky130_fd_sc_hd__conb_1 _365_ (.LO(_100_));
 sky130_fd_sc_hd__conb_1 _366_ (.LO(_101_));
 sky130_fd_sc_hd__conb_1 _367_ (.LO(_102_));
 sky130_fd_sc_hd__conb_1 _368_ (.LO(_103_));
 sky130_fd_sc_hd__conb_1 _369_ (.LO(_104_));
 sky130_fd_sc_hd__conb_1 _370_ (.LO(_105_));
 sky130_fd_sc_hd__conb_1 _371_ (.LO(_106_));
 sky130_fd_sc_hd__conb_1 _372_ (.LO(_107_));
 sky130_fd_sc_hd__conb_1 _373_ (.LO(_108_));
 sky130_fd_sc_hd__conb_1 _374_ (.LO(_109_));
 sky130_fd_sc_hd__conb_1 _375_ (.LO(_110_));
 sky130_fd_sc_hd__conb_1 _376_ (.LO(_111_));
 sky130_fd_sc_hd__conb_1 _377_ (.LO(_112_));
 sky130_fd_sc_hd__conb_1 _378_ (.LO(_113_));
 sky130_fd_sc_hd__conb_1 _379_ (.LO(_114_));
 sky130_fd_sc_hd__conb_1 _380_ (.LO(_115_));
 sky130_fd_sc_hd__conb_1 _381_ (.LO(_116_));
 sky130_fd_sc_hd__conb_1 _382_ (.LO(_117_));
 sky130_fd_sc_hd__conb_1 _383_ (.LO(_118_));
 sky130_fd_sc_hd__conb_1 _384_ (.LO(_119_));
 sky130_fd_sc_hd__conb_1 _385_ (.LO(_120_));
 sky130_fd_sc_hd__conb_1 _386_ (.LO(_121_));
 sky130_fd_sc_hd__conb_1 _387_ (.LO(_122_));
 sky130_fd_sc_hd__conb_1 _388_ (.LO(_123_));
 sky130_fd_sc_hd__conb_1 _389_ (.LO(_124_));
 sky130_fd_sc_hd__conb_1 _390_ (.LO(_125_));
 sky130_fd_sc_hd__conb_1 _391_ (.LO(_126_));
 sky130_fd_sc_hd__conb_1 _392_ (.LO(_127_));
 sky130_fd_sc_hd__conb_1 _393_ (.LO(_128_));
 sky130_fd_sc_hd__conb_1 _394_ (.LO(_129_));
 sky130_fd_sc_hd__conb_1 _395_ (.LO(_130_));
 sky130_fd_sc_hd__conb_1 _396_ (.LO(_131_));
 sky130_fd_sc_hd__conb_1 _397_ (.LO(_132_));
 sky130_fd_sc_hd__conb_1 _398_ (.LO(_133_));
 sky130_fd_sc_hd__conb_1 _399_ (.LO(_134_));
 sky130_fd_sc_hd__conb_1 _400_ (.LO(_135_));
 sky130_fd_sc_hd__conb_1 _401_ (.LO(_136_));
 sky130_fd_sc_hd__conb_1 _402_ (.LO(_137_));
 sky130_fd_sc_hd__conb_1 _403_ (.LO(_138_));
 sky130_fd_sc_hd__conb_1 _404_ (.LO(_139_));
 sky130_fd_sc_hd__conb_1 _405_ (.LO(_140_));
 sky130_fd_sc_hd__conb_1 _406_ (.LO(_141_));
 sky130_fd_sc_hd__conb_1 _407_ (.LO(_142_));
 sky130_fd_sc_hd__conb_1 _408_ (.LO(_143_));
 sky130_fd_sc_hd__conb_1 _409_ (.LO(_144_));
 sky130_fd_sc_hd__conb_1 _410_ (.LO(_145_));
 sky130_fd_sc_hd__conb_1 _411_ (.LO(_146_));
 sky130_fd_sc_hd__conb_1 _412_ (.LO(_147_));
 sky130_fd_sc_hd__conb_1 _413_ (.LO(_148_));
 sky130_fd_sc_hd__conb_1 _414_ (.LO(_149_));
 sky130_fd_sc_hd__conb_1 _415_ (.LO(_150_));
 sky130_fd_sc_hd__conb_1 _416_ (.LO(_151_));
 sky130_fd_sc_hd__conb_1 _417_ (.LO(_152_));
 sky130_fd_sc_hd__conb_1 _418_ (.LO(_153_));
 sky130_fd_sc_hd__conb_1 _419_ (.LO(_154_));
 sky130_fd_sc_hd__conb_1 _420_ (.LO(_155_));
 sky130_fd_sc_hd__conb_1 _421_ (.LO(_156_));
 sky130_fd_sc_hd__conb_1 _422_ (.LO(_157_));
 sky130_fd_sc_hd__conb_1 _423_ (.LO(_158_));
 sky130_fd_sc_hd__conb_1 _424_ (.LO(_159_));
 sky130_fd_sc_hd__conb_1 _425_ (.LO(_160_));
 sky130_fd_sc_hd__conb_1 _426_ (.LO(_161_));
 sky130_fd_sc_hd__conb_1 _427_ (.LO(_162_));
 sky130_fd_sc_hd__conb_1 _428_ (.LO(_163_));
 sky130_fd_sc_hd__conb_1 _429_ (.LO(_164_));
 sky130_fd_sc_hd__conb_1 _430_ (.LO(_165_));
 sky130_fd_sc_hd__conb_1 _431_ (.LO(_166_));
 sky130_fd_sc_hd__conb_1 _432_ (.LO(_167_));
 sky130_fd_sc_hd__conb_1 _433_ (.LO(_168_));
 sky130_fd_sc_hd__conb_1 _434_ (.LO(_169_));
 sky130_fd_sc_hd__conb_1 _435_ (.LO(_170_));
 sky130_fd_sc_hd__conb_1 _436_ (.LO(_171_));
 sky130_fd_sc_hd__conb_1 _437_ (.LO(_172_));
 sky130_fd_sc_hd__conb_1 _438_ (.LO(_173_));
 sky130_fd_sc_hd__conb_1 _439_ (.LO(_174_));
 sky130_fd_sc_hd__conb_1 _440_ (.LO(_175_));
 sky130_fd_sc_hd__conb_1 _441_ (.LO(_176_));
 sky130_fd_sc_hd__conb_1 _442_ (.LO(_177_));
 sky130_fd_sc_hd__conb_1 _443_ (.LO(_178_));
 sky130_fd_sc_hd__conb_1 _444_ (.LO(_179_));
 sky130_fd_sc_hd__conb_1 _445_ (.LO(_180_));
 sky130_fd_sc_hd__conb_1 _446_ (.LO(_181_));
 sky130_fd_sc_hd__conb_1 _447_ (.LO(_182_));
 sky130_fd_sc_hd__conb_1 _448_ (.LO(_183_));
 sky130_fd_sc_hd__conb_1 _449_ (.LO(_184_));
 sky130_fd_sc_hd__conb_1 _450_ (.LO(_185_));
 sky130_fd_sc_hd__conb_1 _451_ (.LO(_186_));
 sky130_fd_sc_hd__conb_1 _452_ (.LO(_187_));
 sky130_fd_sc_hd__conb_1 _453_ (.LO(_188_));
 sky130_fd_sc_hd__conb_1 _454_ (.LO(_189_));
 sky130_fd_sc_hd__conb_1 _455_ (.LO(_190_));
 sky130_fd_sc_hd__conb_1 _456_ (.LO(_191_));
 sky130_fd_sc_hd__conb_1 _457_ (.LO(_192_));
 sky130_fd_sc_hd__conb_1 _458_ (.LO(_193_));
 sky130_fd_sc_hd__conb_1 _459_ (.LO(_194_));
 sky130_fd_sc_hd__conb_1 _460_ (.LO(_195_));
 sky130_fd_sc_hd__conb_1 _461_ (.LO(_196_));
 sky130_fd_sc_hd__conb_1 _462_ (.LO(_197_));
 sky130_fd_sc_hd__conb_1 _463_ (.LO(_198_));
 sky130_fd_sc_hd__conb_1 _464_ (.LO(_199_));
 sky130_fd_sc_hd__conb_1 _465_ (.LO(_200_));
 sky130_fd_sc_hd__conb_1 _466_ (.LO(_201_));
 sky130_fd_sc_hd__conb_1 _467_ (.LO(_202_));
 sky130_fd_sc_hd__conb_1 _468_ (.LO(_203_));
 sky130_fd_sc_hd__conb_1 _469_ (.LO(_204_));
 sky130_fd_sc_hd__conb_1 _470_ (.LO(_205_));
 sky130_fd_sc_hd__conb_1 _471_ (.LO(_206_));
 sky130_fd_sc_hd__conb_1 _472_ (.LO(_207_));
 sky130_fd_sc_hd__conb_1 _473_ (.LO(_208_));
 sky130_fd_sc_hd__conb_1 _474_ (.LO(_209_));
 sky130_fd_sc_hd__conb_1 _475_ (.LO(_210_));
 sky130_fd_sc_hd__conb_1 _476_ (.LO(_211_));
 sky130_fd_sc_hd__conb_1 _477_ (.LO(_212_));
 sky130_fd_sc_hd__conb_1 _478_ (.LO(_213_));
 sky130_fd_sc_hd__conb_1 _479_ (.LO(_214_));
 sky130_fd_sc_hd__conb_1 _480_ (.LO(_215_));
 sky130_fd_sc_hd__conb_1 _481_ (.LO(_216_));
 sky130_fd_sc_hd__conb_1 _482_ (.LO(_217_));
 sky130_fd_sc_hd__conb_1 _483_ (.LO(_218_));
 sky130_fd_sc_hd__conb_1 _484_ (.LO(_219_));
 sky130_fd_sc_hd__conb_1 _485_ (.LO(_220_));
 sky130_fd_sc_hd__conb_1 _486_ (.LO(_221_));
 sky130_fd_sc_hd__conb_1 _487_ (.LO(_222_));
 sky130_fd_sc_hd__conb_1 _488_ (.LO(_223_));
 sky130_fd_sc_hd__conb_1 _489_ (.LO(_224_));
 sky130_fd_sc_hd__conb_1 _490_ (.LO(_225_));
 sky130_fd_sc_hd__conb_1 _491_ (.LO(_226_));
 sky130_fd_sc_hd__conb_1 _492_ (.LO(_227_));
 sky130_fd_sc_hd__conb_1 _493_ (.LO(_228_));
 sky130_fd_sc_hd__conb_1 _494_ (.LO(_229_));
 sky130_fd_sc_hd__conb_1 _495_ (.LO(_230_));
 sky130_fd_sc_hd__conb_1 _496_ (.LO(_231_));
 wishbone_configuratorinator_00 wishbonatron_00 (.cen(\wb_cen_out[0] ),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(\wbs_ack_o_internal[0] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .set_out({\wb_set_out[0][3] ,
    \wb_set_out[0][2] ,
    \wb_set_out[0][1] ,
    \wb_set_out[0][0] }),
    .shift_out({\wb_shift_out[0][3] ,
    \wb_shift_out[0][2] ,
    \wb_shift_out[0][1] ,
    \wb_shift_out[0][0] }),
    .wbs_addr_i({wbs_addr_i[31],
    wbs_addr_i[30],
    wbs_addr_i[29],
    wbs_addr_i[28],
    wbs_addr_i[27],
    wbs_addr_i[26],
    wbs_addr_i[25],
    wbs_addr_i[24],
    wbs_addr_i[23],
    wbs_addr_i[22],
    wbs_addr_i[21],
    wbs_addr_i[20],
    wbs_addr_i[19],
    wbs_addr_i[18],
    wbs_addr_i[17],
    wbs_addr_i[16],
    wbs_addr_i[15],
    wbs_addr_i[14],
    wbs_addr_i[13],
    wbs_addr_i[12],
    wbs_addr_i[11],
    wbs_addr_i[10],
    wbs_addr_i[9],
    wbs_addr_i[8],
    wbs_addr_i[7],
    wbs_addr_i[6],
    wbs_addr_i[5],
    wbs_addr_i[4],
    wbs_addr_i[3],
    wbs_addr_i[2],
    wbs_addr_i[1],
    wbs_addr_i[0]}),
    .wbs_data_i({wbs_data_i[31],
    wbs_data_i[30],
    wbs_data_i[29],
    wbs_data_i[28],
    wbs_data_i[27],
    wbs_data_i[26],
    wbs_data_i[25],
    wbs_data_i[24],
    wbs_data_i[23],
    wbs_data_i[22],
    wbs_data_i[21],
    wbs_data_i[20],
    wbs_data_i[19],
    wbs_data_i[18],
    wbs_data_i[17],
    wbs_data_i[16],
    wbs_data_i[15],
    wbs_data_i[14],
    wbs_data_i[13],
    wbs_data_i[12],
    wbs_data_i[11],
    wbs_data_i[10],
    wbs_data_i[9],
    wbs_data_i[8],
    wbs_data_i[7],
    wbs_data_i[6],
    wbs_data_i[5],
    wbs_data_i[4],
    wbs_data_i[3],
    wbs_data_i[2],
    wbs_data_i[1],
    wbs_data_i[0]}),
    .wbs_data_o({\wbs_data_o_internal[0][31] ,
    \wbs_data_o_internal[0][30] ,
    \wbs_data_o_internal[0][29] ,
    \wbs_data_o_internal[0][28] ,
    \wbs_data_o_internal[0][27] ,
    \wbs_data_o_internal[0][26] ,
    \wbs_data_o_internal[0][25] ,
    \wbs_data_o_internal[0][24] ,
    \wbs_data_o_internal[0][23] ,
    \wbs_data_o_internal[0][22] ,
    \wbs_data_o_internal[0][21] ,
    \wbs_data_o_internal[0][20] ,
    \wbs_data_o_internal[0][19] ,
    \wbs_data_o_internal[0][18] ,
    \wbs_data_o_internal[0][17] ,
    \wbs_data_o_internal[0][16] ,
    \wbs_data_o_internal[0][15] ,
    \wbs_data_o_internal[0][14] ,
    \wbs_data_o_internal[0][13] ,
    \wbs_data_o_internal[0][12] ,
    \wbs_data_o_internal[0][11] ,
    \wbs_data_o_internal[0][10] ,
    \wbs_data_o_internal[0][9] ,
    \wbs_data_o_internal[0][8] ,
    \wbs_data_o_internal[0][7] ,
    \wbs_data_o_internal[0][6] ,
    \wbs_data_o_internal[0][5] ,
    \wbs_data_o_internal[0][4] ,
    \wbs_data_o_internal[0][3] ,
    \wbs_data_o_internal[0][2] ,
    \wbs_data_o_internal[0][1] ,
    \wbs_data_o_internal[0][0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 wishbone_configuratorinator_10 wishbonatron_10 (.cen(\wb_cen_out[1] ),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(\wbs_ack_o_internal[1] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .set_out({\wb_set_out[1][3] ,
    \wb_set_out[1][2] ,
    \wb_set_out[1][1] ,
    \wb_set_out[1][0] }),
    .shift_out({\wb_shift_out[1][3] ,
    \wb_shift_out[1][2] ,
    \wb_shift_out[1][1] ,
    \wb_shift_out[1][0] }),
    .wbs_addr_i({wbs_addr_i[31],
    wbs_addr_i[30],
    wbs_addr_i[29],
    wbs_addr_i[28],
    wbs_addr_i[27],
    wbs_addr_i[26],
    wbs_addr_i[25],
    wbs_addr_i[24],
    wbs_addr_i[23],
    wbs_addr_i[22],
    wbs_addr_i[21],
    wbs_addr_i[20],
    wbs_addr_i[19],
    wbs_addr_i[18],
    wbs_addr_i[17],
    wbs_addr_i[16],
    wbs_addr_i[15],
    wbs_addr_i[14],
    wbs_addr_i[13],
    wbs_addr_i[12],
    wbs_addr_i[11],
    wbs_addr_i[10],
    wbs_addr_i[9],
    wbs_addr_i[8],
    wbs_addr_i[7],
    wbs_addr_i[6],
    wbs_addr_i[5],
    wbs_addr_i[4],
    wbs_addr_i[3],
    wbs_addr_i[2],
    wbs_addr_i[1],
    wbs_addr_i[0]}),
    .wbs_data_i({wbs_data_i[31],
    wbs_data_i[30],
    wbs_data_i[29],
    wbs_data_i[28],
    wbs_data_i[27],
    wbs_data_i[26],
    wbs_data_i[25],
    wbs_data_i[24],
    wbs_data_i[23],
    wbs_data_i[22],
    wbs_data_i[21],
    wbs_data_i[20],
    wbs_data_i[19],
    wbs_data_i[18],
    wbs_data_i[17],
    wbs_data_i[16],
    wbs_data_i[15],
    wbs_data_i[14],
    wbs_data_i[13],
    wbs_data_i[12],
    wbs_data_i[11],
    wbs_data_i[10],
    wbs_data_i[9],
    wbs_data_i[8],
    wbs_data_i[7],
    wbs_data_i[6],
    wbs_data_i[5],
    wbs_data_i[4],
    wbs_data_i[3],
    wbs_data_i[2],
    wbs_data_i[1],
    wbs_data_i[0]}),
    .wbs_data_o({\wbs_data_o_internal[1][31] ,
    \wbs_data_o_internal[1][30] ,
    \wbs_data_o_internal[1][29] ,
    \wbs_data_o_internal[1][28] ,
    \wbs_data_o_internal[1][27] ,
    \wbs_data_o_internal[1][26] ,
    \wbs_data_o_internal[1][25] ,
    \wbs_data_o_internal[1][24] ,
    \wbs_data_o_internal[1][23] ,
    \wbs_data_o_internal[1][22] ,
    \wbs_data_o_internal[1][21] ,
    \wbs_data_o_internal[1][20] ,
    \wbs_data_o_internal[1][19] ,
    \wbs_data_o_internal[1][18] ,
    \wbs_data_o_internal[1][17] ,
    \wbs_data_o_internal[1][16] ,
    \wbs_data_o_internal[1][15] ,
    \wbs_data_o_internal[1][14] ,
    \wbs_data_o_internal[1][13] ,
    \wbs_data_o_internal[1][12] ,
    \wbs_data_o_internal[1][11] ,
    \wbs_data_o_internal[1][10] ,
    \wbs_data_o_internal[1][9] ,
    \wbs_data_o_internal[1][8] ,
    \wbs_data_o_internal[1][7] ,
    \wbs_data_o_internal[1][6] ,
    \wbs_data_o_internal[1][5] ,
    \wbs_data_o_internal[1][4] ,
    \wbs_data_o_internal[1][3] ,
    \wbs_data_o_internal[1][2] ,
    \wbs_data_o_internal[1][1] ,
    \wbs_data_o_internal[1][0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_1306 ();
 sky130_fd_sc_hd__decap_3 PHY_1307 ();
 sky130_fd_sc_hd__decap_3 PHY_1308 ();
 sky130_fd_sc_hd__decap_3 PHY_1309 ();
 sky130_fd_sc_hd__decap_3 PHY_1310 ();
 sky130_fd_sc_hd__decap_3 PHY_1311 ();
 sky130_fd_sc_hd__decap_3 PHY_1312 ();
 sky130_fd_sc_hd__decap_3 PHY_1313 ();
 sky130_fd_sc_hd__decap_3 PHY_1314 ();
 sky130_fd_sc_hd__decap_3 PHY_1315 ();
 sky130_fd_sc_hd__decap_3 PHY_1316 ();
 sky130_fd_sc_hd__decap_3 PHY_1317 ();
 sky130_fd_sc_hd__decap_3 PHY_1318 ();
 sky130_fd_sc_hd__decap_3 PHY_1319 ();
 sky130_fd_sc_hd__decap_3 PHY_1320 ();
 sky130_fd_sc_hd__decap_3 PHY_1321 ();
 sky130_fd_sc_hd__decap_3 PHY_1322 ();
 sky130_fd_sc_hd__decap_3 PHY_1323 ();
 sky130_fd_sc_hd__decap_3 PHY_1324 ();
 sky130_fd_sc_hd__decap_3 PHY_1325 ();
 sky130_fd_sc_hd__decap_3 PHY_1326 ();
 sky130_fd_sc_hd__decap_3 PHY_1327 ();
 sky130_fd_sc_hd__decap_3 PHY_1328 ();
 sky130_fd_sc_hd__decap_3 PHY_1329 ();
 sky130_fd_sc_hd__decap_3 PHY_1330 ();
 sky130_fd_sc_hd__decap_3 PHY_1331 ();
 sky130_fd_sc_hd__decap_3 PHY_1332 ();
 sky130_fd_sc_hd__decap_3 PHY_1333 ();
 sky130_fd_sc_hd__decap_3 PHY_1334 ();
 sky130_fd_sc_hd__decap_3 PHY_1335 ();
 sky130_fd_sc_hd__decap_3 PHY_1336 ();
 sky130_fd_sc_hd__decap_3 PHY_1337 ();
 sky130_fd_sc_hd__decap_3 PHY_1338 ();
 sky130_fd_sc_hd__decap_3 PHY_1339 ();
 sky130_fd_sc_hd__decap_3 PHY_1340 ();
 sky130_fd_sc_hd__decap_3 PHY_1341 ();
 sky130_fd_sc_hd__decap_3 PHY_1342 ();
 sky130_fd_sc_hd__decap_3 PHY_1343 ();
 sky130_fd_sc_hd__decap_3 PHY_1344 ();
 sky130_fd_sc_hd__decap_3 PHY_1345 ();
 sky130_fd_sc_hd__decap_3 PHY_1346 ();
 sky130_fd_sc_hd__decap_3 PHY_1347 ();
 sky130_fd_sc_hd__decap_3 PHY_1348 ();
 sky130_fd_sc_hd__decap_3 PHY_1349 ();
 sky130_fd_sc_hd__decap_3 PHY_1350 ();
 sky130_fd_sc_hd__decap_3 PHY_1351 ();
 sky130_fd_sc_hd__decap_3 PHY_1352 ();
 sky130_fd_sc_hd__decap_3 PHY_1353 ();
 sky130_fd_sc_hd__decap_3 PHY_1354 ();
 sky130_fd_sc_hd__decap_3 PHY_1355 ();
 sky130_fd_sc_hd__decap_3 PHY_1356 ();
 sky130_fd_sc_hd__decap_3 PHY_1357 ();
 sky130_fd_sc_hd__decap_3 PHY_1358 ();
 sky130_fd_sc_hd__decap_3 PHY_1359 ();
 sky130_fd_sc_hd__decap_3 PHY_1360 ();
 sky130_fd_sc_hd__decap_3 PHY_1361 ();
 sky130_fd_sc_hd__decap_3 PHY_1362 ();
 sky130_fd_sc_hd__decap_3 PHY_1363 ();
 sky130_fd_sc_hd__decap_3 PHY_1364 ();
 sky130_fd_sc_hd__decap_3 PHY_1365 ();
 sky130_fd_sc_hd__decap_3 PHY_1366 ();
 sky130_fd_sc_hd__decap_3 PHY_1367 ();
 sky130_fd_sc_hd__decap_3 PHY_1368 ();
 sky130_fd_sc_hd__decap_3 PHY_1369 ();
 sky130_fd_sc_hd__decap_3 PHY_1370 ();
 sky130_fd_sc_hd__decap_3 PHY_1371 ();
 sky130_fd_sc_hd__decap_3 PHY_1372 ();
 sky130_fd_sc_hd__decap_3 PHY_1373 ();
 sky130_fd_sc_hd__decap_3 PHY_1374 ();
 sky130_fd_sc_hd__decap_3 PHY_1375 ();
 sky130_fd_sc_hd__decap_3 PHY_1376 ();
 sky130_fd_sc_hd__decap_3 PHY_1377 ();
 sky130_fd_sc_hd__decap_3 PHY_1378 ();
 sky130_fd_sc_hd__decap_3 PHY_1379 ();
 sky130_fd_sc_hd__decap_3 PHY_1380 ();
 sky130_fd_sc_hd__decap_3 PHY_1381 ();
 sky130_fd_sc_hd__decap_3 PHY_1382 ();
 sky130_fd_sc_hd__decap_3 PHY_1383 ();
 sky130_fd_sc_hd__decap_3 PHY_1384 ();
 sky130_fd_sc_hd__decap_3 PHY_1385 ();
 sky130_fd_sc_hd__decap_3 PHY_1386 ();
 sky130_fd_sc_hd__decap_3 PHY_1387 ();
 sky130_fd_sc_hd__decap_3 PHY_1388 ();
 sky130_fd_sc_hd__decap_3 PHY_1389 ();
 sky130_fd_sc_hd__decap_3 PHY_1390 ();
 sky130_fd_sc_hd__decap_3 PHY_1391 ();
 sky130_fd_sc_hd__decap_3 PHY_1392 ();
 sky130_fd_sc_hd__decap_3 PHY_1393 ();
 sky130_fd_sc_hd__decap_3 PHY_1394 ();
 sky130_fd_sc_hd__decap_3 PHY_1395 ();
 sky130_fd_sc_hd__decap_3 PHY_1396 ();
 sky130_fd_sc_hd__decap_3 PHY_1397 ();
 sky130_fd_sc_hd__decap_3 PHY_1398 ();
 sky130_fd_sc_hd__decap_3 PHY_1399 ();
 sky130_fd_sc_hd__decap_3 PHY_1400 ();
 sky130_fd_sc_hd__decap_3 PHY_1401 ();
 sky130_fd_sc_hd__decap_3 PHY_1402 ();
 sky130_fd_sc_hd__decap_3 PHY_1403 ();
 sky130_fd_sc_hd__decap_3 PHY_1404 ();
 sky130_fd_sc_hd__decap_3 PHY_1405 ();
 sky130_fd_sc_hd__decap_3 PHY_1406 ();
 sky130_fd_sc_hd__decap_3 PHY_1407 ();
 sky130_fd_sc_hd__decap_3 PHY_1408 ();
 sky130_fd_sc_hd__decap_3 PHY_1409 ();
 sky130_fd_sc_hd__decap_3 PHY_1410 ();
 sky130_fd_sc_hd__decap_3 PHY_1411 ();
 sky130_fd_sc_hd__decap_3 PHY_1412 ();
 sky130_fd_sc_hd__decap_3 PHY_1413 ();
 sky130_fd_sc_hd__decap_3 PHY_1414 ();
 sky130_fd_sc_hd__decap_3 PHY_1415 ();
 sky130_fd_sc_hd__decap_3 PHY_1416 ();
 sky130_fd_sc_hd__decap_3 PHY_1417 ();
 sky130_fd_sc_hd__decap_3 PHY_1418 ();
 sky130_fd_sc_hd__decap_3 PHY_1419 ();
 sky130_fd_sc_hd__decap_3 PHY_1420 ();
 sky130_fd_sc_hd__decap_3 PHY_1421 ();
 sky130_fd_sc_hd__decap_3 PHY_1422 ();
 sky130_fd_sc_hd__decap_3 PHY_1423 ();
 sky130_fd_sc_hd__decap_3 PHY_1424 ();
 sky130_fd_sc_hd__decap_3 PHY_1425 ();
 sky130_fd_sc_hd__decap_3 PHY_1426 ();
 sky130_fd_sc_hd__decap_3 PHY_1427 ();
 sky130_fd_sc_hd__decap_3 PHY_1428 ();
 sky130_fd_sc_hd__decap_3 PHY_1429 ();
 sky130_fd_sc_hd__decap_3 PHY_1430 ();
 sky130_fd_sc_hd__decap_3 PHY_1431 ();
 sky130_fd_sc_hd__decap_3 PHY_1432 ();
 sky130_fd_sc_hd__decap_3 PHY_1433 ();
 sky130_fd_sc_hd__decap_3 PHY_1434 ();
 sky130_fd_sc_hd__decap_3 PHY_1435 ();
 sky130_fd_sc_hd__decap_3 PHY_1436 ();
 sky130_fd_sc_hd__decap_3 PHY_1437 ();
 sky130_fd_sc_hd__decap_3 PHY_1438 ();
 sky130_fd_sc_hd__decap_3 PHY_1439 ();
 sky130_fd_sc_hd__decap_3 PHY_1440 ();
 sky130_fd_sc_hd__decap_3 PHY_1441 ();
 sky130_fd_sc_hd__decap_3 PHY_1442 ();
 sky130_fd_sc_hd__decap_3 PHY_1443 ();
 sky130_fd_sc_hd__decap_3 PHY_1444 ();
 sky130_fd_sc_hd__decap_3 PHY_1445 ();
 sky130_fd_sc_hd__decap_3 PHY_1446 ();
 sky130_fd_sc_hd__decap_3 PHY_1447 ();
 sky130_fd_sc_hd__decap_3 PHY_1448 ();
 sky130_fd_sc_hd__decap_3 PHY_1449 ();
 sky130_fd_sc_hd__decap_3 PHY_1450 ();
 sky130_fd_sc_hd__decap_3 PHY_1451 ();
 sky130_fd_sc_hd__decap_3 PHY_1452 ();
 sky130_fd_sc_hd__decap_3 PHY_1453 ();
 sky130_fd_sc_hd__decap_3 PHY_1454 ();
 sky130_fd_sc_hd__decap_3 PHY_1455 ();
 sky130_fd_sc_hd__decap_3 PHY_1456 ();
 sky130_fd_sc_hd__decap_3 PHY_1457 ();
 sky130_fd_sc_hd__decap_3 PHY_1458 ();
 sky130_fd_sc_hd__decap_3 PHY_1459 ();
 sky130_fd_sc_hd__decap_3 PHY_1460 ();
 sky130_fd_sc_hd__decap_3 PHY_1461 ();
 sky130_fd_sc_hd__decap_3 PHY_1462 ();
 sky130_fd_sc_hd__decap_3 PHY_1463 ();
 sky130_fd_sc_hd__decap_3 PHY_1464 ();
 sky130_fd_sc_hd__decap_3 PHY_1465 ();
 sky130_fd_sc_hd__decap_3 PHY_1466 ();
 sky130_fd_sc_hd__decap_3 PHY_1467 ();
 sky130_fd_sc_hd__decap_3 PHY_1468 ();
 sky130_fd_sc_hd__decap_3 PHY_1469 ();
 sky130_fd_sc_hd__decap_3 PHY_1470 ();
 sky130_fd_sc_hd__decap_3 PHY_1471 ();
 sky130_fd_sc_hd__decap_3 PHY_1472 ();
 sky130_fd_sc_hd__decap_3 PHY_1473 ();
 sky130_fd_sc_hd__decap_3 PHY_1474 ();
 sky130_fd_sc_hd__decap_3 PHY_1475 ();
 sky130_fd_sc_hd__decap_3 PHY_1476 ();
 sky130_fd_sc_hd__decap_3 PHY_1477 ();
 sky130_fd_sc_hd__decap_3 PHY_1478 ();
 sky130_fd_sc_hd__decap_3 PHY_1479 ();
 sky130_fd_sc_hd__decap_3 PHY_1480 ();
 sky130_fd_sc_hd__decap_3 PHY_1481 ();
 sky130_fd_sc_hd__decap_3 PHY_1482 ();
 sky130_fd_sc_hd__decap_3 PHY_1483 ();
 sky130_fd_sc_hd__decap_3 PHY_1484 ();
 sky130_fd_sc_hd__decap_3 PHY_1485 ();
 sky130_fd_sc_hd__decap_3 PHY_1486 ();
 sky130_fd_sc_hd__decap_3 PHY_1487 ();
 sky130_fd_sc_hd__decap_3 PHY_1488 ();
 sky130_fd_sc_hd__decap_3 PHY_1489 ();
 sky130_fd_sc_hd__decap_3 PHY_1490 ();
 sky130_fd_sc_hd__decap_3 PHY_1491 ();
 sky130_fd_sc_hd__decap_3 PHY_1492 ();
 sky130_fd_sc_hd__decap_3 PHY_1493 ();
 sky130_fd_sc_hd__decap_3 PHY_1494 ();
 sky130_fd_sc_hd__decap_3 PHY_1495 ();
 sky130_fd_sc_hd__decap_3 PHY_1496 ();
 sky130_fd_sc_hd__decap_3 PHY_1497 ();
 sky130_fd_sc_hd__decap_3 PHY_1498 ();
 sky130_fd_sc_hd__decap_3 PHY_1499 ();
 sky130_fd_sc_hd__decap_3 PHY_1500 ();
 sky130_fd_sc_hd__decap_3 PHY_1501 ();
 sky130_fd_sc_hd__decap_3 PHY_1502 ();
 sky130_fd_sc_hd__decap_3 PHY_1503 ();
 sky130_fd_sc_hd__decap_3 PHY_1504 ();
 sky130_fd_sc_hd__decap_3 PHY_1505 ();
 sky130_fd_sc_hd__decap_3 PHY_1506 ();
 sky130_fd_sc_hd__decap_3 PHY_1507 ();
 sky130_fd_sc_hd__decap_3 PHY_1508 ();
 sky130_fd_sc_hd__decap_3 PHY_1509 ();
 sky130_fd_sc_hd__decap_3 PHY_1510 ();
 sky130_fd_sc_hd__decap_3 PHY_1511 ();
 sky130_fd_sc_hd__decap_3 PHY_1512 ();
 sky130_fd_sc_hd__decap_3 PHY_1513 ();
 sky130_fd_sc_hd__decap_3 PHY_1514 ();
 sky130_fd_sc_hd__decap_3 PHY_1515 ();
 sky130_fd_sc_hd__decap_3 PHY_1516 ();
 sky130_fd_sc_hd__decap_3 PHY_1517 ();
 sky130_fd_sc_hd__decap_3 PHY_1518 ();
 sky130_fd_sc_hd__decap_3 PHY_1519 ();
 sky130_fd_sc_hd__decap_3 PHY_1520 ();
 sky130_fd_sc_hd__decap_3 PHY_1521 ();
 sky130_fd_sc_hd__decap_3 PHY_1522 ();
 sky130_fd_sc_hd__decap_3 PHY_1523 ();
 sky130_fd_sc_hd__decap_3 PHY_1524 ();
 sky130_fd_sc_hd__decap_3 PHY_1525 ();
 sky130_fd_sc_hd__decap_3 PHY_1526 ();
 sky130_fd_sc_hd__decap_3 PHY_1527 ();
 sky130_fd_sc_hd__decap_3 PHY_1528 ();
 sky130_fd_sc_hd__decap_3 PHY_1529 ();
 sky130_fd_sc_hd__decap_3 PHY_1530 ();
 sky130_fd_sc_hd__decap_3 PHY_1531 ();
 sky130_fd_sc_hd__decap_3 PHY_1532 ();
 sky130_fd_sc_hd__decap_3 PHY_1533 ();
 sky130_fd_sc_hd__decap_3 PHY_1534 ();
 sky130_fd_sc_hd__decap_3 PHY_1535 ();
 sky130_fd_sc_hd__decap_3 PHY_1536 ();
 sky130_fd_sc_hd__decap_3 PHY_1537 ();
 sky130_fd_sc_hd__decap_3 PHY_1538 ();
 sky130_fd_sc_hd__decap_3 PHY_1539 ();
 sky130_fd_sc_hd__decap_3 PHY_1540 ();
 sky130_fd_sc_hd__decap_3 PHY_1541 ();
 sky130_fd_sc_hd__decap_3 PHY_1542 ();
 sky130_fd_sc_hd__decap_3 PHY_1543 ();
 sky130_fd_sc_hd__decap_3 PHY_1544 ();
 sky130_fd_sc_hd__decap_3 PHY_1545 ();
 sky130_fd_sc_hd__decap_3 PHY_1546 ();
 sky130_fd_sc_hd__decap_3 PHY_1547 ();
 sky130_fd_sc_hd__decap_3 PHY_1548 ();
 sky130_fd_sc_hd__decap_3 PHY_1549 ();
 sky130_fd_sc_hd__decap_3 PHY_1550 ();
 sky130_fd_sc_hd__decap_3 PHY_1551 ();
 sky130_fd_sc_hd__decap_3 PHY_1552 ();
 sky130_fd_sc_hd__decap_3 PHY_1553 ();
 sky130_fd_sc_hd__decap_3 PHY_1554 ();
 sky130_fd_sc_hd__decap_3 PHY_1555 ();
 sky130_fd_sc_hd__decap_3 PHY_1556 ();
 sky130_fd_sc_hd__decap_3 PHY_1557 ();
 sky130_fd_sc_hd__decap_3 PHY_1558 ();
 sky130_fd_sc_hd__decap_3 PHY_1559 ();
 sky130_fd_sc_hd__decap_3 PHY_1560 ();
 sky130_fd_sc_hd__decap_3 PHY_1561 ();
 sky130_fd_sc_hd__decap_3 PHY_1562 ();
 sky130_fd_sc_hd__decap_3 PHY_1563 ();
 sky130_fd_sc_hd__decap_3 PHY_1564 ();
 sky130_fd_sc_hd__decap_3 PHY_1565 ();
 sky130_fd_sc_hd__decap_3 PHY_1566 ();
 sky130_fd_sc_hd__decap_3 PHY_1567 ();
 sky130_fd_sc_hd__decap_3 PHY_1568 ();
 sky130_fd_sc_hd__decap_3 PHY_1569 ();
 sky130_fd_sc_hd__decap_3 PHY_1570 ();
 sky130_fd_sc_hd__decap_3 PHY_1571 ();
 sky130_fd_sc_hd__decap_3 PHY_1572 ();
 sky130_fd_sc_hd__decap_3 PHY_1573 ();
 sky130_fd_sc_hd__decap_3 PHY_1574 ();
 sky130_fd_sc_hd__decap_3 PHY_1575 ();
 sky130_fd_sc_hd__decap_3 PHY_1576 ();
 sky130_fd_sc_hd__decap_3 PHY_1577 ();
 sky130_fd_sc_hd__decap_3 PHY_1578 ();
 sky130_fd_sc_hd__decap_3 PHY_1579 ();
 sky130_fd_sc_hd__decap_3 PHY_1580 ();
 sky130_fd_sc_hd__decap_3 PHY_1581 ();
 sky130_fd_sc_hd__decap_3 PHY_1582 ();
 sky130_fd_sc_hd__decap_3 PHY_1583 ();
 sky130_fd_sc_hd__decap_3 PHY_1584 ();
 sky130_fd_sc_hd__decap_3 PHY_1585 ();
 sky130_fd_sc_hd__decap_3 PHY_1586 ();
 sky130_fd_sc_hd__decap_3 PHY_1587 ();
 sky130_fd_sc_hd__decap_3 PHY_1588 ();
 sky130_fd_sc_hd__decap_3 PHY_1589 ();
 sky130_fd_sc_hd__decap_3 PHY_1590 ();
 sky130_fd_sc_hd__decap_3 PHY_1591 ();
 sky130_fd_sc_hd__decap_3 PHY_1592 ();
 sky130_fd_sc_hd__decap_3 PHY_1593 ();
 sky130_fd_sc_hd__decap_3 PHY_1594 ();
 sky130_fd_sc_hd__decap_3 PHY_1595 ();
 sky130_fd_sc_hd__decap_3 PHY_1596 ();
 sky130_fd_sc_hd__decap_3 PHY_1597 ();
 sky130_fd_sc_hd__decap_3 PHY_1598 ();
 sky130_fd_sc_hd__decap_3 PHY_1599 ();
 sky130_fd_sc_hd__decap_3 PHY_1600 ();
 sky130_fd_sc_hd__decap_3 PHY_1601 ();
 sky130_fd_sc_hd__decap_3 PHY_1602 ();
 sky130_fd_sc_hd__decap_3 PHY_1603 ();
 sky130_fd_sc_hd__decap_3 PHY_1604 ();
 sky130_fd_sc_hd__decap_3 PHY_1605 ();
 sky130_fd_sc_hd__decap_3 PHY_1606 ();
 sky130_fd_sc_hd__decap_3 PHY_1607 ();
 sky130_fd_sc_hd__decap_3 PHY_1608 ();
 sky130_fd_sc_hd__decap_3 PHY_1609 ();
 sky130_fd_sc_hd__decap_3 PHY_1610 ();
 sky130_fd_sc_hd__decap_3 PHY_1611 ();
 sky130_fd_sc_hd__decap_3 PHY_1612 ();
 sky130_fd_sc_hd__decap_3 PHY_1613 ();
 sky130_fd_sc_hd__decap_3 PHY_1614 ();
 sky130_fd_sc_hd__decap_3 PHY_1615 ();
 sky130_fd_sc_hd__decap_3 PHY_1616 ();
 sky130_fd_sc_hd__decap_3 PHY_1617 ();
 sky130_fd_sc_hd__decap_3 PHY_1618 ();
 sky130_fd_sc_hd__decap_3 PHY_1619 ();
 sky130_fd_sc_hd__decap_3 PHY_1620 ();
 sky130_fd_sc_hd__decap_3 PHY_1621 ();
 sky130_fd_sc_hd__decap_3 PHY_1622 ();
 sky130_fd_sc_hd__decap_3 PHY_1623 ();
 sky130_fd_sc_hd__decap_3 PHY_1624 ();
 sky130_fd_sc_hd__decap_3 PHY_1625 ();
 sky130_fd_sc_hd__decap_3 PHY_1626 ();
 sky130_fd_sc_hd__decap_3 PHY_1627 ();
 sky130_fd_sc_hd__decap_3 PHY_1628 ();
 sky130_fd_sc_hd__decap_3 PHY_1629 ();
 sky130_fd_sc_hd__decap_3 PHY_1630 ();
 sky130_fd_sc_hd__decap_3 PHY_1631 ();
 sky130_fd_sc_hd__decap_3 PHY_1632 ();
 sky130_fd_sc_hd__decap_3 PHY_1633 ();
 sky130_fd_sc_hd__decap_3 PHY_1634 ();
 sky130_fd_sc_hd__decap_3 PHY_1635 ();
 sky130_fd_sc_hd__decap_3 PHY_1636 ();
 sky130_fd_sc_hd__decap_3 PHY_1637 ();
 sky130_fd_sc_hd__decap_3 PHY_1638 ();
 sky130_fd_sc_hd__decap_3 PHY_1639 ();
 sky130_fd_sc_hd__decap_3 PHY_1640 ();
 sky130_fd_sc_hd__decap_3 PHY_1641 ();
 sky130_fd_sc_hd__decap_3 PHY_1642 ();
 sky130_fd_sc_hd__decap_3 PHY_1643 ();
 sky130_fd_sc_hd__decap_3 PHY_1644 ();
 sky130_fd_sc_hd__decap_3 PHY_1645 ();
 sky130_fd_sc_hd__decap_3 PHY_1646 ();
 sky130_fd_sc_hd__decap_3 PHY_1647 ();
 sky130_fd_sc_hd__decap_3 PHY_1648 ();
 sky130_fd_sc_hd__decap_3 PHY_1649 ();
 sky130_fd_sc_hd__decap_3 PHY_1650 ();
 sky130_fd_sc_hd__decap_3 PHY_1651 ();
 sky130_fd_sc_hd__decap_3 PHY_1652 ();
 sky130_fd_sc_hd__decap_3 PHY_1653 ();
 sky130_fd_sc_hd__decap_3 PHY_1654 ();
 sky130_fd_sc_hd__decap_3 PHY_1655 ();
 sky130_fd_sc_hd__decap_3 PHY_1656 ();
 sky130_fd_sc_hd__decap_3 PHY_1657 ();
 sky130_fd_sc_hd__decap_3 PHY_1658 ();
 sky130_fd_sc_hd__decap_3 PHY_1659 ();
 sky130_fd_sc_hd__decap_3 PHY_1660 ();
 sky130_fd_sc_hd__decap_3 PHY_1661 ();
 sky130_fd_sc_hd__decap_3 PHY_1662 ();
 sky130_fd_sc_hd__decap_3 PHY_1663 ();
 sky130_fd_sc_hd__decap_3 PHY_1664 ();
 sky130_fd_sc_hd__decap_3 PHY_1665 ();
 sky130_fd_sc_hd__decap_3 PHY_1666 ();
 sky130_fd_sc_hd__decap_3 PHY_1667 ();
 sky130_fd_sc_hd__decap_3 PHY_1668 ();
 sky130_fd_sc_hd__decap_3 PHY_1669 ();
 sky130_fd_sc_hd__decap_3 PHY_1670 ();
 sky130_fd_sc_hd__decap_3 PHY_1671 ();
 sky130_fd_sc_hd__decap_3 PHY_1672 ();
 sky130_fd_sc_hd__decap_3 PHY_1673 ();
 sky130_fd_sc_hd__decap_3 PHY_1674 ();
 sky130_fd_sc_hd__decap_3 PHY_1675 ();
 sky130_fd_sc_hd__decap_3 PHY_1676 ();
 sky130_fd_sc_hd__decap_3 PHY_1677 ();
 sky130_fd_sc_hd__decap_3 PHY_1678 ();
 sky130_fd_sc_hd__decap_3 PHY_1679 ();
 sky130_fd_sc_hd__decap_3 PHY_1680 ();
 sky130_fd_sc_hd__decap_3 PHY_1681 ();
 sky130_fd_sc_hd__decap_3 PHY_1682 ();
 sky130_fd_sc_hd__decap_3 PHY_1683 ();
 sky130_fd_sc_hd__decap_3 PHY_1684 ();
 sky130_fd_sc_hd__decap_3 PHY_1685 ();
 sky130_fd_sc_hd__decap_3 PHY_1686 ();
 sky130_fd_sc_hd__decap_3 PHY_1687 ();
 sky130_fd_sc_hd__decap_3 PHY_1688 ();
 sky130_fd_sc_hd__decap_3 PHY_1689 ();
 sky130_fd_sc_hd__decap_3 PHY_1690 ();
 sky130_fd_sc_hd__decap_3 PHY_1691 ();
 sky130_fd_sc_hd__decap_3 PHY_1692 ();
 sky130_fd_sc_hd__decap_3 PHY_1693 ();
 sky130_fd_sc_hd__decap_3 PHY_1694 ();
 sky130_fd_sc_hd__decap_3 PHY_1695 ();
 sky130_fd_sc_hd__decap_3 PHY_1696 ();
 sky130_fd_sc_hd__decap_3 PHY_1697 ();
 sky130_fd_sc_hd__decap_3 PHY_1698 ();
 sky130_fd_sc_hd__decap_3 PHY_1699 ();
 sky130_fd_sc_hd__decap_3 PHY_1700 ();
 sky130_fd_sc_hd__decap_3 PHY_1701 ();
 sky130_fd_sc_hd__decap_3 PHY_1702 ();
 sky130_fd_sc_hd__decap_3 PHY_1703 ();
 sky130_fd_sc_hd__decap_3 PHY_1704 ();
 sky130_fd_sc_hd__decap_3 PHY_1705 ();
 sky130_fd_sc_hd__decap_3 PHY_1706 ();
 sky130_fd_sc_hd__decap_3 PHY_1707 ();
 sky130_fd_sc_hd__decap_3 PHY_1708 ();
 sky130_fd_sc_hd__decap_3 PHY_1709 ();
 sky130_fd_sc_hd__decap_3 PHY_1710 ();
 sky130_fd_sc_hd__decap_3 PHY_1711 ();
 sky130_fd_sc_hd__decap_3 PHY_1712 ();
 sky130_fd_sc_hd__decap_3 PHY_1713 ();
 sky130_fd_sc_hd__decap_3 PHY_1714 ();
 sky130_fd_sc_hd__decap_3 PHY_1715 ();
 sky130_fd_sc_hd__decap_3 PHY_1716 ();
 sky130_fd_sc_hd__decap_3 PHY_1717 ();
 sky130_fd_sc_hd__decap_3 PHY_1718 ();
 sky130_fd_sc_hd__decap_3 PHY_1719 ();
 sky130_fd_sc_hd__decap_3 PHY_1720 ();
 sky130_fd_sc_hd__decap_3 PHY_1721 ();
 sky130_fd_sc_hd__decap_3 PHY_1722 ();
 sky130_fd_sc_hd__decap_3 PHY_1723 ();
 sky130_fd_sc_hd__decap_3 PHY_1724 ();
 sky130_fd_sc_hd__decap_3 PHY_1725 ();
 sky130_fd_sc_hd__decap_3 PHY_1726 ();
 sky130_fd_sc_hd__decap_3 PHY_1727 ();
 sky130_fd_sc_hd__decap_3 PHY_1728 ();
 sky130_fd_sc_hd__decap_3 PHY_1729 ();
 sky130_fd_sc_hd__decap_3 PHY_1730 ();
 sky130_fd_sc_hd__decap_3 PHY_1731 ();
 sky130_fd_sc_hd__decap_3 PHY_1732 ();
 sky130_fd_sc_hd__decap_3 PHY_1733 ();
 sky130_fd_sc_hd__decap_3 PHY_1734 ();
 sky130_fd_sc_hd__decap_3 PHY_1735 ();
 sky130_fd_sc_hd__decap_3 PHY_1736 ();
 sky130_fd_sc_hd__decap_3 PHY_1737 ();
 sky130_fd_sc_hd__decap_3 PHY_1738 ();
 sky130_fd_sc_hd__decap_3 PHY_1739 ();
 sky130_fd_sc_hd__decap_3 PHY_1740 ();
 sky130_fd_sc_hd__decap_3 PHY_1741 ();
 sky130_fd_sc_hd__decap_3 PHY_1742 ();
 sky130_fd_sc_hd__decap_3 PHY_1743 ();
 sky130_fd_sc_hd__decap_3 PHY_1744 ();
 sky130_fd_sc_hd__decap_3 PHY_1745 ();
 sky130_fd_sc_hd__decap_3 PHY_1746 ();
 sky130_fd_sc_hd__decap_3 PHY_1747 ();
 sky130_fd_sc_hd__decap_3 PHY_1748 ();
 sky130_fd_sc_hd__decap_3 PHY_1749 ();
 sky130_fd_sc_hd__decap_3 PHY_1750 ();
 sky130_fd_sc_hd__decap_3 PHY_1751 ();
 sky130_fd_sc_hd__decap_3 PHY_1752 ();
 sky130_fd_sc_hd__decap_3 PHY_1753 ();
 sky130_fd_sc_hd__decap_3 PHY_1754 ();
 sky130_fd_sc_hd__decap_3 PHY_1755 ();
 sky130_fd_sc_hd__decap_3 PHY_1756 ();
 sky130_fd_sc_hd__decap_3 PHY_1757 ();
 sky130_fd_sc_hd__decap_3 PHY_1758 ();
 sky130_fd_sc_hd__decap_3 PHY_1759 ();
 sky130_fd_sc_hd__decap_3 PHY_1760 ();
 sky130_fd_sc_hd__decap_3 PHY_1761 ();
 sky130_fd_sc_hd__decap_3 PHY_1762 ();
 sky130_fd_sc_hd__decap_3 PHY_1763 ();
 sky130_fd_sc_hd__decap_3 PHY_1764 ();
 sky130_fd_sc_hd__decap_3 PHY_1765 ();
 sky130_fd_sc_hd__decap_3 PHY_1766 ();
 sky130_fd_sc_hd__decap_3 PHY_1767 ();
 sky130_fd_sc_hd__decap_3 PHY_1768 ();
 sky130_fd_sc_hd__decap_3 PHY_1769 ();
 sky130_fd_sc_hd__decap_3 PHY_1770 ();
 sky130_fd_sc_hd__decap_3 PHY_1771 ();
 sky130_fd_sc_hd__decap_3 PHY_1772 ();
 sky130_fd_sc_hd__decap_3 PHY_1773 ();
 sky130_fd_sc_hd__decap_3 PHY_1774 ();
 sky130_fd_sc_hd__decap_3 PHY_1775 ();
 sky130_fd_sc_hd__decap_3 PHY_1776 ();
 sky130_fd_sc_hd__decap_3 PHY_1777 ();
 sky130_fd_sc_hd__decap_3 PHY_1778 ();
 sky130_fd_sc_hd__decap_3 PHY_1779 ();
 sky130_fd_sc_hd__decap_3 PHY_1780 ();
 sky130_fd_sc_hd__decap_3 PHY_1781 ();
 sky130_fd_sc_hd__decap_3 PHY_1782 ();
 sky130_fd_sc_hd__decap_3 PHY_1783 ();
 sky130_fd_sc_hd__decap_3 PHY_1784 ();
 sky130_fd_sc_hd__decap_3 PHY_1785 ();
 sky130_fd_sc_hd__decap_3 PHY_1786 ();
 sky130_fd_sc_hd__decap_3 PHY_1787 ();
 sky130_fd_sc_hd__decap_3 PHY_1788 ();
 sky130_fd_sc_hd__decap_3 PHY_1789 ();
 sky130_fd_sc_hd__decap_3 PHY_1790 ();
 sky130_fd_sc_hd__decap_3 PHY_1791 ();
 sky130_fd_sc_hd__decap_3 PHY_1792 ();
 sky130_fd_sc_hd__decap_3 PHY_1793 ();
 sky130_fd_sc_hd__decap_3 PHY_1794 ();
 sky130_fd_sc_hd__decap_3 PHY_1795 ();
 sky130_fd_sc_hd__decap_3 PHY_1796 ();
 sky130_fd_sc_hd__decap_3 PHY_1797 ();
 sky130_fd_sc_hd__decap_3 PHY_1798 ();
 sky130_fd_sc_hd__decap_3 PHY_1799 ();
 sky130_fd_sc_hd__decap_3 PHY_1800 ();
 sky130_fd_sc_hd__decap_3 PHY_1801 ();
 sky130_fd_sc_hd__decap_3 PHY_1802 ();
 sky130_fd_sc_hd__decap_3 PHY_1803 ();
 sky130_fd_sc_hd__decap_3 PHY_1804 ();
 sky130_fd_sc_hd__decap_3 PHY_1805 ();
 sky130_fd_sc_hd__decap_3 PHY_1806 ();
 sky130_fd_sc_hd__decap_3 PHY_1807 ();
 sky130_fd_sc_hd__decap_3 PHY_1808 ();
 sky130_fd_sc_hd__decap_3 PHY_1809 ();
 sky130_fd_sc_hd__decap_3 PHY_1810 ();
 sky130_fd_sc_hd__decap_3 PHY_1811 ();
 sky130_fd_sc_hd__decap_3 PHY_1812 ();
 sky130_fd_sc_hd__decap_3 PHY_1813 ();
 sky130_fd_sc_hd__decap_3 PHY_1814 ();
 sky130_fd_sc_hd__decap_3 PHY_1815 ();
 sky130_fd_sc_hd__decap_3 PHY_1816 ();
 sky130_fd_sc_hd__decap_3 PHY_1817 ();
 sky130_fd_sc_hd__decap_3 PHY_1818 ();
 sky130_fd_sc_hd__decap_3 PHY_1819 ();
 sky130_fd_sc_hd__decap_3 PHY_1820 ();
 sky130_fd_sc_hd__decap_3 PHY_1821 ();
 sky130_fd_sc_hd__decap_3 PHY_1822 ();
 sky130_fd_sc_hd__decap_3 PHY_1823 ();
 sky130_fd_sc_hd__decap_3 PHY_1824 ();
 sky130_fd_sc_hd__decap_3 PHY_1825 ();
 sky130_fd_sc_hd__decap_3 PHY_1826 ();
 sky130_fd_sc_hd__decap_3 PHY_1827 ();
 sky130_fd_sc_hd__decap_3 PHY_1828 ();
 sky130_fd_sc_hd__decap_3 PHY_1829 ();
 sky130_fd_sc_hd__decap_3 PHY_1830 ();
 sky130_fd_sc_hd__decap_3 PHY_1831 ();
 sky130_fd_sc_hd__decap_3 PHY_1832 ();
 sky130_fd_sc_hd__decap_3 PHY_1833 ();
 sky130_fd_sc_hd__decap_3 PHY_1834 ();
 sky130_fd_sc_hd__decap_3 PHY_1835 ();
 sky130_fd_sc_hd__decap_3 PHY_1836 ();
 sky130_fd_sc_hd__decap_3 PHY_1837 ();
 sky130_fd_sc_hd__decap_3 PHY_1838 ();
 sky130_fd_sc_hd__decap_3 PHY_1839 ();
 sky130_fd_sc_hd__decap_3 PHY_1840 ();
 sky130_fd_sc_hd__decap_3 PHY_1841 ();
 sky130_fd_sc_hd__decap_3 PHY_1842 ();
 sky130_fd_sc_hd__decap_3 PHY_1843 ();
 sky130_fd_sc_hd__decap_3 PHY_1844 ();
 sky130_fd_sc_hd__decap_3 PHY_1845 ();
 sky130_fd_sc_hd__decap_3 PHY_1846 ();
 sky130_fd_sc_hd__decap_3 PHY_1847 ();
 sky130_fd_sc_hd__decap_3 PHY_1848 ();
 sky130_fd_sc_hd__decap_3 PHY_1849 ();
 sky130_fd_sc_hd__decap_3 PHY_1850 ();
 sky130_fd_sc_hd__decap_3 PHY_1851 ();
 sky130_fd_sc_hd__decap_3 PHY_1852 ();
 sky130_fd_sc_hd__decap_3 PHY_1853 ();
 sky130_fd_sc_hd__decap_3 PHY_1854 ();
 sky130_fd_sc_hd__decap_3 PHY_1855 ();
 sky130_fd_sc_hd__decap_3 PHY_1856 ();
 sky130_fd_sc_hd__decap_3 PHY_1857 ();
 sky130_fd_sc_hd__decap_3 PHY_1858 ();
 sky130_fd_sc_hd__decap_3 PHY_1859 ();
 sky130_fd_sc_hd__decap_3 PHY_1860 ();
 sky130_fd_sc_hd__decap_3 PHY_1861 ();
 sky130_fd_sc_hd__decap_3 PHY_1862 ();
 sky130_fd_sc_hd__decap_3 PHY_1863 ();
 sky130_fd_sc_hd__decap_3 PHY_1864 ();
 sky130_fd_sc_hd__decap_3 PHY_1865 ();
 sky130_fd_sc_hd__decap_3 PHY_1866 ();
 sky130_fd_sc_hd__decap_3 PHY_1867 ();
 sky130_fd_sc_hd__decap_3 PHY_1868 ();
 sky130_fd_sc_hd__decap_3 PHY_1869 ();
 sky130_fd_sc_hd__decap_3 PHY_1870 ();
 sky130_fd_sc_hd__decap_3 PHY_1871 ();
 sky130_fd_sc_hd__decap_3 PHY_1872 ();
 sky130_fd_sc_hd__decap_3 PHY_1873 ();
 sky130_fd_sc_hd__decap_3 PHY_1874 ();
 sky130_fd_sc_hd__decap_3 PHY_1875 ();
 sky130_fd_sc_hd__decap_3 PHY_1876 ();
 sky130_fd_sc_hd__decap_3 PHY_1877 ();
 sky130_fd_sc_hd__decap_3 PHY_1878 ();
 sky130_fd_sc_hd__decap_3 PHY_1879 ();
 sky130_fd_sc_hd__decap_3 PHY_1880 ();
 sky130_fd_sc_hd__decap_3 PHY_1881 ();
 sky130_fd_sc_hd__decap_3 PHY_1882 ();
 sky130_fd_sc_hd__decap_3 PHY_1883 ();
 sky130_fd_sc_hd__decap_3 PHY_1884 ();
 sky130_fd_sc_hd__decap_3 PHY_1885 ();
 sky130_fd_sc_hd__decap_3 PHY_1886 ();
 sky130_fd_sc_hd__decap_3 PHY_1887 ();
 sky130_fd_sc_hd__decap_3 PHY_1888 ();
 sky130_fd_sc_hd__decap_3 PHY_1889 ();
 sky130_fd_sc_hd__decap_3 PHY_1890 ();
 sky130_fd_sc_hd__decap_3 PHY_1891 ();
 sky130_fd_sc_hd__decap_3 PHY_1892 ();
 sky130_fd_sc_hd__decap_3 PHY_1893 ();
 sky130_fd_sc_hd__decap_3 PHY_1894 ();
 sky130_fd_sc_hd__decap_3 PHY_1895 ();
 sky130_fd_sc_hd__decap_3 PHY_1896 ();
 sky130_fd_sc_hd__decap_3 PHY_1897 ();
 sky130_fd_sc_hd__decap_3 PHY_1898 ();
 sky130_fd_sc_hd__decap_3 PHY_1899 ();
 sky130_fd_sc_hd__decap_3 PHY_1900 ();
 sky130_fd_sc_hd__decap_3 PHY_1901 ();
 sky130_fd_sc_hd__decap_3 PHY_1902 ();
 sky130_fd_sc_hd__decap_3 PHY_1903 ();
 sky130_fd_sc_hd__decap_3 PHY_1904 ();
 sky130_fd_sc_hd__decap_3 PHY_1905 ();
 sky130_fd_sc_hd__decap_3 PHY_1906 ();
 sky130_fd_sc_hd__decap_3 PHY_1907 ();
 sky130_fd_sc_hd__decap_3 PHY_1908 ();
 sky130_fd_sc_hd__decap_3 PHY_1909 ();
 sky130_fd_sc_hd__decap_3 PHY_1910 ();
 sky130_fd_sc_hd__decap_3 PHY_1911 ();
 sky130_fd_sc_hd__decap_3 PHY_1912 ();
 sky130_fd_sc_hd__decap_3 PHY_1913 ();
 sky130_fd_sc_hd__decap_3 PHY_1914 ();
 sky130_fd_sc_hd__decap_3 PHY_1915 ();
 sky130_fd_sc_hd__decap_3 PHY_1916 ();
 sky130_fd_sc_hd__decap_3 PHY_1917 ();
 sky130_fd_sc_hd__decap_3 PHY_1918 ();
 sky130_fd_sc_hd__decap_3 PHY_1919 ();
 sky130_fd_sc_hd__decap_3 PHY_1920 ();
 sky130_fd_sc_hd__decap_3 PHY_1921 ();
 sky130_fd_sc_hd__decap_3 PHY_1922 ();
 sky130_fd_sc_hd__decap_3 PHY_1923 ();
 sky130_fd_sc_hd__decap_3 PHY_1924 ();
 sky130_fd_sc_hd__decap_3 PHY_1925 ();
 sky130_fd_sc_hd__decap_3 PHY_1926 ();
 sky130_fd_sc_hd__decap_3 PHY_1927 ();
 sky130_fd_sc_hd__decap_3 PHY_1928 ();
 sky130_fd_sc_hd__decap_3 PHY_1929 ();
 sky130_fd_sc_hd__decap_3 PHY_1930 ();
 sky130_fd_sc_hd__decap_3 PHY_1931 ();
 sky130_fd_sc_hd__decap_3 PHY_1932 ();
 sky130_fd_sc_hd__decap_3 PHY_1933 ();
 sky130_fd_sc_hd__decap_3 PHY_1934 ();
 sky130_fd_sc_hd__decap_3 PHY_1935 ();
 sky130_fd_sc_hd__decap_3 PHY_1936 ();
 sky130_fd_sc_hd__decap_3 PHY_1937 ();
 sky130_fd_sc_hd__decap_3 PHY_1938 ();
 sky130_fd_sc_hd__decap_3 PHY_1939 ();
 sky130_fd_sc_hd__decap_3 PHY_1940 ();
 sky130_fd_sc_hd__decap_3 PHY_1941 ();
 sky130_fd_sc_hd__decap_3 PHY_1942 ();
 sky130_fd_sc_hd__decap_3 PHY_1943 ();
 sky130_fd_sc_hd__decap_3 PHY_1944 ();
 sky130_fd_sc_hd__decap_3 PHY_1945 ();
 sky130_fd_sc_hd__decap_3 PHY_1946 ();
 sky130_fd_sc_hd__decap_3 PHY_1947 ();
 sky130_fd_sc_hd__decap_3 PHY_1948 ();
 sky130_fd_sc_hd__decap_3 PHY_1949 ();
 sky130_fd_sc_hd__decap_3 PHY_1950 ();
 sky130_fd_sc_hd__decap_3 PHY_1951 ();
 sky130_fd_sc_hd__decap_3 PHY_1952 ();
 sky130_fd_sc_hd__decap_3 PHY_1953 ();
 sky130_fd_sc_hd__decap_3 PHY_1954 ();
 sky130_fd_sc_hd__decap_3 PHY_1955 ();
 sky130_fd_sc_hd__decap_3 PHY_1956 ();
 sky130_fd_sc_hd__decap_3 PHY_1957 ();
 sky130_fd_sc_hd__decap_3 PHY_1958 ();
 sky130_fd_sc_hd__decap_3 PHY_1959 ();
 sky130_fd_sc_hd__decap_3 PHY_1960 ();
 sky130_fd_sc_hd__decap_3 PHY_1961 ();
 sky130_fd_sc_hd__decap_3 PHY_1962 ();
 sky130_fd_sc_hd__decap_3 PHY_1963 ();
 sky130_fd_sc_hd__decap_3 PHY_1964 ();
 sky130_fd_sc_hd__decap_3 PHY_1965 ();
 sky130_fd_sc_hd__decap_3 PHY_1966 ();
 sky130_fd_sc_hd__decap_3 PHY_1967 ();
 sky130_fd_sc_hd__decap_3 PHY_1968 ();
 sky130_fd_sc_hd__decap_3 PHY_1969 ();
 sky130_fd_sc_hd__decap_3 PHY_1970 ();
 sky130_fd_sc_hd__decap_3 PHY_1971 ();
 sky130_fd_sc_hd__decap_3 PHY_1972 ();
 sky130_fd_sc_hd__decap_3 PHY_1973 ();
 sky130_fd_sc_hd__decap_3 PHY_1974 ();
 sky130_fd_sc_hd__decap_3 PHY_1975 ();
 sky130_fd_sc_hd__decap_3 PHY_1976 ();
 sky130_fd_sc_hd__decap_3 PHY_1977 ();
 sky130_fd_sc_hd__decap_3 PHY_1978 ();
 sky130_fd_sc_hd__decap_3 PHY_1979 ();
 sky130_fd_sc_hd__decap_3 PHY_1980 ();
 sky130_fd_sc_hd__decap_3 PHY_1981 ();
 sky130_fd_sc_hd__decap_3 PHY_1982 ();
 sky130_fd_sc_hd__decap_3 PHY_1983 ();
 sky130_fd_sc_hd__decap_3 PHY_1984 ();
 sky130_fd_sc_hd__decap_3 PHY_1985 ();
 sky130_fd_sc_hd__decap_3 PHY_1986 ();
 sky130_fd_sc_hd__decap_3 PHY_1987 ();
 sky130_fd_sc_hd__decap_3 PHY_1988 ();
 sky130_fd_sc_hd__decap_3 PHY_1989 ();
 sky130_fd_sc_hd__decap_3 PHY_1990 ();
 sky130_fd_sc_hd__decap_3 PHY_1991 ();
 sky130_fd_sc_hd__decap_3 PHY_1992 ();
 sky130_fd_sc_hd__decap_3 PHY_1993 ();
 sky130_fd_sc_hd__decap_3 PHY_1994 ();
 sky130_fd_sc_hd__decap_3 PHY_1995 ();
 sky130_fd_sc_hd__decap_3 PHY_1996 ();
 sky130_fd_sc_hd__decap_3 PHY_1997 ();
 sky130_fd_sc_hd__decap_3 PHY_1998 ();
 sky130_fd_sc_hd__decap_3 PHY_1999 ();
 sky130_fd_sc_hd__decap_3 PHY_2000 ();
 sky130_fd_sc_hd__decap_3 PHY_2001 ();
 sky130_fd_sc_hd__decap_3 PHY_2002 ();
 sky130_fd_sc_hd__decap_3 PHY_2003 ();
 sky130_fd_sc_hd__decap_3 PHY_2004 ();
 sky130_fd_sc_hd__decap_3 PHY_2005 ();
 sky130_fd_sc_hd__decap_3 PHY_2006 ();
 sky130_fd_sc_hd__decap_3 PHY_2007 ();
 sky130_fd_sc_hd__decap_3 PHY_2008 ();
 sky130_fd_sc_hd__decap_3 PHY_2009 ();
 sky130_fd_sc_hd__decap_3 PHY_2010 ();
 sky130_fd_sc_hd__decap_3 PHY_2011 ();
 sky130_fd_sc_hd__decap_3 PHY_2012 ();
 sky130_fd_sc_hd__decap_3 PHY_2013 ();
 sky130_fd_sc_hd__decap_3 PHY_2014 ();
 sky130_fd_sc_hd__decap_3 PHY_2015 ();
 sky130_fd_sc_hd__decap_3 PHY_2016 ();
 sky130_fd_sc_hd__decap_3 PHY_2017 ();
 sky130_fd_sc_hd__decap_3 PHY_2018 ();
 sky130_fd_sc_hd__decap_3 PHY_2019 ();
 sky130_fd_sc_hd__decap_3 PHY_2020 ();
 sky130_fd_sc_hd__decap_3 PHY_2021 ();
 sky130_fd_sc_hd__decap_3 PHY_2022 ();
 sky130_fd_sc_hd__decap_3 PHY_2023 ();
 sky130_fd_sc_hd__decap_3 PHY_2024 ();
 sky130_fd_sc_hd__decap_3 PHY_2025 ();
 sky130_fd_sc_hd__decap_3 PHY_2026 ();
 sky130_fd_sc_hd__decap_3 PHY_2027 ();
 sky130_fd_sc_hd__decap_3 PHY_2028 ();
 sky130_fd_sc_hd__decap_3 PHY_2029 ();
 sky130_fd_sc_hd__decap_3 PHY_2030 ();
 sky130_fd_sc_hd__decap_3 PHY_2031 ();
 sky130_fd_sc_hd__decap_3 PHY_2032 ();
 sky130_fd_sc_hd__decap_3 PHY_2033 ();
 sky130_fd_sc_hd__decap_3 PHY_2034 ();
 sky130_fd_sc_hd__decap_3 PHY_2035 ();
 sky130_fd_sc_hd__decap_3 PHY_2036 ();
 sky130_fd_sc_hd__decap_3 PHY_2037 ();
 sky130_fd_sc_hd__decap_3 PHY_2038 ();
 sky130_fd_sc_hd__decap_3 PHY_2039 ();
 sky130_fd_sc_hd__decap_3 PHY_2040 ();
 sky130_fd_sc_hd__decap_3 PHY_2041 ();
 sky130_fd_sc_hd__decap_3 PHY_2042 ();
 sky130_fd_sc_hd__decap_3 PHY_2043 ();
 sky130_fd_sc_hd__decap_3 PHY_2044 ();
 sky130_fd_sc_hd__decap_3 PHY_2045 ();
 sky130_fd_sc_hd__decap_3 PHY_2046 ();
 sky130_fd_sc_hd__decap_3 PHY_2047 ();
 sky130_fd_sc_hd__decap_3 PHY_2048 ();
 sky130_fd_sc_hd__decap_3 PHY_2049 ();
 sky130_fd_sc_hd__decap_3 PHY_2050 ();
 sky130_fd_sc_hd__decap_3 PHY_2051 ();
 sky130_fd_sc_hd__decap_3 PHY_2052 ();
 sky130_fd_sc_hd__decap_3 PHY_2053 ();
 sky130_fd_sc_hd__decap_3 PHY_2054 ();
 sky130_fd_sc_hd__decap_3 PHY_2055 ();
 sky130_fd_sc_hd__decap_3 PHY_2056 ();
 sky130_fd_sc_hd__decap_3 PHY_2057 ();
 sky130_fd_sc_hd__decap_3 PHY_2058 ();
 sky130_fd_sc_hd__decap_3 PHY_2059 ();
 sky130_fd_sc_hd__decap_3 PHY_2060 ();
 sky130_fd_sc_hd__decap_3 PHY_2061 ();
 sky130_fd_sc_hd__decap_3 PHY_2062 ();
 sky130_fd_sc_hd__decap_3 PHY_2063 ();
 sky130_fd_sc_hd__decap_3 PHY_2064 ();
 sky130_fd_sc_hd__decap_3 PHY_2065 ();
 sky130_fd_sc_hd__decap_3 PHY_2066 ();
 sky130_fd_sc_hd__decap_3 PHY_2067 ();
 sky130_fd_sc_hd__decap_3 PHY_2068 ();
 sky130_fd_sc_hd__decap_3 PHY_2069 ();
 sky130_fd_sc_hd__decap_3 PHY_2070 ();
 sky130_fd_sc_hd__decap_3 PHY_2071 ();
 sky130_fd_sc_hd__decap_3 PHY_2072 ();
 sky130_fd_sc_hd__decap_3 PHY_2073 ();
 sky130_fd_sc_hd__decap_3 PHY_2074 ();
 sky130_fd_sc_hd__decap_3 PHY_2075 ();
 sky130_fd_sc_hd__decap_3 PHY_2076 ();
 sky130_fd_sc_hd__decap_3 PHY_2077 ();
 sky130_fd_sc_hd__decap_3 PHY_2078 ();
 sky130_fd_sc_hd__decap_3 PHY_2079 ();
 sky130_fd_sc_hd__decap_3 PHY_2080 ();
 sky130_fd_sc_hd__decap_3 PHY_2081 ();
 sky130_fd_sc_hd__decap_3 PHY_2082 ();
 sky130_fd_sc_hd__decap_3 PHY_2083 ();
 sky130_fd_sc_hd__decap_3 PHY_2084 ();
 sky130_fd_sc_hd__decap_3 PHY_2085 ();
 sky130_fd_sc_hd__decap_3 PHY_2086 ();
 sky130_fd_sc_hd__decap_3 PHY_2087 ();
 sky130_fd_sc_hd__decap_3 PHY_2088 ();
 sky130_fd_sc_hd__decap_3 PHY_2089 ();
 sky130_fd_sc_hd__decap_3 PHY_2090 ();
 sky130_fd_sc_hd__decap_3 PHY_2091 ();
 sky130_fd_sc_hd__decap_3 PHY_2092 ();
 sky130_fd_sc_hd__decap_3 PHY_2093 ();
 sky130_fd_sc_hd__decap_3 PHY_2094 ();
 sky130_fd_sc_hd__decap_3 PHY_2095 ();
 sky130_fd_sc_hd__decap_3 PHY_2096 ();
 sky130_fd_sc_hd__decap_3 PHY_2097 ();
 sky130_fd_sc_hd__decap_3 PHY_2098 ();
 sky130_fd_sc_hd__decap_3 PHY_2099 ();
 sky130_fd_sc_hd__decap_3 PHY_2100 ();
 sky130_fd_sc_hd__decap_3 PHY_2101 ();
 sky130_fd_sc_hd__decap_3 PHY_2102 ();
 sky130_fd_sc_hd__decap_3 PHY_2103 ();
 sky130_fd_sc_hd__decap_3 PHY_2104 ();
 sky130_fd_sc_hd__decap_3 PHY_2105 ();
 sky130_fd_sc_hd__decap_3 PHY_2106 ();
 sky130_fd_sc_hd__decap_3 PHY_2107 ();
 sky130_fd_sc_hd__decap_3 PHY_2108 ();
 sky130_fd_sc_hd__decap_3 PHY_2109 ();
 sky130_fd_sc_hd__decap_3 PHY_2110 ();
 sky130_fd_sc_hd__decap_3 PHY_2111 ();
 sky130_fd_sc_hd__decap_3 PHY_2112 ();
 sky130_fd_sc_hd__decap_3 PHY_2113 ();
 sky130_fd_sc_hd__decap_3 PHY_2114 ();
 sky130_fd_sc_hd__decap_3 PHY_2115 ();
 sky130_fd_sc_hd__decap_3 PHY_2116 ();
 sky130_fd_sc_hd__decap_3 PHY_2117 ();
 sky130_fd_sc_hd__decap_3 PHY_2118 ();
 sky130_fd_sc_hd__decap_3 PHY_2119 ();
 sky130_fd_sc_hd__decap_3 PHY_2120 ();
 sky130_fd_sc_hd__decap_3 PHY_2121 ();
 sky130_fd_sc_hd__decap_3 PHY_2122 ();
 sky130_fd_sc_hd__decap_3 PHY_2123 ();
 sky130_fd_sc_hd__decap_3 PHY_2124 ();
 sky130_fd_sc_hd__decap_3 PHY_2125 ();
 sky130_fd_sc_hd__decap_3 PHY_2126 ();
 sky130_fd_sc_hd__decap_3 PHY_2127 ();
 sky130_fd_sc_hd__decap_3 PHY_2128 ();
 sky130_fd_sc_hd__decap_3 PHY_2129 ();
 sky130_fd_sc_hd__decap_3 PHY_2130 ();
 sky130_fd_sc_hd__decap_3 PHY_2131 ();
 sky130_fd_sc_hd__decap_3 PHY_2132 ();
 sky130_fd_sc_hd__decap_3 PHY_2133 ();
 sky130_fd_sc_hd__decap_3 PHY_2134 ();
 sky130_fd_sc_hd__decap_3 PHY_2135 ();
 sky130_fd_sc_hd__decap_3 PHY_2136 ();
 sky130_fd_sc_hd__decap_3 PHY_2137 ();
 sky130_fd_sc_hd__decap_3 PHY_2138 ();
 sky130_fd_sc_hd__decap_3 PHY_2139 ();
 sky130_fd_sc_hd__decap_3 PHY_2140 ();
 sky130_fd_sc_hd__decap_3 PHY_2141 ();
 sky130_fd_sc_hd__decap_3 PHY_2142 ();
 sky130_fd_sc_hd__decap_3 PHY_2143 ();
 sky130_fd_sc_hd__decap_3 PHY_2144 ();
 sky130_fd_sc_hd__decap_3 PHY_2145 ();
 sky130_fd_sc_hd__decap_3 PHY_2146 ();
 sky130_fd_sc_hd__decap_3 PHY_2147 ();
 sky130_fd_sc_hd__decap_3 PHY_2148 ();
 sky130_fd_sc_hd__decap_3 PHY_2149 ();
 sky130_fd_sc_hd__decap_3 PHY_2150 ();
 sky130_fd_sc_hd__decap_3 PHY_2151 ();
 sky130_fd_sc_hd__decap_3 PHY_2152 ();
 sky130_fd_sc_hd__decap_3 PHY_2153 ();
 sky130_fd_sc_hd__decap_3 PHY_2154 ();
 sky130_fd_sc_hd__decap_3 PHY_2155 ();
 sky130_fd_sc_hd__decap_3 PHY_2156 ();
 sky130_fd_sc_hd__decap_3 PHY_2157 ();
 sky130_fd_sc_hd__decap_3 PHY_2158 ();
 sky130_fd_sc_hd__decap_3 PHY_2159 ();
 sky130_fd_sc_hd__decap_3 PHY_2160 ();
 sky130_fd_sc_hd__decap_3 PHY_2161 ();
 sky130_fd_sc_hd__decap_3 PHY_2162 ();
 sky130_fd_sc_hd__decap_3 PHY_2163 ();
 sky130_fd_sc_hd__decap_3 PHY_2164 ();
 sky130_fd_sc_hd__decap_3 PHY_2165 ();
 sky130_fd_sc_hd__decap_3 PHY_2166 ();
 sky130_fd_sc_hd__decap_3 PHY_2167 ();
 sky130_fd_sc_hd__decap_3 PHY_2168 ();
 sky130_fd_sc_hd__decap_3 PHY_2169 ();
 sky130_fd_sc_hd__decap_3 PHY_2170 ();
 sky130_fd_sc_hd__decap_3 PHY_2171 ();
 sky130_fd_sc_hd__decap_3 PHY_2172 ();
 sky130_fd_sc_hd__decap_3 PHY_2173 ();
 sky130_fd_sc_hd__decap_3 PHY_2174 ();
 sky130_fd_sc_hd__decap_3 PHY_2175 ();
 sky130_fd_sc_hd__decap_3 PHY_2176 ();
 sky130_fd_sc_hd__decap_3 PHY_2177 ();
 sky130_fd_sc_hd__decap_3 PHY_2178 ();
 sky130_fd_sc_hd__decap_3 PHY_2179 ();
 sky130_fd_sc_hd__decap_3 PHY_2180 ();
 sky130_fd_sc_hd__decap_3 PHY_2181 ();
 sky130_fd_sc_hd__decap_3 PHY_2182 ();
 sky130_fd_sc_hd__decap_3 PHY_2183 ();
 sky130_fd_sc_hd__decap_3 PHY_2184 ();
 sky130_fd_sc_hd__decap_3 PHY_2185 ();
 sky130_fd_sc_hd__decap_3 PHY_2186 ();
 sky130_fd_sc_hd__decap_3 PHY_2187 ();
 sky130_fd_sc_hd__decap_3 PHY_2188 ();
 sky130_fd_sc_hd__decap_3 PHY_2189 ();
 sky130_fd_sc_hd__decap_3 PHY_2190 ();
 sky130_fd_sc_hd__decap_3 PHY_2191 ();
 sky130_fd_sc_hd__decap_3 PHY_2192 ();
 sky130_fd_sc_hd__decap_3 PHY_2193 ();
 sky130_fd_sc_hd__decap_3 PHY_2194 ();
 sky130_fd_sc_hd__decap_3 PHY_2195 ();
 sky130_fd_sc_hd__decap_3 PHY_2196 ();
 sky130_fd_sc_hd__decap_3 PHY_2197 ();
 sky130_fd_sc_hd__decap_3 PHY_2198 ();
 sky130_fd_sc_hd__decap_3 PHY_2199 ();
 sky130_fd_sc_hd__decap_3 PHY_2200 ();
 sky130_fd_sc_hd__decap_3 PHY_2201 ();
 sky130_fd_sc_hd__decap_3 PHY_2202 ();
 sky130_fd_sc_hd__decap_3 PHY_2203 ();
 sky130_fd_sc_hd__decap_3 PHY_2204 ();
 sky130_fd_sc_hd__decap_3 PHY_2205 ();
 sky130_fd_sc_hd__decap_3 PHY_2206 ();
 sky130_fd_sc_hd__decap_3 PHY_2207 ();
 sky130_fd_sc_hd__decap_3 PHY_2208 ();
 sky130_fd_sc_hd__decap_3 PHY_2209 ();
 sky130_fd_sc_hd__decap_3 PHY_2210 ();
 sky130_fd_sc_hd__decap_3 PHY_2211 ();
 sky130_fd_sc_hd__decap_3 PHY_2212 ();
 sky130_fd_sc_hd__decap_3 PHY_2213 ();
 sky130_fd_sc_hd__decap_3 PHY_2214 ();
 sky130_fd_sc_hd__decap_3 PHY_2215 ();
 sky130_fd_sc_hd__decap_3 PHY_2216 ();
 sky130_fd_sc_hd__decap_3 PHY_2217 ();
 sky130_fd_sc_hd__decap_3 PHY_2218 ();
 sky130_fd_sc_hd__decap_3 PHY_2219 ();
 sky130_fd_sc_hd__decap_3 PHY_2220 ();
 sky130_fd_sc_hd__decap_3 PHY_2221 ();
 sky130_fd_sc_hd__decap_3 PHY_2222 ();
 sky130_fd_sc_hd__decap_3 PHY_2223 ();
 sky130_fd_sc_hd__decap_3 PHY_2224 ();
 sky130_fd_sc_hd__decap_3 PHY_2225 ();
 sky130_fd_sc_hd__decap_3 PHY_2226 ();
 sky130_fd_sc_hd__decap_3 PHY_2227 ();
 sky130_fd_sc_hd__decap_3 PHY_2228 ();
 sky130_fd_sc_hd__decap_3 PHY_2229 ();
 sky130_fd_sc_hd__decap_3 PHY_2230 ();
 sky130_fd_sc_hd__decap_3 PHY_2231 ();
 sky130_fd_sc_hd__decap_3 PHY_2232 ();
 sky130_fd_sc_hd__decap_3 PHY_2233 ();
 sky130_fd_sc_hd__decap_3 PHY_2234 ();
 sky130_fd_sc_hd__decap_3 PHY_2235 ();
 sky130_fd_sc_hd__decap_3 PHY_2236 ();
 sky130_fd_sc_hd__decap_3 PHY_2237 ();
 sky130_fd_sc_hd__decap_3 PHY_2238 ();
 sky130_fd_sc_hd__decap_3 PHY_2239 ();
 sky130_fd_sc_hd__decap_3 PHY_2240 ();
 sky130_fd_sc_hd__decap_3 PHY_2241 ();
 sky130_fd_sc_hd__decap_3 PHY_2242 ();
 sky130_fd_sc_hd__decap_3 PHY_2243 ();
 sky130_fd_sc_hd__decap_3 PHY_2244 ();
 sky130_fd_sc_hd__decap_3 PHY_2245 ();
 sky130_fd_sc_hd__decap_3 PHY_2246 ();
 sky130_fd_sc_hd__decap_3 PHY_2247 ();
 sky130_fd_sc_hd__decap_3 PHY_2248 ();
 sky130_fd_sc_hd__decap_3 PHY_2249 ();
 sky130_fd_sc_hd__decap_3 PHY_2250 ();
 sky130_fd_sc_hd__decap_3 PHY_2251 ();
 sky130_fd_sc_hd__decap_3 PHY_2252 ();
 sky130_fd_sc_hd__decap_3 PHY_2253 ();
 sky130_fd_sc_hd__decap_3 PHY_2254 ();
 sky130_fd_sc_hd__decap_3 PHY_2255 ();
 sky130_fd_sc_hd__decap_3 PHY_2256 ();
 sky130_fd_sc_hd__decap_3 PHY_2257 ();
 sky130_fd_sc_hd__decap_3 PHY_2258 ();
 sky130_fd_sc_hd__decap_3 PHY_2259 ();
 sky130_fd_sc_hd__decap_3 PHY_2260 ();
 sky130_fd_sc_hd__decap_3 PHY_2261 ();
 sky130_fd_sc_hd__decap_3 PHY_2262 ();
 sky130_fd_sc_hd__decap_3 PHY_2263 ();
 sky130_fd_sc_hd__decap_3 PHY_2264 ();
 sky130_fd_sc_hd__decap_3 PHY_2265 ();
 sky130_fd_sc_hd__decap_3 PHY_2266 ();
 sky130_fd_sc_hd__decap_3 PHY_2267 ();
 sky130_fd_sc_hd__decap_3 PHY_2268 ();
 sky130_fd_sc_hd__decap_3 PHY_2269 ();
 sky130_fd_sc_hd__decap_3 PHY_2270 ();
 sky130_fd_sc_hd__decap_3 PHY_2271 ();
 sky130_fd_sc_hd__decap_3 PHY_2272 ();
 sky130_fd_sc_hd__decap_3 PHY_2273 ();
 sky130_fd_sc_hd__decap_3 PHY_2274 ();
 sky130_fd_sc_hd__decap_3 PHY_2275 ();
 sky130_fd_sc_hd__decap_3 PHY_2276 ();
 sky130_fd_sc_hd__decap_3 PHY_2277 ();
 sky130_fd_sc_hd__decap_3 PHY_2278 ();
 sky130_fd_sc_hd__decap_3 PHY_2279 ();
 sky130_fd_sc_hd__decap_3 PHY_2280 ();
 sky130_fd_sc_hd__decap_3 PHY_2281 ();
 sky130_fd_sc_hd__decap_3 PHY_2282 ();
 sky130_fd_sc_hd__decap_3 PHY_2283 ();
 sky130_fd_sc_hd__decap_3 PHY_2284 ();
 sky130_fd_sc_hd__decap_3 PHY_2285 ();
 sky130_fd_sc_hd__decap_3 PHY_2286 ();
 sky130_fd_sc_hd__decap_3 PHY_2287 ();
 sky130_fd_sc_hd__decap_3 PHY_2288 ();
 sky130_fd_sc_hd__decap_3 PHY_2289 ();
 sky130_fd_sc_hd__decap_3 PHY_2290 ();
 sky130_fd_sc_hd__decap_3 PHY_2291 ();
 sky130_fd_sc_hd__decap_3 PHY_2292 ();
 sky130_fd_sc_hd__decap_3 PHY_2293 ();
 sky130_fd_sc_hd__decap_3 PHY_2294 ();
 sky130_fd_sc_hd__decap_3 PHY_2295 ();
 sky130_fd_sc_hd__decap_3 PHY_2296 ();
 sky130_fd_sc_hd__decap_3 PHY_2297 ();
 sky130_fd_sc_hd__decap_3 PHY_2298 ();
 sky130_fd_sc_hd__decap_3 PHY_2299 ();
 sky130_fd_sc_hd__decap_3 PHY_2300 ();
 sky130_fd_sc_hd__decap_3 PHY_2301 ();
 sky130_fd_sc_hd__decap_3 PHY_2302 ();
 sky130_fd_sc_hd__decap_3 PHY_2303 ();
 sky130_fd_sc_hd__decap_3 PHY_2304 ();
 sky130_fd_sc_hd__decap_3 PHY_2305 ();
 sky130_fd_sc_hd__decap_3 PHY_2306 ();
 sky130_fd_sc_hd__decap_3 PHY_2307 ();
 sky130_fd_sc_hd__decap_3 PHY_2308 ();
 sky130_fd_sc_hd__decap_3 PHY_2309 ();
 sky130_fd_sc_hd__decap_3 PHY_2310 ();
 sky130_fd_sc_hd__decap_3 PHY_2311 ();
 sky130_fd_sc_hd__decap_3 PHY_2312 ();
 sky130_fd_sc_hd__decap_3 PHY_2313 ();
 sky130_fd_sc_hd__decap_3 PHY_2314 ();
 sky130_fd_sc_hd__decap_3 PHY_2315 ();
 sky130_fd_sc_hd__decap_3 PHY_2316 ();
 sky130_fd_sc_hd__decap_3 PHY_2317 ();
 sky130_fd_sc_hd__decap_3 PHY_2318 ();
 sky130_fd_sc_hd__decap_3 PHY_2319 ();
 sky130_fd_sc_hd__decap_3 PHY_2320 ();
 sky130_fd_sc_hd__decap_3 PHY_2321 ();
 sky130_fd_sc_hd__decap_3 PHY_2322 ();
 sky130_fd_sc_hd__decap_3 PHY_2323 ();
 sky130_fd_sc_hd__decap_3 PHY_2324 ();
 sky130_fd_sc_hd__decap_3 PHY_2325 ();
 sky130_fd_sc_hd__decap_3 PHY_2326 ();
 sky130_fd_sc_hd__decap_3 PHY_2327 ();
 sky130_fd_sc_hd__decap_3 PHY_2328 ();
 sky130_fd_sc_hd__decap_3 PHY_2329 ();
 sky130_fd_sc_hd__decap_3 PHY_2330 ();
 sky130_fd_sc_hd__decap_3 PHY_2331 ();
 sky130_fd_sc_hd__decap_3 PHY_2332 ();
 sky130_fd_sc_hd__decap_3 PHY_2333 ();
 sky130_fd_sc_hd__decap_3 PHY_2334 ();
 sky130_fd_sc_hd__decap_3 PHY_2335 ();
 sky130_fd_sc_hd__decap_3 PHY_2336 ();
 sky130_fd_sc_hd__decap_3 PHY_2337 ();
 sky130_fd_sc_hd__decap_3 PHY_2338 ();
 sky130_fd_sc_hd__decap_3 PHY_2339 ();
 sky130_fd_sc_hd__decap_3 PHY_2340 ();
 sky130_fd_sc_hd__decap_3 PHY_2341 ();
 sky130_fd_sc_hd__decap_3 PHY_2342 ();
 sky130_fd_sc_hd__decap_3 PHY_2343 ();
 sky130_fd_sc_hd__decap_3 PHY_2344 ();
 sky130_fd_sc_hd__decap_3 PHY_2345 ();
 sky130_fd_sc_hd__decap_3 PHY_2346 ();
 sky130_fd_sc_hd__decap_3 PHY_2347 ();
 sky130_fd_sc_hd__decap_3 PHY_2348 ();
 sky130_fd_sc_hd__decap_3 PHY_2349 ();
 sky130_fd_sc_hd__decap_3 PHY_2350 ();
 sky130_fd_sc_hd__decap_3 PHY_2351 ();
 sky130_fd_sc_hd__decap_3 PHY_2352 ();
 sky130_fd_sc_hd__decap_3 PHY_2353 ();
 sky130_fd_sc_hd__decap_3 PHY_2354 ();
 sky130_fd_sc_hd__decap_3 PHY_2355 ();
 sky130_fd_sc_hd__decap_3 PHY_2356 ();
 sky130_fd_sc_hd__decap_3 PHY_2357 ();
 sky130_fd_sc_hd__decap_3 PHY_2358 ();
 sky130_fd_sc_hd__decap_3 PHY_2359 ();
 sky130_fd_sc_hd__decap_3 PHY_2360 ();
 sky130_fd_sc_hd__decap_3 PHY_2361 ();
 sky130_fd_sc_hd__decap_3 PHY_2362 ();
 sky130_fd_sc_hd__decap_3 PHY_2363 ();
 sky130_fd_sc_hd__decap_3 PHY_2364 ();
 sky130_fd_sc_hd__decap_3 PHY_2365 ();
 sky130_fd_sc_hd__decap_3 PHY_2366 ();
 sky130_fd_sc_hd__decap_3 PHY_2367 ();
 sky130_fd_sc_hd__decap_3 PHY_2368 ();
 sky130_fd_sc_hd__decap_3 PHY_2369 ();
 sky130_fd_sc_hd__decap_3 PHY_2370 ();
 sky130_fd_sc_hd__decap_3 PHY_2371 ();
 sky130_fd_sc_hd__decap_3 PHY_2372 ();
 sky130_fd_sc_hd__decap_3 PHY_2373 ();
 sky130_fd_sc_hd__decap_3 PHY_2374 ();
 sky130_fd_sc_hd__decap_3 PHY_2375 ();
 sky130_fd_sc_hd__decap_3 PHY_2376 ();
 sky130_fd_sc_hd__decap_3 PHY_2377 ();
 sky130_fd_sc_hd__decap_3 PHY_2378 ();
 sky130_fd_sc_hd__decap_3 PHY_2379 ();
 sky130_fd_sc_hd__decap_3 PHY_2380 ();
 sky130_fd_sc_hd__decap_3 PHY_2381 ();
 sky130_fd_sc_hd__decap_3 PHY_2382 ();
 sky130_fd_sc_hd__decap_3 PHY_2383 ();
 sky130_fd_sc_hd__decap_3 PHY_2384 ();
 sky130_fd_sc_hd__decap_3 PHY_2385 ();
 sky130_fd_sc_hd__decap_3 PHY_2386 ();
 sky130_fd_sc_hd__decap_3 PHY_2387 ();
 sky130_fd_sc_hd__decap_3 PHY_2388 ();
 sky130_fd_sc_hd__decap_3 PHY_2389 ();
 sky130_fd_sc_hd__decap_3 PHY_2390 ();
 sky130_fd_sc_hd__decap_3 PHY_2391 ();
 sky130_fd_sc_hd__decap_3 PHY_2392 ();
 sky130_fd_sc_hd__decap_3 PHY_2393 ();
 sky130_fd_sc_hd__decap_3 PHY_2394 ();
 sky130_fd_sc_hd__decap_3 PHY_2395 ();
 sky130_fd_sc_hd__decap_3 PHY_2396 ();
 sky130_fd_sc_hd__decap_3 PHY_2397 ();
 sky130_fd_sc_hd__decap_3 PHY_2398 ();
 sky130_fd_sc_hd__decap_3 PHY_2399 ();
 sky130_fd_sc_hd__decap_3 PHY_2400 ();
 sky130_fd_sc_hd__decap_3 PHY_2401 ();
 sky130_fd_sc_hd__decap_3 PHY_2402 ();
 sky130_fd_sc_hd__decap_3 PHY_2403 ();
 sky130_fd_sc_hd__decap_3 PHY_2404 ();
 sky130_fd_sc_hd__decap_3 PHY_2405 ();
 sky130_fd_sc_hd__decap_3 PHY_2406 ();
 sky130_fd_sc_hd__decap_3 PHY_2407 ();
 sky130_fd_sc_hd__decap_3 PHY_2408 ();
 sky130_fd_sc_hd__decap_3 PHY_2409 ();
 sky130_fd_sc_hd__decap_3 PHY_2410 ();
 sky130_fd_sc_hd__decap_3 PHY_2411 ();
 sky130_fd_sc_hd__decap_3 PHY_2412 ();
 sky130_fd_sc_hd__decap_3 PHY_2413 ();
 sky130_fd_sc_hd__decap_3 PHY_2414 ();
 sky130_fd_sc_hd__decap_3 PHY_2415 ();
 sky130_fd_sc_hd__decap_3 PHY_2416 ();
 sky130_fd_sc_hd__decap_3 PHY_2417 ();
 sky130_fd_sc_hd__decap_3 PHY_2418 ();
 sky130_fd_sc_hd__decap_3 PHY_2419 ();
 sky130_fd_sc_hd__decap_3 PHY_2420 ();
 sky130_fd_sc_hd__decap_3 PHY_2421 ();
 sky130_fd_sc_hd__decap_3 PHY_2422 ();
 sky130_fd_sc_hd__decap_3 PHY_2423 ();
 sky130_fd_sc_hd__decap_3 PHY_2424 ();
 sky130_fd_sc_hd__decap_3 PHY_2425 ();
 sky130_fd_sc_hd__decap_3 PHY_2426 ();
 sky130_fd_sc_hd__decap_3 PHY_2427 ();
 sky130_fd_sc_hd__decap_3 PHY_2428 ();
 sky130_fd_sc_hd__decap_3 PHY_2429 ();
 sky130_fd_sc_hd__decap_3 PHY_2430 ();
 sky130_fd_sc_hd__decap_3 PHY_2431 ();
 sky130_fd_sc_hd__decap_3 PHY_2432 ();
 sky130_fd_sc_hd__decap_3 PHY_2433 ();
 sky130_fd_sc_hd__decap_3 PHY_2434 ();
 sky130_fd_sc_hd__decap_3 PHY_2435 ();
 sky130_fd_sc_hd__decap_3 PHY_2436 ();
 sky130_fd_sc_hd__decap_3 PHY_2437 ();
 sky130_fd_sc_hd__decap_3 PHY_2438 ();
 sky130_fd_sc_hd__decap_3 PHY_2439 ();
 sky130_fd_sc_hd__decap_3 PHY_2440 ();
 sky130_fd_sc_hd__decap_3 PHY_2441 ();
 sky130_fd_sc_hd__decap_3 PHY_2442 ();
 sky130_fd_sc_hd__decap_3 PHY_2443 ();
 sky130_fd_sc_hd__decap_3 PHY_2444 ();
 sky130_fd_sc_hd__decap_3 PHY_2445 ();
 sky130_fd_sc_hd__decap_3 PHY_2446 ();
 sky130_fd_sc_hd__decap_3 PHY_2447 ();
 sky130_fd_sc_hd__decap_3 PHY_2448 ();
 sky130_fd_sc_hd__decap_3 PHY_2449 ();
 sky130_fd_sc_hd__decap_3 PHY_2450 ();
 sky130_fd_sc_hd__decap_3 PHY_2451 ();
 sky130_fd_sc_hd__decap_3 PHY_2452 ();
 sky130_fd_sc_hd__decap_3 PHY_2453 ();
 sky130_fd_sc_hd__decap_3 PHY_2454 ();
 sky130_fd_sc_hd__decap_3 PHY_2455 ();
 sky130_fd_sc_hd__decap_3 PHY_2456 ();
 sky130_fd_sc_hd__decap_3 PHY_2457 ();
 sky130_fd_sc_hd__decap_3 PHY_2458 ();
 sky130_fd_sc_hd__decap_3 PHY_2459 ();
 sky130_fd_sc_hd__decap_3 PHY_2460 ();
 sky130_fd_sc_hd__decap_3 PHY_2461 ();
 sky130_fd_sc_hd__decap_3 PHY_2462 ();
 sky130_fd_sc_hd__decap_3 PHY_2463 ();
 sky130_fd_sc_hd__decap_3 PHY_2464 ();
 sky130_fd_sc_hd__decap_3 PHY_2465 ();
 sky130_fd_sc_hd__decap_3 PHY_2466 ();
 sky130_fd_sc_hd__decap_3 PHY_2467 ();
 sky130_fd_sc_hd__decap_3 PHY_2468 ();
 sky130_fd_sc_hd__decap_3 PHY_2469 ();
 sky130_fd_sc_hd__decap_3 PHY_2470 ();
 sky130_fd_sc_hd__decap_3 PHY_2471 ();
 sky130_fd_sc_hd__decap_3 PHY_2472 ();
 sky130_fd_sc_hd__decap_3 PHY_2473 ();
 sky130_fd_sc_hd__decap_3 PHY_2474 ();
 sky130_fd_sc_hd__decap_3 PHY_2475 ();
 sky130_fd_sc_hd__decap_3 PHY_2476 ();
 sky130_fd_sc_hd__decap_3 PHY_2477 ();
 sky130_fd_sc_hd__decap_3 PHY_2478 ();
 sky130_fd_sc_hd__decap_3 PHY_2479 ();
 sky130_fd_sc_hd__decap_3 PHY_2480 ();
 sky130_fd_sc_hd__decap_3 PHY_2481 ();
 sky130_fd_sc_hd__decap_3 PHY_2482 ();
 sky130_fd_sc_hd__decap_3 PHY_2483 ();
 sky130_fd_sc_hd__decap_3 PHY_2484 ();
 sky130_fd_sc_hd__decap_3 PHY_2485 ();
 sky130_fd_sc_hd__decap_3 PHY_2486 ();
 sky130_fd_sc_hd__decap_3 PHY_2487 ();
 sky130_fd_sc_hd__decap_3 PHY_2488 ();
 sky130_fd_sc_hd__decap_3 PHY_2489 ();
 sky130_fd_sc_hd__decap_3 PHY_2490 ();
 sky130_fd_sc_hd__decap_3 PHY_2491 ();
 sky130_fd_sc_hd__decap_3 PHY_2492 ();
 sky130_fd_sc_hd__decap_3 PHY_2493 ();
 sky130_fd_sc_hd__decap_3 PHY_2494 ();
 sky130_fd_sc_hd__decap_3 PHY_2495 ();
 sky130_fd_sc_hd__decap_3 PHY_2496 ();
 sky130_fd_sc_hd__decap_3 PHY_2497 ();
 sky130_fd_sc_hd__decap_3 PHY_2498 ();
 sky130_fd_sc_hd__decap_3 PHY_2499 ();
 sky130_fd_sc_hd__decap_3 PHY_2500 ();
 sky130_fd_sc_hd__decap_3 PHY_2501 ();
 sky130_fd_sc_hd__decap_3 PHY_2502 ();
 sky130_fd_sc_hd__decap_3 PHY_2503 ();
 sky130_fd_sc_hd__decap_3 PHY_2504 ();
 sky130_fd_sc_hd__decap_3 PHY_2505 ();
 sky130_fd_sc_hd__decap_3 PHY_2506 ();
 sky130_fd_sc_hd__decap_3 PHY_2507 ();
 sky130_fd_sc_hd__decap_3 PHY_2508 ();
 sky130_fd_sc_hd__decap_3 PHY_2509 ();
 sky130_fd_sc_hd__decap_3 PHY_2510 ();
 sky130_fd_sc_hd__decap_3 PHY_2511 ();
 sky130_fd_sc_hd__decap_3 PHY_2512 ();
 sky130_fd_sc_hd__decap_3 PHY_2513 ();
 sky130_fd_sc_hd__decap_3 PHY_2514 ();
 sky130_fd_sc_hd__decap_3 PHY_2515 ();
 sky130_fd_sc_hd__decap_3 PHY_2516 ();
 sky130_fd_sc_hd__decap_3 PHY_2517 ();
 sky130_fd_sc_hd__decap_3 PHY_2518 ();
 sky130_fd_sc_hd__decap_3 PHY_2519 ();
 sky130_fd_sc_hd__decap_3 PHY_2520 ();
 sky130_fd_sc_hd__decap_3 PHY_2521 ();
 sky130_fd_sc_hd__decap_3 PHY_2522 ();
 sky130_fd_sc_hd__decap_3 PHY_2523 ();
 sky130_fd_sc_hd__decap_3 PHY_2524 ();
 sky130_fd_sc_hd__decap_3 PHY_2525 ();
 sky130_fd_sc_hd__decap_3 PHY_2526 ();
 sky130_fd_sc_hd__decap_3 PHY_2527 ();
 sky130_fd_sc_hd__decap_3 PHY_2528 ();
 sky130_fd_sc_hd__decap_3 PHY_2529 ();
 sky130_fd_sc_hd__decap_3 PHY_2530 ();
 sky130_fd_sc_hd__decap_3 PHY_2531 ();
 sky130_fd_sc_hd__decap_3 PHY_2532 ();
 sky130_fd_sc_hd__decap_3 PHY_2533 ();
 sky130_fd_sc_hd__decap_3 PHY_2534 ();
 sky130_fd_sc_hd__decap_3 PHY_2535 ();
 sky130_fd_sc_hd__decap_3 PHY_2536 ();
 sky130_fd_sc_hd__decap_3 PHY_2537 ();
 sky130_fd_sc_hd__decap_3 PHY_2538 ();
 sky130_fd_sc_hd__decap_3 PHY_2539 ();
 sky130_fd_sc_hd__decap_3 PHY_2540 ();
 sky130_fd_sc_hd__decap_3 PHY_2541 ();
 sky130_fd_sc_hd__decap_3 PHY_2542 ();
 sky130_fd_sc_hd__decap_3 PHY_2543 ();
 sky130_fd_sc_hd__decap_3 PHY_2544 ();
 sky130_fd_sc_hd__decap_3 PHY_2545 ();
 sky130_fd_sc_hd__decap_3 PHY_2546 ();
 sky130_fd_sc_hd__decap_3 PHY_2547 ();
 sky130_fd_sc_hd__decap_3 PHY_2548 ();
 sky130_fd_sc_hd__decap_3 PHY_2549 ();
 sky130_fd_sc_hd__decap_3 PHY_2550 ();
 sky130_fd_sc_hd__decap_3 PHY_2551 ();
 sky130_fd_sc_hd__decap_3 PHY_2552 ();
 sky130_fd_sc_hd__decap_3 PHY_2553 ();
 sky130_fd_sc_hd__decap_3 PHY_2554 ();
 sky130_fd_sc_hd__decap_3 PHY_2555 ();
 sky130_fd_sc_hd__decap_3 PHY_2556 ();
 sky130_fd_sc_hd__decap_3 PHY_2557 ();
 sky130_fd_sc_hd__decap_3 PHY_2558 ();
 sky130_fd_sc_hd__decap_3 PHY_2559 ();
 sky130_fd_sc_hd__decap_3 PHY_2560 ();
 sky130_fd_sc_hd__decap_3 PHY_2561 ();
 sky130_fd_sc_hd__decap_3 PHY_2562 ();
 sky130_fd_sc_hd__decap_3 PHY_2563 ();
 sky130_fd_sc_hd__decap_3 PHY_2564 ();
 sky130_fd_sc_hd__decap_3 PHY_2565 ();
 sky130_fd_sc_hd__decap_3 PHY_2566 ();
 sky130_fd_sc_hd__decap_3 PHY_2567 ();
 sky130_fd_sc_hd__decap_3 PHY_2568 ();
 sky130_fd_sc_hd__decap_3 PHY_2569 ();
 sky130_fd_sc_hd__decap_3 PHY_2570 ();
 sky130_fd_sc_hd__decap_3 PHY_2571 ();
 sky130_fd_sc_hd__decap_3 PHY_2572 ();
 sky130_fd_sc_hd__decap_3 PHY_2573 ();
 sky130_fd_sc_hd__decap_3 PHY_2574 ();
 sky130_fd_sc_hd__decap_3 PHY_2575 ();
 sky130_fd_sc_hd__decap_3 PHY_2576 ();
 sky130_fd_sc_hd__decap_3 PHY_2577 ();
 sky130_fd_sc_hd__decap_3 PHY_2578 ();
 sky130_fd_sc_hd__decap_3 PHY_2579 ();
 sky130_fd_sc_hd__decap_3 PHY_2580 ();
 sky130_fd_sc_hd__decap_3 PHY_2581 ();
 sky130_fd_sc_hd__decap_3 PHY_2582 ();
 sky130_fd_sc_hd__decap_3 PHY_2583 ();
 sky130_fd_sc_hd__decap_3 PHY_2584 ();
 sky130_fd_sc_hd__decap_3 PHY_2585 ();
 sky130_fd_sc_hd__decap_3 PHY_2586 ();
 sky130_fd_sc_hd__decap_3 PHY_2587 ();
 sky130_fd_sc_hd__decap_3 PHY_2588 ();
 sky130_fd_sc_hd__decap_3 PHY_2589 ();
 sky130_fd_sc_hd__decap_3 PHY_2590 ();
 sky130_fd_sc_hd__decap_3 PHY_2591 ();
 sky130_fd_sc_hd__decap_3 PHY_2592 ();
 sky130_fd_sc_hd__decap_3 PHY_2593 ();
 sky130_fd_sc_hd__decap_3 PHY_2594 ();
 sky130_fd_sc_hd__decap_3 PHY_2595 ();
 sky130_fd_sc_hd__decap_3 PHY_2596 ();
 sky130_fd_sc_hd__decap_3 PHY_2597 ();
 sky130_fd_sc_hd__decap_3 PHY_2598 ();
 sky130_fd_sc_hd__decap_3 PHY_2599 ();
 sky130_fd_sc_hd__decap_3 PHY_2600 ();
 sky130_fd_sc_hd__decap_3 PHY_2601 ();
 sky130_fd_sc_hd__decap_3 PHY_2602 ();
 sky130_fd_sc_hd__decap_3 PHY_2603 ();
 sky130_fd_sc_hd__decap_3 PHY_2604 ();
 sky130_fd_sc_hd__decap_3 PHY_2605 ();
 sky130_fd_sc_hd__decap_3 PHY_2606 ();
 sky130_fd_sc_hd__decap_3 PHY_2607 ();
 sky130_fd_sc_hd__decap_3 PHY_2608 ();
 sky130_fd_sc_hd__decap_3 PHY_2609 ();
 sky130_fd_sc_hd__decap_3 PHY_2610 ();
 sky130_fd_sc_hd__decap_3 PHY_2611 ();
 sky130_fd_sc_hd__decap_3 PHY_2612 ();
 sky130_fd_sc_hd__decap_3 PHY_2613 ();
 sky130_fd_sc_hd__decap_3 PHY_2614 ();
 sky130_fd_sc_hd__decap_3 PHY_2615 ();
 sky130_fd_sc_hd__decap_3 PHY_2616 ();
 sky130_fd_sc_hd__decap_3 PHY_2617 ();
 sky130_fd_sc_hd__decap_3 PHY_2618 ();
 sky130_fd_sc_hd__decap_3 PHY_2619 ();
 sky130_fd_sc_hd__decap_3 PHY_2620 ();
 sky130_fd_sc_hd__decap_3 PHY_2621 ();
 sky130_fd_sc_hd__decap_3 PHY_2622 ();
 sky130_fd_sc_hd__decap_3 PHY_2623 ();
 sky130_fd_sc_hd__decap_3 PHY_2624 ();
 sky130_fd_sc_hd__decap_3 PHY_2625 ();
 sky130_fd_sc_hd__decap_3 PHY_2626 ();
 sky130_fd_sc_hd__decap_3 PHY_2627 ();
 sky130_fd_sc_hd__decap_3 PHY_2628 ();
 sky130_fd_sc_hd__decap_3 PHY_2629 ();
 sky130_fd_sc_hd__decap_3 PHY_2630 ();
 sky130_fd_sc_hd__decap_3 PHY_2631 ();
 sky130_fd_sc_hd__decap_3 PHY_2632 ();
 sky130_fd_sc_hd__decap_3 PHY_2633 ();
 sky130_fd_sc_hd__decap_3 PHY_2634 ();
 sky130_fd_sc_hd__decap_3 PHY_2635 ();
 sky130_fd_sc_hd__decap_3 PHY_2636 ();
 sky130_fd_sc_hd__decap_3 PHY_2637 ();
 sky130_fd_sc_hd__decap_3 PHY_2638 ();
 sky130_fd_sc_hd__decap_3 PHY_2639 ();
 sky130_fd_sc_hd__decap_3 PHY_2640 ();
 sky130_fd_sc_hd__decap_3 PHY_2641 ();
 sky130_fd_sc_hd__decap_3 PHY_2642 ();
 sky130_fd_sc_hd__decap_3 PHY_2643 ();
 sky130_fd_sc_hd__decap_3 PHY_2644 ();
 sky130_fd_sc_hd__decap_3 PHY_2645 ();
 sky130_fd_sc_hd__decap_3 PHY_2646 ();
 sky130_fd_sc_hd__decap_3 PHY_2647 ();
 sky130_fd_sc_hd__decap_3 PHY_2648 ();
 sky130_fd_sc_hd__decap_3 PHY_2649 ();
 sky130_fd_sc_hd__decap_3 PHY_2650 ();
 sky130_fd_sc_hd__decap_3 PHY_2651 ();
 sky130_fd_sc_hd__decap_3 PHY_2652 ();
 sky130_fd_sc_hd__decap_3 PHY_2653 ();
 sky130_fd_sc_hd__decap_3 PHY_2654 ();
 sky130_fd_sc_hd__decap_3 PHY_2655 ();
 sky130_fd_sc_hd__decap_3 PHY_2656 ();
 sky130_fd_sc_hd__decap_3 PHY_2657 ();
 sky130_fd_sc_hd__decap_3 PHY_2658 ();
 sky130_fd_sc_hd__decap_3 PHY_2659 ();
 sky130_fd_sc_hd__decap_3 PHY_2660 ();
 sky130_fd_sc_hd__decap_3 PHY_2661 ();
 sky130_fd_sc_hd__decap_3 PHY_2662 ();
 sky130_fd_sc_hd__decap_3 PHY_2663 ();
 sky130_fd_sc_hd__decap_3 PHY_2664 ();
 sky130_fd_sc_hd__decap_3 PHY_2665 ();
 sky130_fd_sc_hd__decap_3 PHY_2666 ();
 sky130_fd_sc_hd__decap_3 PHY_2667 ();
 sky130_fd_sc_hd__decap_3 PHY_2668 ();
 sky130_fd_sc_hd__decap_3 PHY_2669 ();
 sky130_fd_sc_hd__decap_3 PHY_2670 ();
 sky130_fd_sc_hd__decap_3 PHY_2671 ();
 sky130_fd_sc_hd__decap_3 PHY_2672 ();
 sky130_fd_sc_hd__decap_3 PHY_2673 ();
 sky130_fd_sc_hd__decap_3 PHY_2674 ();
 sky130_fd_sc_hd__decap_3 PHY_2675 ();
 sky130_fd_sc_hd__decap_3 PHY_2676 ();
 sky130_fd_sc_hd__decap_3 PHY_2677 ();
 sky130_fd_sc_hd__decap_3 PHY_2678 ();
 sky130_fd_sc_hd__decap_3 PHY_2679 ();
 sky130_fd_sc_hd__decap_3 PHY_2680 ();
 sky130_fd_sc_hd__decap_3 PHY_2681 ();
 sky130_fd_sc_hd__decap_3 PHY_2682 ();
 sky130_fd_sc_hd__decap_3 PHY_2683 ();
 sky130_fd_sc_hd__decap_3 PHY_2684 ();
 sky130_fd_sc_hd__decap_3 PHY_2685 ();
 sky130_fd_sc_hd__decap_3 PHY_2686 ();
 sky130_fd_sc_hd__decap_3 PHY_2687 ();
 sky130_fd_sc_hd__decap_3 PHY_2688 ();
 sky130_fd_sc_hd__decap_3 PHY_2689 ();
 sky130_fd_sc_hd__decap_3 PHY_2690 ();
 sky130_fd_sc_hd__decap_3 PHY_2691 ();
 sky130_fd_sc_hd__decap_3 PHY_2692 ();
 sky130_fd_sc_hd__decap_3 PHY_2693 ();
 sky130_fd_sc_hd__decap_3 PHY_2694 ();
 sky130_fd_sc_hd__decap_3 PHY_2695 ();
 sky130_fd_sc_hd__decap_3 PHY_2696 ();
 sky130_fd_sc_hd__decap_3 PHY_2697 ();
 sky130_fd_sc_hd__decap_3 PHY_2698 ();
 sky130_fd_sc_hd__decap_3 PHY_2699 ();
 sky130_fd_sc_hd__decap_3 PHY_2700 ();
 sky130_fd_sc_hd__decap_3 PHY_2701 ();
 sky130_fd_sc_hd__decap_3 PHY_2702 ();
 sky130_fd_sc_hd__decap_3 PHY_2703 ();
 sky130_fd_sc_hd__decap_3 PHY_2704 ();
 sky130_fd_sc_hd__decap_3 PHY_2705 ();
 sky130_fd_sc_hd__decap_3 PHY_2706 ();
 sky130_fd_sc_hd__decap_3 PHY_2707 ();
 sky130_fd_sc_hd__decap_3 PHY_2708 ();
 sky130_fd_sc_hd__decap_3 PHY_2709 ();
 sky130_fd_sc_hd__decap_3 PHY_2710 ();
 sky130_fd_sc_hd__decap_3 PHY_2711 ();
 sky130_fd_sc_hd__decap_3 PHY_2712 ();
 sky130_fd_sc_hd__decap_3 PHY_2713 ();
 sky130_fd_sc_hd__decap_3 PHY_2714 ();
 sky130_fd_sc_hd__decap_3 PHY_2715 ();
 sky130_fd_sc_hd__decap_3 PHY_2716 ();
 sky130_fd_sc_hd__decap_3 PHY_2717 ();
 sky130_fd_sc_hd__decap_3 PHY_2718 ();
 sky130_fd_sc_hd__decap_3 PHY_2719 ();
 sky130_fd_sc_hd__decap_3 PHY_2720 ();
 sky130_fd_sc_hd__decap_3 PHY_2721 ();
 sky130_fd_sc_hd__decap_3 PHY_2722 ();
 sky130_fd_sc_hd__decap_3 PHY_2723 ();
 sky130_fd_sc_hd__decap_3 PHY_2724 ();
 sky130_fd_sc_hd__decap_3 PHY_2725 ();
 sky130_fd_sc_hd__decap_3 PHY_2726 ();
 sky130_fd_sc_hd__decap_3 PHY_2727 ();
 sky130_fd_sc_hd__decap_3 PHY_2728 ();
 sky130_fd_sc_hd__decap_3 PHY_2729 ();
 sky130_fd_sc_hd__decap_3 PHY_2730 ();
 sky130_fd_sc_hd__decap_3 PHY_2731 ();
 sky130_fd_sc_hd__decap_3 PHY_2732 ();
 sky130_fd_sc_hd__decap_3 PHY_2733 ();
 sky130_fd_sc_hd__decap_3 PHY_2734 ();
 sky130_fd_sc_hd__decap_3 PHY_2735 ();
 sky130_fd_sc_hd__decap_3 PHY_2736 ();
 sky130_fd_sc_hd__decap_3 PHY_2737 ();
 sky130_fd_sc_hd__decap_3 PHY_2738 ();
 sky130_fd_sc_hd__decap_3 PHY_2739 ();
 sky130_fd_sc_hd__decap_3 PHY_2740 ();
 sky130_fd_sc_hd__decap_3 PHY_2741 ();
 sky130_fd_sc_hd__decap_3 PHY_2742 ();
 sky130_fd_sc_hd__decap_3 PHY_2743 ();
 sky130_fd_sc_hd__decap_3 PHY_2744 ();
 sky130_fd_sc_hd__decap_3 PHY_2745 ();
 sky130_fd_sc_hd__decap_3 PHY_2746 ();
 sky130_fd_sc_hd__decap_3 PHY_2747 ();
 sky130_fd_sc_hd__decap_3 PHY_2748 ();
 sky130_fd_sc_hd__decap_3 PHY_2749 ();
 sky130_fd_sc_hd__decap_3 PHY_2750 ();
 sky130_fd_sc_hd__decap_3 PHY_2751 ();
 sky130_fd_sc_hd__decap_3 PHY_2752 ();
 sky130_fd_sc_hd__decap_3 PHY_2753 ();
 sky130_fd_sc_hd__decap_3 PHY_2754 ();
 sky130_fd_sc_hd__decap_3 PHY_2755 ();
 sky130_fd_sc_hd__decap_3 PHY_2756 ();
 sky130_fd_sc_hd__decap_3 PHY_2757 ();
 sky130_fd_sc_hd__decap_3 PHY_2758 ();
 sky130_fd_sc_hd__decap_3 PHY_2759 ();
 sky130_fd_sc_hd__decap_3 PHY_2760 ();
 sky130_fd_sc_hd__decap_3 PHY_2761 ();
 sky130_fd_sc_hd__decap_3 PHY_2762 ();
 sky130_fd_sc_hd__decap_3 PHY_2763 ();
 sky130_fd_sc_hd__decap_3 PHY_2764 ();
 sky130_fd_sc_hd__decap_3 PHY_2765 ();
 sky130_fd_sc_hd__decap_3 PHY_2766 ();
 sky130_fd_sc_hd__decap_3 PHY_2767 ();
 sky130_fd_sc_hd__decap_3 PHY_2768 ();
 sky130_fd_sc_hd__decap_3 PHY_2769 ();
 sky130_fd_sc_hd__decap_3 PHY_2770 ();
 sky130_fd_sc_hd__decap_3 PHY_2771 ();
 sky130_fd_sc_hd__decap_3 PHY_2772 ();
 sky130_fd_sc_hd__decap_3 PHY_2773 ();
 sky130_fd_sc_hd__decap_3 PHY_2774 ();
 sky130_fd_sc_hd__decap_3 PHY_2775 ();
 sky130_fd_sc_hd__decap_3 PHY_2776 ();
 sky130_fd_sc_hd__decap_3 PHY_2777 ();
 sky130_fd_sc_hd__decap_3 PHY_2778 ();
 sky130_fd_sc_hd__decap_3 PHY_2779 ();
 sky130_fd_sc_hd__decap_3 PHY_2780 ();
 sky130_fd_sc_hd__decap_3 PHY_2781 ();
 sky130_fd_sc_hd__decap_3 PHY_2782 ();
 sky130_fd_sc_hd__decap_3 PHY_2783 ();
 sky130_fd_sc_hd__decap_3 PHY_2784 ();
 sky130_fd_sc_hd__decap_3 PHY_2785 ();
 sky130_fd_sc_hd__decap_3 PHY_2786 ();
 sky130_fd_sc_hd__decap_3 PHY_2787 ();
 sky130_fd_sc_hd__decap_3 PHY_2788 ();
 sky130_fd_sc_hd__decap_3 PHY_2789 ();
 sky130_fd_sc_hd__decap_3 PHY_2790 ();
 sky130_fd_sc_hd__decap_3 PHY_2791 ();
 sky130_fd_sc_hd__decap_3 PHY_2792 ();
 sky130_fd_sc_hd__decap_3 PHY_2793 ();
 sky130_fd_sc_hd__decap_3 PHY_2794 ();
 sky130_fd_sc_hd__decap_3 PHY_2795 ();
 sky130_fd_sc_hd__decap_3 PHY_2796 ();
 sky130_fd_sc_hd__decap_3 PHY_2797 ();
 sky130_fd_sc_hd__decap_3 PHY_2798 ();
 sky130_fd_sc_hd__decap_3 PHY_2799 ();
 sky130_fd_sc_hd__decap_3 PHY_2800 ();
 sky130_fd_sc_hd__decap_3 PHY_2801 ();
 sky130_fd_sc_hd__decap_3 PHY_2802 ();
 sky130_fd_sc_hd__decap_3 PHY_2803 ();
 sky130_fd_sc_hd__decap_3 PHY_2804 ();
 sky130_fd_sc_hd__decap_3 PHY_2805 ();
 sky130_fd_sc_hd__decap_3 PHY_2806 ();
 sky130_fd_sc_hd__decap_3 PHY_2807 ();
 sky130_fd_sc_hd__decap_3 PHY_2808 ();
 sky130_fd_sc_hd__decap_3 PHY_2809 ();
 sky130_fd_sc_hd__decap_3 PHY_2810 ();
 sky130_fd_sc_hd__decap_3 PHY_2811 ();
 sky130_fd_sc_hd__decap_3 PHY_2812 ();
 sky130_fd_sc_hd__decap_3 PHY_2813 ();
 sky130_fd_sc_hd__decap_3 PHY_2814 ();
 sky130_fd_sc_hd__decap_3 PHY_2815 ();
 sky130_fd_sc_hd__decap_3 PHY_2816 ();
 sky130_fd_sc_hd__decap_3 PHY_2817 ();
 sky130_fd_sc_hd__decap_3 PHY_2818 ();
 sky130_fd_sc_hd__decap_3 PHY_2819 ();
 sky130_fd_sc_hd__decap_3 PHY_2820 ();
 sky130_fd_sc_hd__decap_3 PHY_2821 ();
 sky130_fd_sc_hd__decap_3 PHY_2822 ();
 sky130_fd_sc_hd__decap_3 PHY_2823 ();
 sky130_fd_sc_hd__decap_3 PHY_2824 ();
 sky130_fd_sc_hd__decap_3 PHY_2825 ();
 sky130_fd_sc_hd__decap_3 PHY_2826 ();
 sky130_fd_sc_hd__decap_3 PHY_2827 ();
 sky130_fd_sc_hd__decap_3 PHY_2828 ();
 sky130_fd_sc_hd__decap_3 PHY_2829 ();
 sky130_fd_sc_hd__decap_3 PHY_2830 ();
 sky130_fd_sc_hd__decap_3 PHY_2831 ();
 sky130_fd_sc_hd__decap_3 PHY_2832 ();
 sky130_fd_sc_hd__decap_3 PHY_2833 ();
 sky130_fd_sc_hd__decap_3 PHY_2834 ();
 sky130_fd_sc_hd__decap_3 PHY_2835 ();
 sky130_fd_sc_hd__decap_3 PHY_2836 ();
 sky130_fd_sc_hd__decap_3 PHY_2837 ();
 sky130_fd_sc_hd__decap_3 PHY_2838 ();
 sky130_fd_sc_hd__decap_3 PHY_2839 ();
 sky130_fd_sc_hd__decap_3 PHY_2840 ();
 sky130_fd_sc_hd__decap_3 PHY_2841 ();
 sky130_fd_sc_hd__decap_3 PHY_2842 ();
 sky130_fd_sc_hd__decap_3 PHY_2843 ();
 sky130_fd_sc_hd__decap_3 PHY_2844 ();
 sky130_fd_sc_hd__decap_3 PHY_2845 ();
 sky130_fd_sc_hd__decap_3 PHY_2846 ();
 sky130_fd_sc_hd__decap_3 PHY_2847 ();
 sky130_fd_sc_hd__decap_3 PHY_2848 ();
 sky130_fd_sc_hd__decap_3 PHY_2849 ();
 sky130_fd_sc_hd__decap_3 PHY_2850 ();
 sky130_fd_sc_hd__decap_3 PHY_2851 ();
 sky130_fd_sc_hd__decap_3 PHY_2852 ();
 sky130_fd_sc_hd__decap_3 PHY_2853 ();
 sky130_fd_sc_hd__decap_3 PHY_2854 ();
 sky130_fd_sc_hd__decap_3 PHY_2855 ();
 sky130_fd_sc_hd__decap_3 PHY_2856 ();
 sky130_fd_sc_hd__decap_3 PHY_2857 ();
 sky130_fd_sc_hd__decap_3 PHY_2858 ();
 sky130_fd_sc_hd__decap_3 PHY_2859 ();
 sky130_fd_sc_hd__decap_3 PHY_2860 ();
 sky130_fd_sc_hd__decap_3 PHY_2861 ();
 sky130_fd_sc_hd__decap_3 PHY_2862 ();
 sky130_fd_sc_hd__decap_3 PHY_2863 ();
 sky130_fd_sc_hd__decap_3 PHY_2864 ();
 sky130_fd_sc_hd__decap_3 PHY_2865 ();
 sky130_fd_sc_hd__decap_3 PHY_2866 ();
 sky130_fd_sc_hd__decap_3 PHY_2867 ();
 sky130_fd_sc_hd__decap_3 PHY_2868 ();
 sky130_fd_sc_hd__decap_3 PHY_2869 ();
 sky130_fd_sc_hd__decap_3 PHY_2870 ();
 sky130_fd_sc_hd__decap_3 PHY_2871 ();
 sky130_fd_sc_hd__decap_3 PHY_2872 ();
 sky130_fd_sc_hd__decap_3 PHY_2873 ();
 sky130_fd_sc_hd__decap_3 PHY_2874 ();
 sky130_fd_sc_hd__decap_3 PHY_2875 ();
 sky130_fd_sc_hd__decap_3 PHY_2876 ();
 sky130_fd_sc_hd__decap_3 PHY_2877 ();
 sky130_fd_sc_hd__decap_3 PHY_2878 ();
 sky130_fd_sc_hd__decap_3 PHY_2879 ();
 sky130_fd_sc_hd__decap_3 PHY_2880 ();
 sky130_fd_sc_hd__decap_3 PHY_2881 ();
 sky130_fd_sc_hd__decap_3 PHY_2882 ();
 sky130_fd_sc_hd__decap_3 PHY_2883 ();
 sky130_fd_sc_hd__decap_3 PHY_2884 ();
 sky130_fd_sc_hd__decap_3 PHY_2885 ();
 sky130_fd_sc_hd__decap_3 PHY_2886 ();
 sky130_fd_sc_hd__decap_3 PHY_2887 ();
 sky130_fd_sc_hd__decap_3 PHY_2888 ();
 sky130_fd_sc_hd__decap_3 PHY_2889 ();
 sky130_fd_sc_hd__decap_3 PHY_2890 ();
 sky130_fd_sc_hd__decap_3 PHY_2891 ();
 sky130_fd_sc_hd__decap_3 PHY_2892 ();
 sky130_fd_sc_hd__decap_3 PHY_2893 ();
 sky130_fd_sc_hd__decap_3 PHY_2894 ();
 sky130_fd_sc_hd__decap_3 PHY_2895 ();
 sky130_fd_sc_hd__decap_3 PHY_2896 ();
 sky130_fd_sc_hd__decap_3 PHY_2897 ();
 sky130_fd_sc_hd__decap_3 PHY_2898 ();
 sky130_fd_sc_hd__decap_3 PHY_2899 ();
 sky130_fd_sc_hd__decap_3 PHY_2900 ();
 sky130_fd_sc_hd__decap_3 PHY_2901 ();
 sky130_fd_sc_hd__decap_3 PHY_2902 ();
 sky130_fd_sc_hd__decap_3 PHY_2903 ();
 sky130_fd_sc_hd__decap_3 PHY_2904 ();
 sky130_fd_sc_hd__decap_3 PHY_2905 ();
 sky130_fd_sc_hd__decap_3 PHY_2906 ();
 sky130_fd_sc_hd__decap_3 PHY_2907 ();
 sky130_fd_sc_hd__decap_3 PHY_2908 ();
 sky130_fd_sc_hd__decap_3 PHY_2909 ();
 sky130_fd_sc_hd__decap_3 PHY_2910 ();
 sky130_fd_sc_hd__decap_3 PHY_2911 ();
 sky130_fd_sc_hd__decap_3 PHY_2912 ();
 sky130_fd_sc_hd__decap_3 PHY_2913 ();
 sky130_fd_sc_hd__decap_3 PHY_2914 ();
 sky130_fd_sc_hd__decap_3 PHY_2915 ();
 sky130_fd_sc_hd__decap_3 PHY_2916 ();
 sky130_fd_sc_hd__decap_3 PHY_2917 ();
 sky130_fd_sc_hd__decap_3 PHY_2918 ();
 sky130_fd_sc_hd__decap_3 PHY_2919 ();
 sky130_fd_sc_hd__decap_3 PHY_2920 ();
 sky130_fd_sc_hd__decap_3 PHY_2921 ();
 sky130_fd_sc_hd__decap_3 PHY_2922 ();
 sky130_fd_sc_hd__decap_3 PHY_2923 ();
 sky130_fd_sc_hd__decap_3 PHY_2924 ();
 sky130_fd_sc_hd__decap_3 PHY_2925 ();
 sky130_fd_sc_hd__decap_3 PHY_2926 ();
 sky130_fd_sc_hd__decap_3 PHY_2927 ();
 sky130_fd_sc_hd__decap_3 PHY_2928 ();
 sky130_fd_sc_hd__decap_3 PHY_2929 ();
 sky130_fd_sc_hd__decap_3 PHY_2930 ();
 sky130_fd_sc_hd__decap_3 PHY_2931 ();
 sky130_fd_sc_hd__decap_3 PHY_2932 ();
 sky130_fd_sc_hd__decap_3 PHY_2933 ();
 sky130_fd_sc_hd__decap_3 PHY_2934 ();
 sky130_fd_sc_hd__decap_3 PHY_2935 ();
 sky130_fd_sc_hd__decap_3 PHY_2936 ();
 sky130_fd_sc_hd__decap_3 PHY_2937 ();
 sky130_fd_sc_hd__decap_3 PHY_2938 ();
 sky130_fd_sc_hd__decap_3 PHY_2939 ();
 sky130_fd_sc_hd__decap_3 PHY_2940 ();
 sky130_fd_sc_hd__decap_3 PHY_2941 ();
 sky130_fd_sc_hd__decap_3 PHY_2942 ();
 sky130_fd_sc_hd__decap_3 PHY_2943 ();
 sky130_fd_sc_hd__decap_3 PHY_2944 ();
 sky130_fd_sc_hd__decap_3 PHY_2945 ();
 sky130_fd_sc_hd__decap_3 PHY_2946 ();
 sky130_fd_sc_hd__decap_3 PHY_2947 ();
 sky130_fd_sc_hd__decap_3 PHY_2948 ();
 sky130_fd_sc_hd__decap_3 PHY_2949 ();
 sky130_fd_sc_hd__decap_3 PHY_2950 ();
 sky130_fd_sc_hd__decap_3 PHY_2951 ();
 sky130_fd_sc_hd__decap_3 PHY_2952 ();
 sky130_fd_sc_hd__decap_3 PHY_2953 ();
 sky130_fd_sc_hd__decap_3 PHY_2954 ();
 sky130_fd_sc_hd__decap_3 PHY_2955 ();
 sky130_fd_sc_hd__decap_3 PHY_2956 ();
 sky130_fd_sc_hd__decap_3 PHY_2957 ();
 sky130_fd_sc_hd__decap_3 PHY_2958 ();
 sky130_fd_sc_hd__decap_3 PHY_2959 ();
 sky130_fd_sc_hd__decap_3 PHY_2960 ();
 sky130_fd_sc_hd__decap_3 PHY_2961 ();
 sky130_fd_sc_hd__decap_3 PHY_2962 ();
 sky130_fd_sc_hd__decap_3 PHY_2963 ();
 sky130_fd_sc_hd__decap_3 PHY_2964 ();
 sky130_fd_sc_hd__decap_3 PHY_2965 ();
 sky130_fd_sc_hd__decap_3 PHY_2966 ();
 sky130_fd_sc_hd__decap_3 PHY_2967 ();
 sky130_fd_sc_hd__decap_3 PHY_2968 ();
 sky130_fd_sc_hd__decap_3 PHY_2969 ();
 sky130_fd_sc_hd__decap_3 PHY_2970 ();
 sky130_fd_sc_hd__decap_3 PHY_2971 ();
 sky130_fd_sc_hd__decap_3 PHY_2972 ();
 sky130_fd_sc_hd__decap_3 PHY_2973 ();
 sky130_fd_sc_hd__decap_3 PHY_2974 ();
 sky130_fd_sc_hd__decap_3 PHY_2975 ();
 sky130_fd_sc_hd__decap_3 PHY_2976 ();
 sky130_fd_sc_hd__decap_3 PHY_2977 ();
 sky130_fd_sc_hd__decap_3 PHY_2978 ();
 sky130_fd_sc_hd__decap_3 PHY_2979 ();
 sky130_fd_sc_hd__decap_3 PHY_2980 ();
 sky130_fd_sc_hd__decap_3 PHY_2981 ();
 sky130_fd_sc_hd__decap_3 PHY_2982 ();
 sky130_fd_sc_hd__decap_3 PHY_2983 ();
 sky130_fd_sc_hd__decap_3 PHY_2984 ();
 sky130_fd_sc_hd__decap_3 PHY_2985 ();
 sky130_fd_sc_hd__decap_3 PHY_2986 ();
 sky130_fd_sc_hd__decap_3 PHY_2987 ();
 sky130_fd_sc_hd__decap_3 PHY_2988 ();
 sky130_fd_sc_hd__decap_3 PHY_2989 ();
 sky130_fd_sc_hd__decap_3 PHY_2990 ();
 sky130_fd_sc_hd__decap_3 PHY_2991 ();
 sky130_fd_sc_hd__decap_3 PHY_2992 ();
 sky130_fd_sc_hd__decap_3 PHY_2993 ();
 sky130_fd_sc_hd__decap_3 PHY_2994 ();
 sky130_fd_sc_hd__decap_3 PHY_2995 ();
 sky130_fd_sc_hd__decap_3 PHY_2996 ();
 sky130_fd_sc_hd__decap_3 PHY_2997 ();
 sky130_fd_sc_hd__decap_3 PHY_2998 ();
 sky130_fd_sc_hd__decap_3 PHY_2999 ();
 sky130_fd_sc_hd__decap_3 PHY_3000 ();
 sky130_fd_sc_hd__decap_3 PHY_3001 ();
 sky130_fd_sc_hd__decap_3 PHY_3002 ();
 sky130_fd_sc_hd__decap_3 PHY_3003 ();
 sky130_fd_sc_hd__decap_3 PHY_3004 ();
 sky130_fd_sc_hd__decap_3 PHY_3005 ();
 sky130_fd_sc_hd__decap_3 PHY_3006 ();
 sky130_fd_sc_hd__decap_3 PHY_3007 ();
 sky130_fd_sc_hd__decap_3 PHY_3008 ();
 sky130_fd_sc_hd__decap_3 PHY_3009 ();
 sky130_fd_sc_hd__decap_3 PHY_3010 ();
 sky130_fd_sc_hd__decap_3 PHY_3011 ();
 sky130_fd_sc_hd__decap_3 PHY_3012 ();
 sky130_fd_sc_hd__decap_3 PHY_3013 ();
 sky130_fd_sc_hd__decap_3 PHY_3014 ();
 sky130_fd_sc_hd__decap_3 PHY_3015 ();
 sky130_fd_sc_hd__decap_3 PHY_3016 ();
 sky130_fd_sc_hd__decap_3 PHY_3017 ();
 sky130_fd_sc_hd__decap_3 PHY_3018 ();
 sky130_fd_sc_hd__decap_3 PHY_3019 ();
 sky130_fd_sc_hd__decap_3 PHY_3020 ();
 sky130_fd_sc_hd__decap_3 PHY_3021 ();
 sky130_fd_sc_hd__decap_3 PHY_3022 ();
 sky130_fd_sc_hd__decap_3 PHY_3023 ();
 sky130_fd_sc_hd__decap_3 PHY_3024 ();
 sky130_fd_sc_hd__decap_3 PHY_3025 ();
 sky130_fd_sc_hd__decap_3 PHY_3026 ();
 sky130_fd_sc_hd__decap_3 PHY_3027 ();
 sky130_fd_sc_hd__decap_3 PHY_3028 ();
 sky130_fd_sc_hd__decap_3 PHY_3029 ();
 sky130_fd_sc_hd__decap_3 PHY_3030 ();
 sky130_fd_sc_hd__decap_3 PHY_3031 ();
 sky130_fd_sc_hd__decap_3 PHY_3032 ();
 sky130_fd_sc_hd__decap_3 PHY_3033 ();
 sky130_fd_sc_hd__decap_3 PHY_3034 ();
 sky130_fd_sc_hd__decap_3 PHY_3035 ();
 sky130_fd_sc_hd__decap_3 PHY_3036 ();
 sky130_fd_sc_hd__decap_3 PHY_3037 ();
 sky130_fd_sc_hd__decap_3 PHY_3038 ();
 sky130_fd_sc_hd__decap_3 PHY_3039 ();
 sky130_fd_sc_hd__decap_3 PHY_3040 ();
 sky130_fd_sc_hd__decap_3 PHY_3041 ();
 sky130_fd_sc_hd__decap_3 PHY_3042 ();
 sky130_fd_sc_hd__decap_3 PHY_3043 ();
 sky130_fd_sc_hd__decap_3 PHY_3044 ();
 sky130_fd_sc_hd__decap_3 PHY_3045 ();
 sky130_fd_sc_hd__decap_3 PHY_3046 ();
 sky130_fd_sc_hd__decap_3 PHY_3047 ();
 sky130_fd_sc_hd__decap_3 PHY_3048 ();
 sky130_fd_sc_hd__decap_3 PHY_3049 ();
 sky130_fd_sc_hd__decap_3 PHY_3050 ();
 sky130_fd_sc_hd__decap_3 PHY_3051 ();
 sky130_fd_sc_hd__decap_3 PHY_3052 ();
 sky130_fd_sc_hd__decap_3 PHY_3053 ();
 sky130_fd_sc_hd__decap_3 PHY_3054 ();
 sky130_fd_sc_hd__decap_3 PHY_3055 ();
 sky130_fd_sc_hd__decap_3 PHY_3056 ();
 sky130_fd_sc_hd__decap_3 PHY_3057 ();
 sky130_fd_sc_hd__decap_3 PHY_3058 ();
 sky130_fd_sc_hd__decap_3 PHY_3059 ();
 sky130_fd_sc_hd__decap_3 PHY_3060 ();
 sky130_fd_sc_hd__decap_3 PHY_3061 ();
 sky130_fd_sc_hd__decap_3 PHY_3062 ();
 sky130_fd_sc_hd__decap_3 PHY_3063 ();
 sky130_fd_sc_hd__decap_3 PHY_3064 ();
 sky130_fd_sc_hd__decap_3 PHY_3065 ();
 sky130_fd_sc_hd__decap_3 PHY_3066 ();
 sky130_fd_sc_hd__decap_3 PHY_3067 ();
 sky130_fd_sc_hd__decap_3 PHY_3068 ();
 sky130_fd_sc_hd__decap_3 PHY_3069 ();
 sky130_fd_sc_hd__decap_3 PHY_3070 ();
 sky130_fd_sc_hd__decap_3 PHY_3071 ();
 sky130_fd_sc_hd__decap_3 PHY_3072 ();
 sky130_fd_sc_hd__decap_3 PHY_3073 ();
 sky130_fd_sc_hd__decap_3 PHY_3074 ();
 sky130_fd_sc_hd__decap_3 PHY_3075 ();
 sky130_fd_sc_hd__decap_3 PHY_3076 ();
 sky130_fd_sc_hd__decap_3 PHY_3077 ();
 sky130_fd_sc_hd__decap_3 PHY_3078 ();
 sky130_fd_sc_hd__decap_3 PHY_3079 ();
 sky130_fd_sc_hd__decap_3 PHY_3080 ();
 sky130_fd_sc_hd__decap_3 PHY_3081 ();
 sky130_fd_sc_hd__decap_3 PHY_3082 ();
 sky130_fd_sc_hd__decap_3 PHY_3083 ();
 sky130_fd_sc_hd__decap_3 PHY_3084 ();
 sky130_fd_sc_hd__decap_3 PHY_3085 ();
 sky130_fd_sc_hd__decap_3 PHY_3086 ();
 sky130_fd_sc_hd__decap_3 PHY_3087 ();
 sky130_fd_sc_hd__decap_3 PHY_3088 ();
 sky130_fd_sc_hd__decap_3 PHY_3089 ();
 sky130_fd_sc_hd__decap_3 PHY_3090 ();
 sky130_fd_sc_hd__decap_3 PHY_3091 ();
 sky130_fd_sc_hd__decap_3 PHY_3092 ();
 sky130_fd_sc_hd__decap_3 PHY_3093 ();
 sky130_fd_sc_hd__decap_3 PHY_3094 ();
 sky130_fd_sc_hd__decap_3 PHY_3095 ();
 sky130_fd_sc_hd__decap_3 PHY_3096 ();
 sky130_fd_sc_hd__decap_3 PHY_3097 ();
 sky130_fd_sc_hd__decap_3 PHY_3098 ();
 sky130_fd_sc_hd__decap_3 PHY_3099 ();
 sky130_fd_sc_hd__decap_3 PHY_3100 ();
 sky130_fd_sc_hd__decap_3 PHY_3101 ();
 sky130_fd_sc_hd__decap_3 PHY_3102 ();
 sky130_fd_sc_hd__decap_3 PHY_3103 ();
 sky130_fd_sc_hd__decap_3 PHY_3104 ();
 sky130_fd_sc_hd__decap_3 PHY_3105 ();
 sky130_fd_sc_hd__decap_3 PHY_3106 ();
 sky130_fd_sc_hd__decap_3 PHY_3107 ();
 sky130_fd_sc_hd__decap_3 PHY_3108 ();
 sky130_fd_sc_hd__decap_3 PHY_3109 ();
 sky130_fd_sc_hd__decap_3 PHY_3110 ();
 sky130_fd_sc_hd__decap_3 PHY_3111 ();
 sky130_fd_sc_hd__decap_3 PHY_3112 ();
 sky130_fd_sc_hd__decap_3 PHY_3113 ();
 sky130_fd_sc_hd__decap_3 PHY_3114 ();
 sky130_fd_sc_hd__decap_3 PHY_3115 ();
 sky130_fd_sc_hd__decap_3 PHY_3116 ();
 sky130_fd_sc_hd__decap_3 PHY_3117 ();
 sky130_fd_sc_hd__decap_3 PHY_3118 ();
 sky130_fd_sc_hd__decap_3 PHY_3119 ();
 sky130_fd_sc_hd__decap_3 PHY_3120 ();
 sky130_fd_sc_hd__decap_3 PHY_3121 ();
 sky130_fd_sc_hd__decap_3 PHY_3122 ();
 sky130_fd_sc_hd__decap_3 PHY_3123 ();
 sky130_fd_sc_hd__decap_3 PHY_3124 ();
 sky130_fd_sc_hd__decap_3 PHY_3125 ();
 sky130_fd_sc_hd__decap_3 PHY_3126 ();
 sky130_fd_sc_hd__decap_3 PHY_3127 ();
 sky130_fd_sc_hd__decap_3 PHY_3128 ();
 sky130_fd_sc_hd__decap_3 PHY_3129 ();
 sky130_fd_sc_hd__decap_3 PHY_3130 ();
 sky130_fd_sc_hd__decap_3 PHY_3131 ();
 sky130_fd_sc_hd__decap_3 PHY_3132 ();
 sky130_fd_sc_hd__decap_3 PHY_3133 ();
 sky130_fd_sc_hd__decap_3 PHY_3134 ();
 sky130_fd_sc_hd__decap_3 PHY_3135 ();
 sky130_fd_sc_hd__decap_3 PHY_3136 ();
 sky130_fd_sc_hd__decap_3 PHY_3137 ();
 sky130_fd_sc_hd__decap_3 PHY_3138 ();
 sky130_fd_sc_hd__decap_3 PHY_3139 ();
 sky130_fd_sc_hd__decap_3 PHY_3140 ();
 sky130_fd_sc_hd__decap_3 PHY_3141 ();
 sky130_fd_sc_hd__decap_3 PHY_3142 ();
 sky130_fd_sc_hd__decap_3 PHY_3143 ();
 sky130_fd_sc_hd__decap_3 PHY_3144 ();
 sky130_fd_sc_hd__decap_3 PHY_3145 ();
 sky130_fd_sc_hd__decap_3 PHY_3146 ();
 sky130_fd_sc_hd__decap_3 PHY_3147 ();
 sky130_fd_sc_hd__decap_3 PHY_3148 ();
 sky130_fd_sc_hd__decap_3 PHY_3149 ();
 sky130_fd_sc_hd__decap_3 PHY_3150 ();
 sky130_fd_sc_hd__decap_3 PHY_3151 ();
 sky130_fd_sc_hd__decap_3 PHY_3152 ();
 sky130_fd_sc_hd__decap_3 PHY_3153 ();
 sky130_fd_sc_hd__decap_3 PHY_3154 ();
 sky130_fd_sc_hd__decap_3 PHY_3155 ();
 sky130_fd_sc_hd__decap_3 PHY_3156 ();
 sky130_fd_sc_hd__decap_3 PHY_3157 ();
 sky130_fd_sc_hd__decap_3 PHY_3158 ();
 sky130_fd_sc_hd__decap_3 PHY_3159 ();
 sky130_fd_sc_hd__decap_3 PHY_3160 ();
 sky130_fd_sc_hd__decap_3 PHY_3161 ();
 sky130_fd_sc_hd__decap_3 PHY_3162 ();
 sky130_fd_sc_hd__decap_3 PHY_3163 ();
 sky130_fd_sc_hd__decap_3 PHY_3164 ();
 sky130_fd_sc_hd__decap_3 PHY_3165 ();
 sky130_fd_sc_hd__decap_3 PHY_3166 ();
 sky130_fd_sc_hd__decap_3 PHY_3167 ();
 sky130_fd_sc_hd__decap_3 PHY_3168 ();
 sky130_fd_sc_hd__decap_3 PHY_3169 ();
 sky130_fd_sc_hd__decap_3 PHY_3170 ();
 sky130_fd_sc_hd__decap_3 PHY_3171 ();
 sky130_fd_sc_hd__decap_3 PHY_3172 ();
 sky130_fd_sc_hd__decap_3 PHY_3173 ();
 sky130_fd_sc_hd__decap_3 PHY_3174 ();
 sky130_fd_sc_hd__decap_3 PHY_3175 ();
 sky130_fd_sc_hd__decap_3 PHY_3176 ();
 sky130_fd_sc_hd__decap_3 PHY_3177 ();
 sky130_fd_sc_hd__decap_3 PHY_3178 ();
 sky130_fd_sc_hd__decap_3 PHY_3179 ();
 sky130_fd_sc_hd__decap_3 PHY_3180 ();
 sky130_fd_sc_hd__decap_3 PHY_3181 ();
 sky130_fd_sc_hd__decap_3 PHY_3182 ();
 sky130_fd_sc_hd__decap_3 PHY_3183 ();
 sky130_fd_sc_hd__decap_3 PHY_3184 ();
 sky130_fd_sc_hd__decap_3 PHY_3185 ();
 sky130_fd_sc_hd__decap_3 PHY_3186 ();
 sky130_fd_sc_hd__decap_3 PHY_3187 ();
 sky130_fd_sc_hd__decap_3 PHY_3188 ();
 sky130_fd_sc_hd__decap_3 PHY_3189 ();
 sky130_fd_sc_hd__decap_3 PHY_3190 ();
 sky130_fd_sc_hd__decap_3 PHY_3191 ();
 sky130_fd_sc_hd__decap_3 PHY_3192 ();
 sky130_fd_sc_hd__decap_3 PHY_3193 ();
 sky130_fd_sc_hd__decap_3 PHY_3194 ();
 sky130_fd_sc_hd__decap_3 PHY_3195 ();
 sky130_fd_sc_hd__decap_3 PHY_3196 ();
 sky130_fd_sc_hd__decap_3 PHY_3197 ();
 sky130_fd_sc_hd__decap_3 PHY_3198 ();
 sky130_fd_sc_hd__decap_3 PHY_3199 ();
 sky130_fd_sc_hd__decap_3 PHY_3200 ();
 sky130_fd_sc_hd__decap_3 PHY_3201 ();
 sky130_fd_sc_hd__decap_3 PHY_3202 ();
 sky130_fd_sc_hd__decap_3 PHY_3203 ();
 sky130_fd_sc_hd__decap_3 PHY_3204 ();
 sky130_fd_sc_hd__decap_3 PHY_3205 ();
 sky130_fd_sc_hd__decap_3 PHY_3206 ();
 sky130_fd_sc_hd__decap_3 PHY_3207 ();
 sky130_fd_sc_hd__decap_3 PHY_3208 ();
 sky130_fd_sc_hd__decap_3 PHY_3209 ();
 sky130_fd_sc_hd__decap_3 PHY_3210 ();
 sky130_fd_sc_hd__decap_3 PHY_3211 ();
 sky130_fd_sc_hd__decap_3 PHY_3212 ();
 sky130_fd_sc_hd__decap_3 PHY_3213 ();
 sky130_fd_sc_hd__decap_3 PHY_3214 ();
 sky130_fd_sc_hd__decap_3 PHY_3215 ();
 sky130_fd_sc_hd__decap_3 PHY_3216 ();
 sky130_fd_sc_hd__decap_3 PHY_3217 ();
 sky130_fd_sc_hd__decap_3 PHY_3218 ();
 sky130_fd_sc_hd__decap_3 PHY_3219 ();
 sky130_fd_sc_hd__decap_3 PHY_3220 ();
 sky130_fd_sc_hd__decap_3 PHY_3221 ();
 sky130_fd_sc_hd__decap_3 PHY_3222 ();
 sky130_fd_sc_hd__decap_3 PHY_3223 ();
 sky130_fd_sc_hd__decap_3 PHY_3224 ();
 sky130_fd_sc_hd__decap_3 PHY_3225 ();
 sky130_fd_sc_hd__decap_3 PHY_3226 ();
 sky130_fd_sc_hd__decap_3 PHY_3227 ();
 sky130_fd_sc_hd__decap_3 PHY_3228 ();
 sky130_fd_sc_hd__decap_3 PHY_3229 ();
 sky130_fd_sc_hd__decap_3 PHY_3230 ();
 sky130_fd_sc_hd__decap_3 PHY_3231 ();
 sky130_fd_sc_hd__decap_3 PHY_3232 ();
 sky130_fd_sc_hd__decap_3 PHY_3233 ();
 sky130_fd_sc_hd__decap_3 PHY_3234 ();
 sky130_fd_sc_hd__decap_3 PHY_3235 ();
 sky130_fd_sc_hd__decap_3 PHY_3236 ();
 sky130_fd_sc_hd__decap_3 PHY_3237 ();
 sky130_fd_sc_hd__decap_3 PHY_3238 ();
 sky130_fd_sc_hd__decap_3 PHY_3239 ();
 sky130_fd_sc_hd__decap_3 PHY_3240 ();
 sky130_fd_sc_hd__decap_3 PHY_3241 ();
 sky130_fd_sc_hd__decap_3 PHY_3242 ();
 sky130_fd_sc_hd__decap_3 PHY_3243 ();
 sky130_fd_sc_hd__decap_3 PHY_3244 ();
 sky130_fd_sc_hd__decap_3 PHY_3245 ();
 sky130_fd_sc_hd__decap_3 PHY_3246 ();
 sky130_fd_sc_hd__decap_3 PHY_3247 ();
 sky130_fd_sc_hd__decap_3 PHY_3248 ();
 sky130_fd_sc_hd__decap_3 PHY_3249 ();
 sky130_fd_sc_hd__decap_3 PHY_3250 ();
 sky130_fd_sc_hd__decap_3 PHY_3251 ();
 sky130_fd_sc_hd__decap_3 PHY_3252 ();
 sky130_fd_sc_hd__decap_3 PHY_3253 ();
 sky130_fd_sc_hd__decap_3 PHY_3254 ();
 sky130_fd_sc_hd__decap_3 PHY_3255 ();
 sky130_fd_sc_hd__decap_3 PHY_3256 ();
 sky130_fd_sc_hd__decap_3 PHY_3257 ();
 sky130_fd_sc_hd__decap_3 PHY_3258 ();
 sky130_fd_sc_hd__decap_3 PHY_3259 ();
 sky130_fd_sc_hd__decap_3 PHY_3260 ();
 sky130_fd_sc_hd__decap_3 PHY_3261 ();
 sky130_fd_sc_hd__decap_3 PHY_3262 ();
 sky130_fd_sc_hd__decap_3 PHY_3263 ();
 sky130_fd_sc_hd__decap_3 PHY_3264 ();
 sky130_fd_sc_hd__decap_3 PHY_3265 ();
 sky130_fd_sc_hd__decap_3 PHY_3266 ();
 sky130_fd_sc_hd__decap_3 PHY_3267 ();
 sky130_fd_sc_hd__decap_3 PHY_3268 ();
 sky130_fd_sc_hd__decap_3 PHY_3269 ();
 sky130_fd_sc_hd__decap_3 PHY_3270 ();
 sky130_fd_sc_hd__decap_3 PHY_3271 ();
 sky130_fd_sc_hd__decap_3 PHY_3272 ();
 sky130_fd_sc_hd__decap_3 PHY_3273 ();
 sky130_fd_sc_hd__decap_3 PHY_3274 ();
 sky130_fd_sc_hd__decap_3 PHY_3275 ();
 sky130_fd_sc_hd__decap_3 PHY_3276 ();
 sky130_fd_sc_hd__decap_3 PHY_3277 ();
 sky130_fd_sc_hd__decap_3 PHY_3278 ();
 sky130_fd_sc_hd__decap_3 PHY_3279 ();
 sky130_fd_sc_hd__decap_3 PHY_3280 ();
 sky130_fd_sc_hd__decap_3 PHY_3281 ();
 sky130_fd_sc_hd__decap_3 PHY_3282 ();
 sky130_fd_sc_hd__decap_3 PHY_3283 ();
 sky130_fd_sc_hd__decap_3 PHY_3284 ();
 sky130_fd_sc_hd__decap_3 PHY_3285 ();
 sky130_fd_sc_hd__decap_3 PHY_3286 ();
 sky130_fd_sc_hd__decap_3 PHY_3287 ();
 sky130_fd_sc_hd__decap_3 PHY_3288 ();
 sky130_fd_sc_hd__decap_3 PHY_3289 ();
 sky130_fd_sc_hd__decap_3 PHY_3290 ();
 sky130_fd_sc_hd__decap_3 PHY_3291 ();
 sky130_fd_sc_hd__decap_3 PHY_3292 ();
 sky130_fd_sc_hd__decap_3 PHY_3293 ();
 sky130_fd_sc_hd__decap_3 PHY_3294 ();
 sky130_fd_sc_hd__decap_3 PHY_3295 ();
 sky130_fd_sc_hd__decap_3 PHY_3296 ();
 sky130_fd_sc_hd__decap_3 PHY_3297 ();
 sky130_fd_sc_hd__decap_3 PHY_3298 ();
 sky130_fd_sc_hd__decap_3 PHY_3299 ();
 sky130_fd_sc_hd__decap_3 PHY_3300 ();
 sky130_fd_sc_hd__decap_3 PHY_3301 ();
 sky130_fd_sc_hd__decap_3 PHY_3302 ();
 sky130_fd_sc_hd__decap_3 PHY_3303 ();
 sky130_fd_sc_hd__decap_3 PHY_3304 ();
 sky130_fd_sc_hd__decap_3 PHY_3305 ();
 sky130_fd_sc_hd__decap_3 PHY_3306 ();
 sky130_fd_sc_hd__decap_3 PHY_3307 ();
 sky130_fd_sc_hd__decap_3 PHY_3308 ();
 sky130_fd_sc_hd__decap_3 PHY_3309 ();
 sky130_fd_sc_hd__decap_3 PHY_3310 ();
 sky130_fd_sc_hd__decap_3 PHY_3311 ();
 sky130_fd_sc_hd__decap_3 PHY_3312 ();
 sky130_fd_sc_hd__decap_3 PHY_3313 ();
 sky130_fd_sc_hd__decap_3 PHY_3314 ();
 sky130_fd_sc_hd__decap_3 PHY_3315 ();
 sky130_fd_sc_hd__decap_3 PHY_3316 ();
 sky130_fd_sc_hd__decap_3 PHY_3317 ();
 sky130_fd_sc_hd__decap_3 PHY_3318 ();
 sky130_fd_sc_hd__decap_3 PHY_3319 ();
 sky130_fd_sc_hd__decap_3 PHY_3320 ();
 sky130_fd_sc_hd__decap_3 PHY_3321 ();
 sky130_fd_sc_hd__decap_3 PHY_3322 ();
 sky130_fd_sc_hd__decap_3 PHY_3323 ();
 sky130_fd_sc_hd__decap_3 PHY_3324 ();
 sky130_fd_sc_hd__decap_3 PHY_3325 ();
 sky130_fd_sc_hd__decap_3 PHY_3326 ();
 sky130_fd_sc_hd__decap_3 PHY_3327 ();
 sky130_fd_sc_hd__decap_3 PHY_3328 ();
 sky130_fd_sc_hd__decap_3 PHY_3329 ();
 sky130_fd_sc_hd__decap_3 PHY_3330 ();
 sky130_fd_sc_hd__decap_3 PHY_3331 ();
 sky130_fd_sc_hd__decap_3 PHY_3332 ();
 sky130_fd_sc_hd__decap_3 PHY_3333 ();
 sky130_fd_sc_hd__decap_3 PHY_3334 ();
 sky130_fd_sc_hd__decap_3 PHY_3335 ();
 sky130_fd_sc_hd__decap_3 PHY_3336 ();
 sky130_fd_sc_hd__decap_3 PHY_3337 ();
 sky130_fd_sc_hd__decap_3 PHY_3338 ();
 sky130_fd_sc_hd__decap_3 PHY_3339 ();
 sky130_fd_sc_hd__decap_3 PHY_3340 ();
 sky130_fd_sc_hd__decap_3 PHY_3341 ();
 sky130_fd_sc_hd__decap_3 PHY_3342 ();
 sky130_fd_sc_hd__decap_3 PHY_3343 ();
 sky130_fd_sc_hd__decap_3 PHY_3344 ();
 sky130_fd_sc_hd__decap_3 PHY_3345 ();
 sky130_fd_sc_hd__decap_3 PHY_3346 ();
 sky130_fd_sc_hd__decap_3 PHY_3347 ();
 sky130_fd_sc_hd__decap_3 PHY_3348 ();
 sky130_fd_sc_hd__decap_3 PHY_3349 ();
 sky130_fd_sc_hd__decap_3 PHY_3350 ();
 sky130_fd_sc_hd__decap_3 PHY_3351 ();
 sky130_fd_sc_hd__decap_3 PHY_3352 ();
 sky130_fd_sc_hd__decap_3 PHY_3353 ();
 sky130_fd_sc_hd__decap_3 PHY_3354 ();
 sky130_fd_sc_hd__decap_3 PHY_3355 ();
 sky130_fd_sc_hd__decap_3 PHY_3356 ();
 sky130_fd_sc_hd__decap_3 PHY_3357 ();
 sky130_fd_sc_hd__decap_3 PHY_3358 ();
 sky130_fd_sc_hd__decap_3 PHY_3359 ();
 sky130_fd_sc_hd__decap_3 PHY_3360 ();
 sky130_fd_sc_hd__decap_3 PHY_3361 ();
 sky130_fd_sc_hd__decap_3 PHY_3362 ();
 sky130_fd_sc_hd__decap_3 PHY_3363 ();
 sky130_fd_sc_hd__decap_3 PHY_3364 ();
 sky130_fd_sc_hd__decap_3 PHY_3365 ();
 sky130_fd_sc_hd__decap_3 PHY_3366 ();
 sky130_fd_sc_hd__decap_3 PHY_3367 ();
 sky130_fd_sc_hd__decap_3 PHY_3368 ();
 sky130_fd_sc_hd__decap_3 PHY_3369 ();
 sky130_fd_sc_hd__decap_3 PHY_3370 ();
 sky130_fd_sc_hd__decap_3 PHY_3371 ();
 sky130_fd_sc_hd__decap_3 PHY_3372 ();
 sky130_fd_sc_hd__decap_3 PHY_3373 ();
 sky130_fd_sc_hd__decap_3 PHY_3374 ();
 sky130_fd_sc_hd__decap_3 PHY_3375 ();
 sky130_fd_sc_hd__decap_3 PHY_3376 ();
 sky130_fd_sc_hd__decap_3 PHY_3377 ();
 sky130_fd_sc_hd__decap_3 PHY_3378 ();
 sky130_fd_sc_hd__decap_3 PHY_3379 ();
 sky130_fd_sc_hd__decap_3 PHY_3380 ();
 sky130_fd_sc_hd__decap_3 PHY_3381 ();
 sky130_fd_sc_hd__decap_3 PHY_3382 ();
 sky130_fd_sc_hd__decap_3 PHY_3383 ();
 sky130_fd_sc_hd__decap_3 PHY_3384 ();
 sky130_fd_sc_hd__decap_3 PHY_3385 ();
 sky130_fd_sc_hd__decap_3 PHY_3386 ();
 sky130_fd_sc_hd__decap_3 PHY_3387 ();
 sky130_fd_sc_hd__decap_3 PHY_3388 ();
 sky130_fd_sc_hd__decap_3 PHY_3389 ();
 sky130_fd_sc_hd__decap_3 PHY_3390 ();
 sky130_fd_sc_hd__decap_3 PHY_3391 ();
 sky130_fd_sc_hd__decap_3 PHY_3392 ();
 sky130_fd_sc_hd__decap_3 PHY_3393 ();
 sky130_fd_sc_hd__decap_3 PHY_3394 ();
 sky130_fd_sc_hd__decap_3 PHY_3395 ();
 sky130_fd_sc_hd__decap_3 PHY_3396 ();
 sky130_fd_sc_hd__decap_3 PHY_3397 ();
 sky130_fd_sc_hd__decap_3 PHY_3398 ();
 sky130_fd_sc_hd__decap_3 PHY_3399 ();
 sky130_fd_sc_hd__decap_3 PHY_3400 ();
 sky130_fd_sc_hd__decap_3 PHY_3401 ();
 sky130_fd_sc_hd__decap_3 PHY_3402 ();
 sky130_fd_sc_hd__decap_3 PHY_3403 ();
 sky130_fd_sc_hd__decap_3 PHY_3404 ();
 sky130_fd_sc_hd__decap_3 PHY_3405 ();
 sky130_fd_sc_hd__decap_3 PHY_3406 ();
 sky130_fd_sc_hd__decap_3 PHY_3407 ();
 sky130_fd_sc_hd__decap_3 PHY_3408 ();
 sky130_fd_sc_hd__decap_3 PHY_3409 ();
 sky130_fd_sc_hd__decap_3 PHY_3410 ();
 sky130_fd_sc_hd__decap_3 PHY_3411 ();
 sky130_fd_sc_hd__decap_3 PHY_3412 ();
 sky130_fd_sc_hd__decap_3 PHY_3413 ();
 sky130_fd_sc_hd__decap_3 PHY_3414 ();
 sky130_fd_sc_hd__decap_3 PHY_3415 ();
 sky130_fd_sc_hd__decap_3 PHY_3416 ();
 sky130_fd_sc_hd__decap_3 PHY_3417 ();
 sky130_fd_sc_hd__decap_3 PHY_3418 ();
 sky130_fd_sc_hd__decap_3 PHY_3419 ();
 sky130_fd_sc_hd__decap_3 PHY_3420 ();
 sky130_fd_sc_hd__decap_3 PHY_3421 ();
 sky130_fd_sc_hd__decap_3 PHY_3422 ();
 sky130_fd_sc_hd__decap_3 PHY_3423 ();
 sky130_fd_sc_hd__decap_3 PHY_3424 ();
 sky130_fd_sc_hd__decap_3 PHY_3425 ();
 sky130_fd_sc_hd__decap_3 PHY_3426 ();
 sky130_fd_sc_hd__decap_3 PHY_3427 ();
 sky130_fd_sc_hd__decap_3 PHY_3428 ();
 sky130_fd_sc_hd__decap_3 PHY_3429 ();
 sky130_fd_sc_hd__decap_3 PHY_3430 ();
 sky130_fd_sc_hd__decap_3 PHY_3431 ();
 sky130_fd_sc_hd__decap_3 PHY_3432 ();
 sky130_fd_sc_hd__decap_3 PHY_3433 ();
 sky130_fd_sc_hd__decap_3 PHY_3434 ();
 sky130_fd_sc_hd__decap_3 PHY_3435 ();
 sky130_fd_sc_hd__decap_3 PHY_3436 ();
 sky130_fd_sc_hd__decap_3 PHY_3437 ();
 sky130_fd_sc_hd__decap_3 PHY_3438 ();
 sky130_fd_sc_hd__decap_3 PHY_3439 ();
 sky130_fd_sc_hd__decap_3 PHY_3440 ();
 sky130_fd_sc_hd__decap_3 PHY_3441 ();
 sky130_fd_sc_hd__decap_3 PHY_3442 ();
 sky130_fd_sc_hd__decap_3 PHY_3443 ();
 sky130_fd_sc_hd__decap_3 PHY_3444 ();
 sky130_fd_sc_hd__decap_3 PHY_3445 ();
 sky130_fd_sc_hd__decap_3 PHY_3446 ();
 sky130_fd_sc_hd__decap_3 PHY_3447 ();
 sky130_fd_sc_hd__decap_3 PHY_3448 ();
 sky130_fd_sc_hd__decap_3 PHY_3449 ();
 sky130_fd_sc_hd__decap_3 PHY_3450 ();
 sky130_fd_sc_hd__decap_3 PHY_3451 ();
 sky130_fd_sc_hd__decap_3 PHY_3452 ();
 sky130_fd_sc_hd__decap_3 PHY_3453 ();
 sky130_fd_sc_hd__decap_3 PHY_3454 ();
 sky130_fd_sc_hd__decap_3 PHY_3455 ();
 sky130_fd_sc_hd__decap_3 PHY_3456 ();
 sky130_fd_sc_hd__decap_3 PHY_3457 ();
 sky130_fd_sc_hd__decap_3 PHY_3458 ();
 sky130_fd_sc_hd__decap_3 PHY_3459 ();
 sky130_fd_sc_hd__decap_3 PHY_3460 ();
 sky130_fd_sc_hd__decap_3 PHY_3461 ();
 sky130_fd_sc_hd__decap_3 PHY_3462 ();
 sky130_fd_sc_hd__decap_3 PHY_3463 ();
 sky130_fd_sc_hd__decap_3 PHY_3464 ();
 sky130_fd_sc_hd__decap_3 PHY_3465 ();
 sky130_fd_sc_hd__decap_3 PHY_3466 ();
 sky130_fd_sc_hd__decap_3 PHY_3467 ();
 sky130_fd_sc_hd__decap_3 PHY_3468 ();
 sky130_fd_sc_hd__decap_3 PHY_3469 ();
 sky130_fd_sc_hd__decap_3 PHY_3470 ();
 sky130_fd_sc_hd__decap_3 PHY_3471 ();
 sky130_fd_sc_hd__decap_3 PHY_3472 ();
 sky130_fd_sc_hd__decap_3 PHY_3473 ();
 sky130_fd_sc_hd__decap_3 PHY_3474 ();
 sky130_fd_sc_hd__decap_3 PHY_3475 ();
 sky130_fd_sc_hd__decap_3 PHY_3476 ();
 sky130_fd_sc_hd__decap_3 PHY_3477 ();
 sky130_fd_sc_hd__decap_3 PHY_3478 ();
 sky130_fd_sc_hd__decap_3 PHY_3479 ();
 sky130_fd_sc_hd__decap_3 PHY_3480 ();
 sky130_fd_sc_hd__decap_3 PHY_3481 ();
 sky130_fd_sc_hd__decap_3 PHY_3482 ();
 sky130_fd_sc_hd__decap_3 PHY_3483 ();
 sky130_fd_sc_hd__decap_3 PHY_3484 ();
 sky130_fd_sc_hd__decap_3 PHY_3485 ();
 sky130_fd_sc_hd__decap_3 PHY_3486 ();
 sky130_fd_sc_hd__decap_3 PHY_3487 ();
 sky130_fd_sc_hd__decap_3 PHY_3488 ();
 sky130_fd_sc_hd__decap_3 PHY_3489 ();
 sky130_fd_sc_hd__decap_3 PHY_3490 ();
 sky130_fd_sc_hd__decap_3 PHY_3491 ();
 sky130_fd_sc_hd__decap_3 PHY_3492 ();
 sky130_fd_sc_hd__decap_3 PHY_3493 ();
 sky130_fd_sc_hd__decap_3 PHY_3494 ();
 sky130_fd_sc_hd__decap_3 PHY_3495 ();
 sky130_fd_sc_hd__decap_3 PHY_3496 ();
 sky130_fd_sc_hd__decap_3 PHY_3497 ();
 sky130_fd_sc_hd__decap_3 PHY_3498 ();
 sky130_fd_sc_hd__decap_3 PHY_3499 ();
 sky130_fd_sc_hd__decap_3 PHY_3500 ();
 sky130_fd_sc_hd__decap_3 PHY_3501 ();
 sky130_fd_sc_hd__decap_3 PHY_3502 ();
 sky130_fd_sc_hd__decap_3 PHY_3503 ();
 sky130_fd_sc_hd__decap_3 PHY_3504 ();
 sky130_fd_sc_hd__decap_3 PHY_3505 ();
 sky130_fd_sc_hd__decap_3 PHY_3506 ();
 sky130_fd_sc_hd__decap_3 PHY_3507 ();
 sky130_fd_sc_hd__decap_3 PHY_3508 ();
 sky130_fd_sc_hd__decap_3 PHY_3509 ();
 sky130_fd_sc_hd__decap_3 PHY_3510 ();
 sky130_fd_sc_hd__decap_3 PHY_3511 ();
 sky130_fd_sc_hd__decap_3 PHY_3512 ();
 sky130_fd_sc_hd__decap_3 PHY_3513 ();
 sky130_fd_sc_hd__decap_3 PHY_3514 ();
 sky130_fd_sc_hd__decap_3 PHY_3515 ();
 sky130_fd_sc_hd__decap_3 PHY_3516 ();
 sky130_fd_sc_hd__decap_3 PHY_3517 ();
 sky130_fd_sc_hd__decap_3 PHY_3518 ();
 sky130_fd_sc_hd__decap_3 PHY_3519 ();
 sky130_fd_sc_hd__decap_3 PHY_3520 ();
 sky130_fd_sc_hd__decap_3 PHY_3521 ();
 sky130_fd_sc_hd__decap_3 PHY_3522 ();
 sky130_fd_sc_hd__decap_3 PHY_3523 ();
 sky130_fd_sc_hd__decap_3 PHY_3524 ();
 sky130_fd_sc_hd__decap_3 PHY_3525 ();
 sky130_fd_sc_hd__decap_3 PHY_3526 ();
 sky130_fd_sc_hd__decap_3 PHY_3527 ();
 sky130_fd_sc_hd__decap_3 PHY_3528 ();
 sky130_fd_sc_hd__decap_3 PHY_3529 ();
 sky130_fd_sc_hd__decap_3 PHY_3530 ();
 sky130_fd_sc_hd__decap_3 PHY_3531 ();
 sky130_fd_sc_hd__decap_3 PHY_3532 ();
 sky130_fd_sc_hd__decap_3 PHY_3533 ();
 sky130_fd_sc_hd__decap_3 PHY_3534 ();
 sky130_fd_sc_hd__decap_3 PHY_3535 ();
 sky130_fd_sc_hd__decap_3 PHY_3536 ();
 sky130_fd_sc_hd__decap_3 PHY_3537 ();
 sky130_fd_sc_hd__decap_3 PHY_3538 ();
 sky130_fd_sc_hd__decap_3 PHY_3539 ();
 sky130_fd_sc_hd__decap_3 PHY_3540 ();
 sky130_fd_sc_hd__decap_3 PHY_3541 ();
 sky130_fd_sc_hd__decap_3 PHY_3542 ();
 sky130_fd_sc_hd__decap_3 PHY_3543 ();
 sky130_fd_sc_hd__decap_3 PHY_3544 ();
 sky130_fd_sc_hd__decap_3 PHY_3545 ();
 sky130_fd_sc_hd__decap_3 PHY_3546 ();
 sky130_fd_sc_hd__decap_3 PHY_3547 ();
 sky130_fd_sc_hd__decap_3 PHY_3548 ();
 sky130_fd_sc_hd__decap_3 PHY_3549 ();
 sky130_fd_sc_hd__decap_3 PHY_3550 ();
 sky130_fd_sc_hd__decap_3 PHY_3551 ();
 sky130_fd_sc_hd__decap_3 PHY_3552 ();
 sky130_fd_sc_hd__decap_3 PHY_3553 ();
 sky130_fd_sc_hd__decap_3 PHY_3554 ();
 sky130_fd_sc_hd__decap_3 PHY_3555 ();
 sky130_fd_sc_hd__decap_3 PHY_3556 ();
 sky130_fd_sc_hd__decap_3 PHY_3557 ();
 sky130_fd_sc_hd__decap_3 PHY_3558 ();
 sky130_fd_sc_hd__decap_3 PHY_3559 ();
 sky130_fd_sc_hd__decap_3 PHY_3560 ();
 sky130_fd_sc_hd__decap_3 PHY_3561 ();
 sky130_fd_sc_hd__decap_3 PHY_3562 ();
 sky130_fd_sc_hd__decap_3 PHY_3563 ();
 sky130_fd_sc_hd__decap_3 PHY_3564 ();
 sky130_fd_sc_hd__decap_3 PHY_3565 ();
 sky130_fd_sc_hd__decap_3 PHY_3566 ();
 sky130_fd_sc_hd__decap_3 PHY_3567 ();
 sky130_fd_sc_hd__decap_3 PHY_3568 ();
 sky130_fd_sc_hd__decap_3 PHY_3569 ();
 sky130_fd_sc_hd__decap_3 PHY_3570 ();
 sky130_fd_sc_hd__decap_3 PHY_3571 ();
 sky130_fd_sc_hd__decap_3 PHY_3572 ();
 sky130_fd_sc_hd__decap_3 PHY_3573 ();
 sky130_fd_sc_hd__decap_3 PHY_3574 ();
 sky130_fd_sc_hd__decap_3 PHY_3575 ();
 sky130_fd_sc_hd__decap_3 PHY_3576 ();
 sky130_fd_sc_hd__decap_3 PHY_3577 ();
 sky130_fd_sc_hd__decap_3 PHY_3578 ();
 sky130_fd_sc_hd__decap_3 PHY_3579 ();
 sky130_fd_sc_hd__decap_3 PHY_3580 ();
 sky130_fd_sc_hd__decap_3 PHY_3581 ();
 sky130_fd_sc_hd__decap_3 PHY_3582 ();
 sky130_fd_sc_hd__decap_3 PHY_3583 ();
 sky130_fd_sc_hd__decap_3 PHY_3584 ();
 sky130_fd_sc_hd__decap_3 PHY_3585 ();
 sky130_fd_sc_hd__decap_3 PHY_3586 ();
 sky130_fd_sc_hd__decap_3 PHY_3587 ();
 sky130_fd_sc_hd__decap_3 PHY_3588 ();
 sky130_fd_sc_hd__decap_3 PHY_3589 ();
 sky130_fd_sc_hd__decap_3 PHY_3590 ();
 sky130_fd_sc_hd__decap_3 PHY_3591 ();
 sky130_fd_sc_hd__decap_3 PHY_3592 ();
 sky130_fd_sc_hd__decap_3 PHY_3593 ();
 sky130_fd_sc_hd__decap_3 PHY_3594 ();
 sky130_fd_sc_hd__decap_3 PHY_3595 ();
 sky130_fd_sc_hd__decap_3 PHY_3596 ();
 sky130_fd_sc_hd__decap_3 PHY_3597 ();
 sky130_fd_sc_hd__decap_3 PHY_3598 ();
 sky130_fd_sc_hd__decap_3 PHY_3599 ();
 sky130_fd_sc_hd__decap_3 PHY_3600 ();
 sky130_fd_sc_hd__decap_3 PHY_3601 ();
 sky130_fd_sc_hd__decap_3 PHY_3602 ();
 sky130_fd_sc_hd__decap_3 PHY_3603 ();
 sky130_fd_sc_hd__decap_3 PHY_3604 ();
 sky130_fd_sc_hd__decap_3 PHY_3605 ();
 sky130_fd_sc_hd__decap_3 PHY_3606 ();
 sky130_fd_sc_hd__decap_3 PHY_3607 ();
 sky130_fd_sc_hd__decap_3 PHY_3608 ();
 sky130_fd_sc_hd__decap_3 PHY_3609 ();
 sky130_fd_sc_hd__decap_3 PHY_3610 ();
 sky130_fd_sc_hd__decap_3 PHY_3611 ();
 sky130_fd_sc_hd__decap_3 PHY_3612 ();
 sky130_fd_sc_hd__decap_3 PHY_3613 ();
 sky130_fd_sc_hd__decap_3 PHY_3614 ();
 sky130_fd_sc_hd__decap_3 PHY_3615 ();
 sky130_fd_sc_hd__decap_3 PHY_3616 ();
 sky130_fd_sc_hd__decap_3 PHY_3617 ();
 sky130_fd_sc_hd__decap_3 PHY_3618 ();
 sky130_fd_sc_hd__decap_3 PHY_3619 ();
 sky130_fd_sc_hd__decap_3 PHY_3620 ();
 sky130_fd_sc_hd__decap_3 PHY_3621 ();
 sky130_fd_sc_hd__decap_3 PHY_3622 ();
 sky130_fd_sc_hd__decap_3 PHY_3623 ();
 sky130_fd_sc_hd__decap_3 PHY_3624 ();
 sky130_fd_sc_hd__decap_3 PHY_3625 ();
 sky130_fd_sc_hd__decap_3 PHY_3626 ();
 sky130_fd_sc_hd__decap_3 PHY_3627 ();
 sky130_fd_sc_hd__decap_3 PHY_3628 ();
 sky130_fd_sc_hd__decap_3 PHY_3629 ();
 sky130_fd_sc_hd__decap_3 PHY_3630 ();
 sky130_fd_sc_hd__decap_3 PHY_3631 ();
 sky130_fd_sc_hd__decap_3 PHY_3632 ();
 sky130_fd_sc_hd__decap_3 PHY_3633 ();
 sky130_fd_sc_hd__decap_3 PHY_3634 ();
 sky130_fd_sc_hd__decap_3 PHY_3635 ();
 sky130_fd_sc_hd__decap_3 PHY_3636 ();
 sky130_fd_sc_hd__decap_3 PHY_3637 ();
 sky130_fd_sc_hd__decap_3 PHY_3638 ();
 sky130_fd_sc_hd__decap_3 PHY_3639 ();
 sky130_fd_sc_hd__decap_3 PHY_3640 ();
 sky130_fd_sc_hd__decap_3 PHY_3641 ();
 sky130_fd_sc_hd__decap_3 PHY_3642 ();
 sky130_fd_sc_hd__decap_3 PHY_3643 ();
 sky130_fd_sc_hd__decap_3 PHY_3644 ();
 sky130_fd_sc_hd__decap_3 PHY_3645 ();
 sky130_fd_sc_hd__decap_3 PHY_3646 ();
 sky130_fd_sc_hd__decap_3 PHY_3647 ();
 sky130_fd_sc_hd__decap_3 PHY_3648 ();
 sky130_fd_sc_hd__decap_3 PHY_3649 ();
 sky130_fd_sc_hd__decap_3 PHY_3650 ();
 sky130_fd_sc_hd__decap_3 PHY_3651 ();
 sky130_fd_sc_hd__decap_3 PHY_3652 ();
 sky130_fd_sc_hd__decap_3 PHY_3653 ();
 sky130_fd_sc_hd__decap_3 PHY_3654 ();
 sky130_fd_sc_hd__decap_3 PHY_3655 ();
 sky130_fd_sc_hd__decap_3 PHY_3656 ();
 sky130_fd_sc_hd__decap_3 PHY_3657 ();
 sky130_fd_sc_hd__decap_3 PHY_3658 ();
 sky130_fd_sc_hd__decap_3 PHY_3659 ();
 sky130_fd_sc_hd__decap_3 PHY_3660 ();
 sky130_fd_sc_hd__decap_3 PHY_3661 ();
 sky130_fd_sc_hd__decap_3 PHY_3662 ();
 sky130_fd_sc_hd__decap_3 PHY_3663 ();
 sky130_fd_sc_hd__decap_3 PHY_3664 ();
 sky130_fd_sc_hd__decap_3 PHY_3665 ();
 sky130_fd_sc_hd__decap_3 PHY_3666 ();
 sky130_fd_sc_hd__decap_3 PHY_3667 ();
 sky130_fd_sc_hd__decap_3 PHY_3668 ();
 sky130_fd_sc_hd__decap_3 PHY_3669 ();
 sky130_fd_sc_hd__decap_3 PHY_3670 ();
 sky130_fd_sc_hd__decap_3 PHY_3671 ();
 sky130_fd_sc_hd__decap_3 PHY_3672 ();
 sky130_fd_sc_hd__decap_3 PHY_3673 ();
 sky130_fd_sc_hd__decap_3 PHY_3674 ();
 sky130_fd_sc_hd__decap_3 PHY_3675 ();
 sky130_fd_sc_hd__decap_3 PHY_3676 ();
 sky130_fd_sc_hd__decap_3 PHY_3677 ();
 sky130_fd_sc_hd__decap_3 PHY_3678 ();
 sky130_fd_sc_hd__decap_3 PHY_3679 ();
 sky130_fd_sc_hd__decap_3 PHY_3680 ();
 sky130_fd_sc_hd__decap_3 PHY_3681 ();
 sky130_fd_sc_hd__decap_3 PHY_3682 ();
 sky130_fd_sc_hd__decap_3 PHY_3683 ();
 sky130_fd_sc_hd__decap_3 PHY_3684 ();
 sky130_fd_sc_hd__decap_3 PHY_3685 ();
 sky130_fd_sc_hd__decap_3 PHY_3686 ();
 sky130_fd_sc_hd__decap_3 PHY_3687 ();
 sky130_fd_sc_hd__decap_3 PHY_3688 ();
 sky130_fd_sc_hd__decap_3 PHY_3689 ();
 sky130_fd_sc_hd__decap_3 PHY_3690 ();
 sky130_fd_sc_hd__decap_3 PHY_3691 ();
 sky130_fd_sc_hd__decap_3 PHY_3692 ();
 sky130_fd_sc_hd__decap_3 PHY_3693 ();
 sky130_fd_sc_hd__decap_3 PHY_3694 ();
 sky130_fd_sc_hd__decap_3 PHY_3695 ();
 sky130_fd_sc_hd__decap_3 PHY_3696 ();
 sky130_fd_sc_hd__decap_3 PHY_3697 ();
 sky130_fd_sc_hd__decap_3 PHY_3698 ();
 sky130_fd_sc_hd__decap_3 PHY_3699 ();
 sky130_fd_sc_hd__decap_3 PHY_3700 ();
 sky130_fd_sc_hd__decap_3 PHY_3701 ();
 sky130_fd_sc_hd__decap_3 PHY_3702 ();
 sky130_fd_sc_hd__decap_3 PHY_3703 ();
 sky130_fd_sc_hd__decap_3 PHY_3704 ();
 sky130_fd_sc_hd__decap_3 PHY_3705 ();
 sky130_fd_sc_hd__decap_3 PHY_3706 ();
 sky130_fd_sc_hd__decap_3 PHY_3707 ();
 sky130_fd_sc_hd__decap_3 PHY_3708 ();
 sky130_fd_sc_hd__decap_3 PHY_3709 ();
 sky130_fd_sc_hd__decap_3 PHY_3710 ();
 sky130_fd_sc_hd__decap_3 PHY_3711 ();
 sky130_fd_sc_hd__decap_3 PHY_3712 ();
 sky130_fd_sc_hd__decap_3 PHY_3713 ();
 sky130_fd_sc_hd__decap_3 PHY_3714 ();
 sky130_fd_sc_hd__decap_3 PHY_3715 ();
 sky130_fd_sc_hd__decap_3 PHY_3716 ();
 sky130_fd_sc_hd__decap_3 PHY_3717 ();
 sky130_fd_sc_hd__decap_3 PHY_3718 ();
 sky130_fd_sc_hd__decap_3 PHY_3719 ();
 sky130_fd_sc_hd__decap_3 PHY_3720 ();
 sky130_fd_sc_hd__decap_3 PHY_3721 ();
 sky130_fd_sc_hd__decap_3 PHY_3722 ();
 sky130_fd_sc_hd__decap_3 PHY_3723 ();
 sky130_fd_sc_hd__decap_3 PHY_3724 ();
 sky130_fd_sc_hd__decap_3 PHY_3725 ();
 sky130_fd_sc_hd__decap_3 PHY_3726 ();
 sky130_fd_sc_hd__decap_3 PHY_3727 ();
 sky130_fd_sc_hd__decap_3 PHY_3728 ();
 sky130_fd_sc_hd__decap_3 PHY_3729 ();
 sky130_fd_sc_hd__decap_3 PHY_3730 ();
 sky130_fd_sc_hd__decap_3 PHY_3731 ();
 sky130_fd_sc_hd__decap_3 PHY_3732 ();
 sky130_fd_sc_hd__decap_3 PHY_3733 ();
 sky130_fd_sc_hd__decap_3 PHY_3734 ();
 sky130_fd_sc_hd__decap_3 PHY_3735 ();
 sky130_fd_sc_hd__decap_3 PHY_3736 ();
 sky130_fd_sc_hd__decap_3 PHY_3737 ();
 sky130_fd_sc_hd__decap_3 PHY_3738 ();
 sky130_fd_sc_hd__decap_3 PHY_3739 ();
 sky130_fd_sc_hd__decap_3 PHY_3740 ();
 sky130_fd_sc_hd__decap_3 PHY_3741 ();
 sky130_fd_sc_hd__decap_3 PHY_3742 ();
 sky130_fd_sc_hd__decap_3 PHY_3743 ();
 sky130_fd_sc_hd__decap_3 PHY_3744 ();
 sky130_fd_sc_hd__decap_3 PHY_3745 ();
 sky130_fd_sc_hd__decap_3 PHY_3746 ();
 sky130_fd_sc_hd__decap_3 PHY_3747 ();
 sky130_fd_sc_hd__decap_3 PHY_3748 ();
 sky130_fd_sc_hd__decap_3 PHY_3749 ();
 sky130_fd_sc_hd__decap_3 PHY_3750 ();
 sky130_fd_sc_hd__decap_3 PHY_3751 ();
 sky130_fd_sc_hd__decap_3 PHY_3752 ();
 sky130_fd_sc_hd__decap_3 PHY_3753 ();
 sky130_fd_sc_hd__decap_3 PHY_3754 ();
 sky130_fd_sc_hd__decap_3 PHY_3755 ();
 sky130_fd_sc_hd__decap_3 PHY_3756 ();
 sky130_fd_sc_hd__decap_3 PHY_3757 ();
 sky130_fd_sc_hd__decap_3 PHY_3758 ();
 sky130_fd_sc_hd__decap_3 PHY_3759 ();
 sky130_fd_sc_hd__decap_3 PHY_3760 ();
 sky130_fd_sc_hd__decap_3 PHY_3761 ();
 sky130_fd_sc_hd__decap_3 PHY_3762 ();
 sky130_fd_sc_hd__decap_3 PHY_3763 ();
 sky130_fd_sc_hd__decap_3 PHY_3764 ();
 sky130_fd_sc_hd__decap_3 PHY_3765 ();
 sky130_fd_sc_hd__decap_3 PHY_3766 ();
 sky130_fd_sc_hd__decap_3 PHY_3767 ();
 sky130_fd_sc_hd__decap_3 PHY_3768 ();
 sky130_fd_sc_hd__decap_3 PHY_3769 ();
 sky130_fd_sc_hd__decap_3 PHY_3770 ();
 sky130_fd_sc_hd__decap_3 PHY_3771 ();
 sky130_fd_sc_hd__decap_3 PHY_3772 ();
 sky130_fd_sc_hd__decap_3 PHY_3773 ();
 sky130_fd_sc_hd__decap_3 PHY_3774 ();
 sky130_fd_sc_hd__decap_3 PHY_3775 ();
 sky130_fd_sc_hd__decap_3 PHY_3776 ();
 sky130_fd_sc_hd__decap_3 PHY_3777 ();
 sky130_fd_sc_hd__decap_3 PHY_3778 ();
 sky130_fd_sc_hd__decap_3 PHY_3779 ();
 sky130_fd_sc_hd__decap_3 PHY_3780 ();
 sky130_fd_sc_hd__decap_3 PHY_3781 ();
 sky130_fd_sc_hd__decap_3 PHY_3782 ();
 sky130_fd_sc_hd__decap_3 PHY_3783 ();
 sky130_fd_sc_hd__decap_3 PHY_3784 ();
 sky130_fd_sc_hd__decap_3 PHY_3785 ();
 sky130_fd_sc_hd__decap_3 PHY_3786 ();
 sky130_fd_sc_hd__decap_3 PHY_3787 ();
 sky130_fd_sc_hd__decap_3 PHY_3788 ();
 sky130_fd_sc_hd__decap_3 PHY_3789 ();
 sky130_fd_sc_hd__decap_3 PHY_3790 ();
 sky130_fd_sc_hd__decap_3 PHY_3791 ();
 sky130_fd_sc_hd__decap_3 PHY_3792 ();
 sky130_fd_sc_hd__decap_3 PHY_3793 ();
 sky130_fd_sc_hd__decap_3 PHY_3794 ();
 sky130_fd_sc_hd__decap_3 PHY_3795 ();
 sky130_fd_sc_hd__decap_3 PHY_3796 ();
 sky130_fd_sc_hd__decap_3 PHY_3797 ();
 sky130_fd_sc_hd__decap_3 PHY_3798 ();
 sky130_fd_sc_hd__decap_3 PHY_3799 ();
 sky130_fd_sc_hd__decap_3 PHY_3800 ();
 sky130_fd_sc_hd__decap_3 PHY_3801 ();
 sky130_fd_sc_hd__decap_3 PHY_3802 ();
 sky130_fd_sc_hd__decap_3 PHY_3803 ();
 sky130_fd_sc_hd__decap_3 PHY_3804 ();
 sky130_fd_sc_hd__decap_3 PHY_3805 ();
 sky130_fd_sc_hd__decap_3 PHY_3806 ();
 sky130_fd_sc_hd__decap_3 PHY_3807 ();
 sky130_fd_sc_hd__decap_3 PHY_3808 ();
 sky130_fd_sc_hd__decap_3 PHY_3809 ();
 sky130_fd_sc_hd__decap_3 PHY_3810 ();
 sky130_fd_sc_hd__decap_3 PHY_3811 ();
 sky130_fd_sc_hd__decap_3 PHY_3812 ();
 sky130_fd_sc_hd__decap_3 PHY_3813 ();
 sky130_fd_sc_hd__decap_3 PHY_3814 ();
 sky130_fd_sc_hd__decap_3 PHY_3815 ();
 sky130_fd_sc_hd__decap_3 PHY_3816 ();
 sky130_fd_sc_hd__decap_3 PHY_3817 ();
 sky130_fd_sc_hd__decap_3 PHY_3818 ();
 sky130_fd_sc_hd__decap_3 PHY_3819 ();
 sky130_fd_sc_hd__decap_3 PHY_3820 ();
 sky130_fd_sc_hd__decap_3 PHY_3821 ();
 sky130_fd_sc_hd__decap_3 PHY_3822 ();
 sky130_fd_sc_hd__decap_3 PHY_3823 ();
 sky130_fd_sc_hd__decap_3 PHY_3824 ();
 sky130_fd_sc_hd__decap_3 PHY_3825 ();
 sky130_fd_sc_hd__decap_3 PHY_3826 ();
 sky130_fd_sc_hd__decap_3 PHY_3827 ();
 sky130_fd_sc_hd__decap_3 PHY_3828 ();
 sky130_fd_sc_hd__decap_3 PHY_3829 ();
 sky130_fd_sc_hd__decap_3 PHY_3830 ();
 sky130_fd_sc_hd__decap_3 PHY_3831 ();
 sky130_fd_sc_hd__decap_3 PHY_3832 ();
 sky130_fd_sc_hd__decap_3 PHY_3833 ();
 sky130_fd_sc_hd__decap_3 PHY_3834 ();
 sky130_fd_sc_hd__decap_3 PHY_3835 ();
 sky130_fd_sc_hd__decap_3 PHY_3836 ();
 sky130_fd_sc_hd__decap_3 PHY_3837 ();
 sky130_fd_sc_hd__decap_3 PHY_3838 ();
 sky130_fd_sc_hd__decap_3 PHY_3839 ();
 sky130_fd_sc_hd__decap_3 PHY_3840 ();
 sky130_fd_sc_hd__decap_3 PHY_3841 ();
 sky130_fd_sc_hd__decap_3 PHY_3842 ();
 sky130_fd_sc_hd__decap_3 PHY_3843 ();
 sky130_fd_sc_hd__decap_3 PHY_3844 ();
 sky130_fd_sc_hd__decap_3 PHY_3845 ();
 sky130_fd_sc_hd__decap_3 PHY_3846 ();
 sky130_fd_sc_hd__decap_3 PHY_3847 ();
 sky130_fd_sc_hd__decap_3 PHY_3848 ();
 sky130_fd_sc_hd__decap_3 PHY_3849 ();
 sky130_fd_sc_hd__decap_3 PHY_3850 ();
 sky130_fd_sc_hd__decap_3 PHY_3851 ();
 sky130_fd_sc_hd__decap_3 PHY_3852 ();
 sky130_fd_sc_hd__decap_3 PHY_3853 ();
 sky130_fd_sc_hd__decap_3 PHY_3854 ();
 sky130_fd_sc_hd__decap_3 PHY_3855 ();
 sky130_fd_sc_hd__decap_3 PHY_3856 ();
 sky130_fd_sc_hd__decap_3 PHY_3857 ();
 sky130_fd_sc_hd__decap_3 PHY_3858 ();
 sky130_fd_sc_hd__decap_3 PHY_3859 ();
 sky130_fd_sc_hd__decap_3 PHY_3860 ();
 sky130_fd_sc_hd__decap_3 PHY_3861 ();
 sky130_fd_sc_hd__decap_3 PHY_3862 ();
 sky130_fd_sc_hd__decap_3 PHY_3863 ();
 sky130_fd_sc_hd__decap_3 PHY_3864 ();
 sky130_fd_sc_hd__decap_3 PHY_3865 ();
 sky130_fd_sc_hd__decap_3 PHY_3866 ();
 sky130_fd_sc_hd__decap_3 PHY_3867 ();
 sky130_fd_sc_hd__decap_3 PHY_3868 ();
 sky130_fd_sc_hd__decap_3 PHY_3869 ();
 sky130_fd_sc_hd__decap_3 PHY_3870 ();
 sky130_fd_sc_hd__decap_3 PHY_3871 ();
 sky130_fd_sc_hd__decap_3 PHY_3872 ();
 sky130_fd_sc_hd__decap_3 PHY_3873 ();
 sky130_fd_sc_hd__decap_3 PHY_3874 ();
 sky130_fd_sc_hd__decap_3 PHY_3875 ();
 sky130_fd_sc_hd__decap_3 PHY_3876 ();
 sky130_fd_sc_hd__decap_3 PHY_3877 ();
 sky130_fd_sc_hd__decap_3 PHY_3878 ();
 sky130_fd_sc_hd__decap_3 PHY_3879 ();
 sky130_fd_sc_hd__decap_3 PHY_3880 ();
 sky130_fd_sc_hd__decap_3 PHY_3881 ();
 sky130_fd_sc_hd__decap_3 PHY_3882 ();
 sky130_fd_sc_hd__decap_3 PHY_3883 ();
 sky130_fd_sc_hd__decap_3 PHY_3884 ();
 sky130_fd_sc_hd__decap_3 PHY_3885 ();
 sky130_fd_sc_hd__decap_3 PHY_3886 ();
 sky130_fd_sc_hd__decap_3 PHY_3887 ();
 sky130_fd_sc_hd__decap_3 PHY_3888 ();
 sky130_fd_sc_hd__decap_3 PHY_3889 ();
 sky130_fd_sc_hd__decap_3 PHY_3890 ();
 sky130_fd_sc_hd__decap_3 PHY_3891 ();
 sky130_fd_sc_hd__decap_3 PHY_3892 ();
 sky130_fd_sc_hd__decap_3 PHY_3893 ();
 sky130_fd_sc_hd__decap_3 PHY_3894 ();
 sky130_fd_sc_hd__decap_3 PHY_3895 ();
 sky130_fd_sc_hd__decap_3 PHY_3896 ();
 sky130_fd_sc_hd__decap_3 PHY_3897 ();
 sky130_fd_sc_hd__decap_3 PHY_3898 ();
 sky130_fd_sc_hd__decap_3 PHY_3899 ();
 sky130_fd_sc_hd__decap_3 PHY_3900 ();
 sky130_fd_sc_hd__decap_3 PHY_3901 ();
 sky130_fd_sc_hd__decap_3 PHY_3902 ();
 sky130_fd_sc_hd__decap_3 PHY_3903 ();
 sky130_fd_sc_hd__decap_3 PHY_3904 ();
 sky130_fd_sc_hd__decap_3 PHY_3905 ();
 sky130_fd_sc_hd__decap_3 PHY_3906 ();
 sky130_fd_sc_hd__decap_3 PHY_3907 ();
 sky130_fd_sc_hd__decap_3 PHY_3908 ();
 sky130_fd_sc_hd__decap_3 PHY_3909 ();
 sky130_fd_sc_hd__decap_3 PHY_3910 ();
 sky130_fd_sc_hd__decap_3 PHY_3911 ();
 sky130_fd_sc_hd__decap_3 PHY_3912 ();
 sky130_fd_sc_hd__decap_3 PHY_3913 ();
 sky130_fd_sc_hd__decap_3 PHY_3914 ();
 sky130_fd_sc_hd__decap_3 PHY_3915 ();
 sky130_fd_sc_hd__decap_3 PHY_3916 ();
 sky130_fd_sc_hd__decap_3 PHY_3917 ();
 sky130_fd_sc_hd__decap_3 PHY_3918 ();
 sky130_fd_sc_hd__decap_3 PHY_3919 ();
 sky130_fd_sc_hd__decap_3 PHY_3920 ();
 sky130_fd_sc_hd__decap_3 PHY_3921 ();
 sky130_fd_sc_hd__decap_3 PHY_3922 ();
 sky130_fd_sc_hd__decap_3 PHY_3923 ();
 sky130_fd_sc_hd__decap_3 PHY_3924 ();
 sky130_fd_sc_hd__decap_3 PHY_3925 ();
 sky130_fd_sc_hd__decap_3 PHY_3926 ();
 sky130_fd_sc_hd__decap_3 PHY_3927 ();
 sky130_fd_sc_hd__decap_3 PHY_3928 ();
 sky130_fd_sc_hd__decap_3 PHY_3929 ();
 sky130_fd_sc_hd__decap_3 PHY_3930 ();
 sky130_fd_sc_hd__decap_3 PHY_3931 ();
 sky130_fd_sc_hd__decap_3 PHY_3932 ();
 sky130_fd_sc_hd__decap_3 PHY_3933 ();
 sky130_fd_sc_hd__decap_3 PHY_3934 ();
 sky130_fd_sc_hd__decap_3 PHY_3935 ();
 sky130_fd_sc_hd__decap_3 PHY_3936 ();
 sky130_fd_sc_hd__decap_3 PHY_3937 ();
 sky130_fd_sc_hd__decap_3 PHY_3938 ();
 sky130_fd_sc_hd__decap_3 PHY_3939 ();
 sky130_fd_sc_hd__decap_3 PHY_3940 ();
 sky130_fd_sc_hd__decap_3 PHY_3941 ();
 sky130_fd_sc_hd__decap_3 PHY_3942 ();
 sky130_fd_sc_hd__decap_3 PHY_3943 ();
 sky130_fd_sc_hd__decap_3 PHY_3944 ();
 sky130_fd_sc_hd__decap_3 PHY_3945 ();
 sky130_fd_sc_hd__decap_3 PHY_3946 ();
 sky130_fd_sc_hd__decap_3 PHY_3947 ();
 sky130_fd_sc_hd__decap_3 PHY_3948 ();
 sky130_fd_sc_hd__decap_3 PHY_3949 ();
 sky130_fd_sc_hd__decap_3 PHY_3950 ();
 sky130_fd_sc_hd__decap_3 PHY_3951 ();
 sky130_fd_sc_hd__decap_3 PHY_3952 ();
 sky130_fd_sc_hd__decap_3 PHY_3953 ();
 sky130_fd_sc_hd__decap_3 PHY_3954 ();
 sky130_fd_sc_hd__decap_3 PHY_3955 ();
 sky130_fd_sc_hd__decap_3 PHY_3956 ();
 sky130_fd_sc_hd__decap_3 PHY_3957 ();
 sky130_fd_sc_hd__decap_3 PHY_3958 ();
 sky130_fd_sc_hd__decap_3 PHY_3959 ();
 sky130_fd_sc_hd__decap_3 PHY_3960 ();
 sky130_fd_sc_hd__decap_3 PHY_3961 ();
 sky130_fd_sc_hd__decap_3 PHY_3962 ();
 sky130_fd_sc_hd__decap_3 PHY_3963 ();
 sky130_fd_sc_hd__decap_3 PHY_3964 ();
 sky130_fd_sc_hd__decap_3 PHY_3965 ();
 sky130_fd_sc_hd__decap_3 PHY_3966 ();
 sky130_fd_sc_hd__decap_3 PHY_3967 ();
 sky130_fd_sc_hd__decap_3 PHY_3968 ();
 sky130_fd_sc_hd__decap_3 PHY_3969 ();
 sky130_fd_sc_hd__decap_3 PHY_3970 ();
 sky130_fd_sc_hd__decap_3 PHY_3971 ();
 sky130_fd_sc_hd__decap_3 PHY_3972 ();
 sky130_fd_sc_hd__decap_3 PHY_3973 ();
 sky130_fd_sc_hd__decap_3 PHY_3974 ();
 sky130_fd_sc_hd__decap_3 PHY_3975 ();
 sky130_fd_sc_hd__decap_3 PHY_3976 ();
 sky130_fd_sc_hd__decap_3 PHY_3977 ();
 sky130_fd_sc_hd__decap_3 PHY_3978 ();
 sky130_fd_sc_hd__decap_3 PHY_3979 ();
 sky130_fd_sc_hd__decap_3 PHY_3980 ();
 sky130_fd_sc_hd__decap_3 PHY_3981 ();
 sky130_fd_sc_hd__decap_3 PHY_3982 ();
 sky130_fd_sc_hd__decap_3 PHY_3983 ();
 sky130_fd_sc_hd__decap_3 PHY_3984 ();
 sky130_fd_sc_hd__decap_3 PHY_3985 ();
 sky130_fd_sc_hd__decap_3 PHY_3986 ();
 sky130_fd_sc_hd__decap_3 PHY_3987 ();
 sky130_fd_sc_hd__decap_3 PHY_3988 ();
 sky130_fd_sc_hd__decap_3 PHY_3989 ();
 sky130_fd_sc_hd__decap_3 PHY_3990 ();
 sky130_fd_sc_hd__decap_3 PHY_3991 ();
 sky130_fd_sc_hd__decap_3 PHY_3992 ();
 sky130_fd_sc_hd__decap_3 PHY_3993 ();
 sky130_fd_sc_hd__decap_3 PHY_3994 ();
 sky130_fd_sc_hd__decap_3 PHY_3995 ();
 sky130_fd_sc_hd__decap_3 PHY_3996 ();
 sky130_fd_sc_hd__decap_3 PHY_3997 ();
 sky130_fd_sc_hd__decap_3 PHY_3998 ();
 sky130_fd_sc_hd__decap_3 PHY_3999 ();
 sky130_fd_sc_hd__decap_3 PHY_4000 ();
 sky130_fd_sc_hd__decap_3 PHY_4001 ();
 sky130_fd_sc_hd__decap_3 PHY_4002 ();
 sky130_fd_sc_hd__decap_3 PHY_4003 ();
 sky130_fd_sc_hd__decap_3 PHY_4004 ();
 sky130_fd_sc_hd__decap_3 PHY_4005 ();
 sky130_fd_sc_hd__decap_3 PHY_4006 ();
 sky130_fd_sc_hd__decap_3 PHY_4007 ();
 sky130_fd_sc_hd__decap_3 PHY_4008 ();
 sky130_fd_sc_hd__decap_3 PHY_4009 ();
 sky130_fd_sc_hd__decap_3 PHY_4010 ();
 sky130_fd_sc_hd__decap_3 PHY_4011 ();
 sky130_fd_sc_hd__decap_3 PHY_4012 ();
 sky130_fd_sc_hd__decap_3 PHY_4013 ();
 sky130_fd_sc_hd__decap_3 PHY_4014 ();
 sky130_fd_sc_hd__decap_3 PHY_4015 ();
 sky130_fd_sc_hd__decap_3 PHY_4016 ();
 sky130_fd_sc_hd__decap_3 PHY_4017 ();
 sky130_fd_sc_hd__decap_3 PHY_4018 ();
 sky130_fd_sc_hd__decap_3 PHY_4019 ();
 sky130_fd_sc_hd__decap_3 PHY_4020 ();
 sky130_fd_sc_hd__decap_3 PHY_4021 ();
 sky130_fd_sc_hd__decap_3 PHY_4022 ();
 sky130_fd_sc_hd__decap_3 PHY_4023 ();
 sky130_fd_sc_hd__decap_3 PHY_4024 ();
 sky130_fd_sc_hd__decap_3 PHY_4025 ();
 sky130_fd_sc_hd__decap_3 PHY_4026 ();
 sky130_fd_sc_hd__decap_3 PHY_4027 ();
 sky130_fd_sc_hd__decap_3 PHY_4028 ();
 sky130_fd_sc_hd__decap_3 PHY_4029 ();
 sky130_fd_sc_hd__decap_3 PHY_4030 ();
 sky130_fd_sc_hd__decap_3 PHY_4031 ();
 sky130_fd_sc_hd__decap_3 PHY_4032 ();
 sky130_fd_sc_hd__decap_3 PHY_4033 ();
 sky130_fd_sc_hd__decap_3 PHY_4034 ();
 sky130_fd_sc_hd__decap_3 PHY_4035 ();
 sky130_fd_sc_hd__decap_3 PHY_4036 ();
 sky130_fd_sc_hd__decap_3 PHY_4037 ();
 sky130_fd_sc_hd__decap_3 PHY_4038 ();
 sky130_fd_sc_hd__decap_3 PHY_4039 ();
 sky130_fd_sc_hd__decap_3 PHY_4040 ();
 sky130_fd_sc_hd__decap_3 PHY_4041 ();
 sky130_fd_sc_hd__decap_3 PHY_4042 ();
 sky130_fd_sc_hd__decap_3 PHY_4043 ();
 sky130_fd_sc_hd__decap_3 PHY_4044 ();
 sky130_fd_sc_hd__decap_3 PHY_4045 ();
 sky130_fd_sc_hd__decap_3 PHY_4046 ();
 sky130_fd_sc_hd__decap_3 PHY_4047 ();
 sky130_fd_sc_hd__decap_3 PHY_4048 ();
 sky130_fd_sc_hd__decap_3 PHY_4049 ();
 sky130_fd_sc_hd__decap_3 PHY_4050 ();
 sky130_fd_sc_hd__decap_3 PHY_4051 ();
 sky130_fd_sc_hd__decap_3 PHY_4052 ();
 sky130_fd_sc_hd__decap_3 PHY_4053 ();
 sky130_fd_sc_hd__decap_3 PHY_4054 ();
 sky130_fd_sc_hd__decap_3 PHY_4055 ();
 sky130_fd_sc_hd__decap_3 PHY_4056 ();
 sky130_fd_sc_hd__decap_3 PHY_4057 ();
 sky130_fd_sc_hd__decap_3 PHY_4058 ();
 sky130_fd_sc_hd__decap_3 PHY_4059 ();
 sky130_fd_sc_hd__decap_3 PHY_4060 ();
 sky130_fd_sc_hd__decap_3 PHY_4061 ();
 sky130_fd_sc_hd__decap_3 PHY_4062 ();
 sky130_fd_sc_hd__decap_3 PHY_4063 ();
 sky130_fd_sc_hd__decap_3 PHY_4064 ();
 sky130_fd_sc_hd__decap_3 PHY_4065 ();
 sky130_fd_sc_hd__decap_3 PHY_4066 ();
 sky130_fd_sc_hd__decap_3 PHY_4067 ();
 sky130_fd_sc_hd__decap_3 PHY_4068 ();
 sky130_fd_sc_hd__decap_3 PHY_4069 ();
 sky130_fd_sc_hd__decap_3 PHY_4070 ();
 sky130_fd_sc_hd__decap_3 PHY_4071 ();
 sky130_fd_sc_hd__decap_3 PHY_4072 ();
 sky130_fd_sc_hd__decap_3 PHY_4073 ();
 sky130_fd_sc_hd__decap_3 PHY_4074 ();
 sky130_fd_sc_hd__decap_3 PHY_4075 ();
 sky130_fd_sc_hd__decap_3 PHY_4076 ();
 sky130_fd_sc_hd__decap_3 PHY_4077 ();
 sky130_fd_sc_hd__decap_3 PHY_4078 ();
 sky130_fd_sc_hd__decap_3 PHY_4079 ();
 sky130_fd_sc_hd__decap_3 PHY_4080 ();
 sky130_fd_sc_hd__decap_3 PHY_4081 ();
 sky130_fd_sc_hd__decap_3 PHY_4082 ();
 sky130_fd_sc_hd__decap_3 PHY_4083 ();
 sky130_fd_sc_hd__decap_3 PHY_4084 ();
 sky130_fd_sc_hd__decap_3 PHY_4085 ();
 sky130_fd_sc_hd__decap_3 PHY_4086 ();
 sky130_fd_sc_hd__decap_3 PHY_4087 ();
 sky130_fd_sc_hd__decap_3 PHY_4088 ();
 sky130_fd_sc_hd__decap_3 PHY_4089 ();
 sky130_fd_sc_hd__decap_3 PHY_4090 ();
 sky130_fd_sc_hd__decap_3 PHY_4091 ();
 sky130_fd_sc_hd__decap_3 PHY_4092 ();
 sky130_fd_sc_hd__decap_3 PHY_4093 ();
 sky130_fd_sc_hd__decap_3 PHY_4094 ();
 sky130_fd_sc_hd__decap_3 PHY_4095 ();
 sky130_fd_sc_hd__decap_3 PHY_4096 ();
 sky130_fd_sc_hd__decap_3 PHY_4097 ();
 sky130_fd_sc_hd__decap_3 PHY_4098 ();
 sky130_fd_sc_hd__decap_3 PHY_4099 ();
 sky130_fd_sc_hd__decap_3 PHY_4100 ();
 sky130_fd_sc_hd__decap_3 PHY_4101 ();
 sky130_fd_sc_hd__decap_3 PHY_4102 ();
 sky130_fd_sc_hd__decap_3 PHY_4103 ();
 sky130_fd_sc_hd__decap_3 PHY_4104 ();
 sky130_fd_sc_hd__decap_3 PHY_4105 ();
 sky130_fd_sc_hd__decap_3 PHY_4106 ();
 sky130_fd_sc_hd__decap_3 PHY_4107 ();
 sky130_fd_sc_hd__decap_3 PHY_4108 ();
 sky130_fd_sc_hd__decap_3 PHY_4109 ();
 sky130_fd_sc_hd__decap_3 PHY_4110 ();
 sky130_fd_sc_hd__decap_3 PHY_4111 ();
 sky130_fd_sc_hd__decap_3 PHY_4112 ();
 sky130_fd_sc_hd__decap_3 PHY_4113 ();
 sky130_fd_sc_hd__decap_3 PHY_4114 ();
 sky130_fd_sc_hd__decap_3 PHY_4115 ();
 sky130_fd_sc_hd__decap_3 PHY_4116 ();
 sky130_fd_sc_hd__decap_3 PHY_4117 ();
 sky130_fd_sc_hd__decap_3 PHY_4118 ();
 sky130_fd_sc_hd__decap_3 PHY_4119 ();
 sky130_fd_sc_hd__decap_3 PHY_4120 ();
 sky130_fd_sc_hd__decap_3 PHY_4121 ();
 sky130_fd_sc_hd__decap_3 PHY_4122 ();
 sky130_fd_sc_hd__decap_3 PHY_4123 ();
 sky130_fd_sc_hd__decap_3 PHY_4124 ();
 sky130_fd_sc_hd__decap_3 PHY_4125 ();
 sky130_fd_sc_hd__decap_3 PHY_4126 ();
 sky130_fd_sc_hd__decap_3 PHY_4127 ();
 sky130_fd_sc_hd__decap_3 PHY_4128 ();
 sky130_fd_sc_hd__decap_3 PHY_4129 ();
 sky130_fd_sc_hd__decap_3 PHY_4130 ();
 sky130_fd_sc_hd__decap_3 PHY_4131 ();
 sky130_fd_sc_hd__decap_3 PHY_4132 ();
 sky130_fd_sc_hd__decap_3 PHY_4133 ();
 sky130_fd_sc_hd__decap_3 PHY_4134 ();
 sky130_fd_sc_hd__decap_3 PHY_4135 ();
 sky130_fd_sc_hd__decap_3 PHY_4136 ();
 sky130_fd_sc_hd__decap_3 PHY_4137 ();
 sky130_fd_sc_hd__decap_3 PHY_4138 ();
 sky130_fd_sc_hd__decap_3 PHY_4139 ();
 sky130_fd_sc_hd__decap_3 PHY_4140 ();
 sky130_fd_sc_hd__decap_3 PHY_4141 ();
 sky130_fd_sc_hd__decap_3 PHY_4142 ();
 sky130_fd_sc_hd__decap_3 PHY_4143 ();
 sky130_fd_sc_hd__decap_3 PHY_4144 ();
 sky130_fd_sc_hd__decap_3 PHY_4145 ();
 sky130_fd_sc_hd__decap_3 PHY_4146 ();
 sky130_fd_sc_hd__decap_3 PHY_4147 ();
 sky130_fd_sc_hd__decap_3 PHY_4148 ();
 sky130_fd_sc_hd__decap_3 PHY_4149 ();
 sky130_fd_sc_hd__decap_3 PHY_4150 ();
 sky130_fd_sc_hd__decap_3 PHY_4151 ();
 sky130_fd_sc_hd__decap_3 PHY_4152 ();
 sky130_fd_sc_hd__decap_3 PHY_4153 ();
 sky130_fd_sc_hd__decap_3 PHY_4154 ();
 sky130_fd_sc_hd__decap_3 PHY_4155 ();
 sky130_fd_sc_hd__decap_3 PHY_4156 ();
 sky130_fd_sc_hd__decap_3 PHY_4157 ();
 sky130_fd_sc_hd__decap_3 PHY_4158 ();
 sky130_fd_sc_hd__decap_3 PHY_4159 ();
 sky130_fd_sc_hd__decap_3 PHY_4160 ();
 sky130_fd_sc_hd__decap_3 PHY_4161 ();
 sky130_fd_sc_hd__decap_3 PHY_4162 ();
 sky130_fd_sc_hd__decap_3 PHY_4163 ();
 sky130_fd_sc_hd__decap_3 PHY_4164 ();
 sky130_fd_sc_hd__decap_3 PHY_4165 ();
 sky130_fd_sc_hd__decap_3 PHY_4166 ();
 sky130_fd_sc_hd__decap_3 PHY_4167 ();
 sky130_fd_sc_hd__decap_3 PHY_4168 ();
 sky130_fd_sc_hd__decap_3 PHY_4169 ();
 sky130_fd_sc_hd__decap_3 PHY_4170 ();
 sky130_fd_sc_hd__decap_3 PHY_4171 ();
 sky130_fd_sc_hd__decap_3 PHY_4172 ();
 sky130_fd_sc_hd__decap_3 PHY_4173 ();
 sky130_fd_sc_hd__decap_3 PHY_4174 ();
 sky130_fd_sc_hd__decap_3 PHY_4175 ();
 sky130_fd_sc_hd__decap_3 PHY_4176 ();
 sky130_fd_sc_hd__decap_3 PHY_4177 ();
 sky130_fd_sc_hd__decap_3 PHY_4178 ();
 sky130_fd_sc_hd__decap_3 PHY_4179 ();
 sky130_fd_sc_hd__decap_3 PHY_4180 ();
 sky130_fd_sc_hd__decap_3 PHY_4181 ();
 sky130_fd_sc_hd__decap_3 PHY_4182 ();
 sky130_fd_sc_hd__decap_3 PHY_4183 ();
 sky130_fd_sc_hd__decap_3 PHY_4184 ();
 sky130_fd_sc_hd__decap_3 PHY_4185 ();
 sky130_fd_sc_hd__decap_3 PHY_4186 ();
 sky130_fd_sc_hd__decap_3 PHY_4187 ();
 sky130_fd_sc_hd__decap_3 PHY_4188 ();
 sky130_fd_sc_hd__decap_3 PHY_4189 ();
 sky130_fd_sc_hd__decap_3 PHY_4190 ();
 sky130_fd_sc_hd__decap_3 PHY_4191 ();
 sky130_fd_sc_hd__decap_3 PHY_4192 ();
 sky130_fd_sc_hd__decap_3 PHY_4193 ();
 sky130_fd_sc_hd__decap_3 PHY_4194 ();
 sky130_fd_sc_hd__decap_3 PHY_4195 ();
 sky130_fd_sc_hd__decap_3 PHY_4196 ();
 sky130_fd_sc_hd__decap_3 PHY_4197 ();
 sky130_fd_sc_hd__decap_3 PHY_4198 ();
 sky130_fd_sc_hd__decap_3 PHY_4199 ();
 sky130_fd_sc_hd__decap_3 PHY_4200 ();
 sky130_fd_sc_hd__decap_3 PHY_4201 ();
 sky130_fd_sc_hd__decap_3 PHY_4202 ();
 sky130_fd_sc_hd__decap_3 PHY_4203 ();
 sky130_fd_sc_hd__decap_3 PHY_4204 ();
 sky130_fd_sc_hd__decap_3 PHY_4205 ();
 sky130_fd_sc_hd__decap_3 PHY_4206 ();
 sky130_fd_sc_hd__decap_3 PHY_4207 ();
 sky130_fd_sc_hd__decap_3 PHY_4208 ();
 sky130_fd_sc_hd__decap_3 PHY_4209 ();
 sky130_fd_sc_hd__decap_3 PHY_4210 ();
 sky130_fd_sc_hd__decap_3 PHY_4211 ();
 sky130_fd_sc_hd__decap_3 PHY_4212 ();
 sky130_fd_sc_hd__decap_3 PHY_4213 ();
 sky130_fd_sc_hd__decap_3 PHY_4214 ();
 sky130_fd_sc_hd__decap_3 PHY_4215 ();
 sky130_fd_sc_hd__decap_3 PHY_4216 ();
 sky130_fd_sc_hd__decap_3 PHY_4217 ();
 sky130_fd_sc_hd__decap_3 PHY_4218 ();
 sky130_fd_sc_hd__decap_3 PHY_4219 ();
 sky130_fd_sc_hd__decap_3 PHY_4220 ();
 sky130_fd_sc_hd__decap_3 PHY_4221 ();
 sky130_fd_sc_hd__decap_3 PHY_4222 ();
 sky130_fd_sc_hd__decap_3 PHY_4223 ();
 sky130_fd_sc_hd__decap_3 PHY_4224 ();
 sky130_fd_sc_hd__decap_3 PHY_4225 ();
 sky130_fd_sc_hd__decap_3 PHY_4226 ();
 sky130_fd_sc_hd__decap_3 PHY_4227 ();
 sky130_fd_sc_hd__decap_3 PHY_4228 ();
 sky130_fd_sc_hd__decap_3 PHY_4229 ();
 sky130_fd_sc_hd__decap_3 PHY_4230 ();
 sky130_fd_sc_hd__decap_3 PHY_4231 ();
 sky130_fd_sc_hd__decap_3 PHY_4232 ();
 sky130_fd_sc_hd__decap_3 PHY_4233 ();
 sky130_fd_sc_hd__decap_3 PHY_4234 ();
 sky130_fd_sc_hd__decap_3 PHY_4235 ();
 sky130_fd_sc_hd__decap_3 PHY_4236 ();
 sky130_fd_sc_hd__decap_3 PHY_4237 ();
 sky130_fd_sc_hd__decap_3 PHY_4238 ();
 sky130_fd_sc_hd__decap_3 PHY_4239 ();
 sky130_fd_sc_hd__decap_3 PHY_4240 ();
 sky130_fd_sc_hd__decap_3 PHY_4241 ();
 sky130_fd_sc_hd__decap_3 PHY_4242 ();
 sky130_fd_sc_hd__decap_3 PHY_4243 ();
 sky130_fd_sc_hd__decap_3 PHY_4244 ();
 sky130_fd_sc_hd__decap_3 PHY_4245 ();
 sky130_fd_sc_hd__decap_3 PHY_4246 ();
 sky130_fd_sc_hd__decap_3 PHY_4247 ();
 sky130_fd_sc_hd__decap_3 PHY_4248 ();
 sky130_fd_sc_hd__decap_3 PHY_4249 ();
 sky130_fd_sc_hd__decap_3 PHY_4250 ();
 sky130_fd_sc_hd__decap_3 PHY_4251 ();
 sky130_fd_sc_hd__decap_3 PHY_4252 ();
 sky130_fd_sc_hd__decap_3 PHY_4253 ();
 sky130_fd_sc_hd__decap_3 PHY_4254 ();
 sky130_fd_sc_hd__decap_3 PHY_4255 ();
 sky130_fd_sc_hd__decap_3 PHY_4256 ();
 sky130_fd_sc_hd__decap_3 PHY_4257 ();
 sky130_fd_sc_hd__decap_3 PHY_4258 ();
 sky130_fd_sc_hd__decap_3 PHY_4259 ();
 sky130_fd_sc_hd__decap_3 PHY_4260 ();
 sky130_fd_sc_hd__decap_3 PHY_4261 ();
 sky130_fd_sc_hd__decap_3 PHY_4262 ();
 sky130_fd_sc_hd__decap_3 PHY_4263 ();
 sky130_fd_sc_hd__decap_3 PHY_4264 ();
 sky130_fd_sc_hd__decap_3 PHY_4265 ();
 sky130_fd_sc_hd__decap_3 PHY_4266 ();
 sky130_fd_sc_hd__decap_3 PHY_4267 ();
 sky130_fd_sc_hd__decap_3 PHY_4268 ();
 sky130_fd_sc_hd__decap_3 PHY_4269 ();
 sky130_fd_sc_hd__decap_3 PHY_4270 ();
 sky130_fd_sc_hd__decap_3 PHY_4271 ();
 sky130_fd_sc_hd__decap_3 PHY_4272 ();
 sky130_fd_sc_hd__decap_3 PHY_4273 ();
 sky130_fd_sc_hd__decap_3 PHY_4274 ();
 sky130_fd_sc_hd__decap_3 PHY_4275 ();
 sky130_fd_sc_hd__decap_3 PHY_4276 ();
 sky130_fd_sc_hd__decap_3 PHY_4277 ();
 sky130_fd_sc_hd__decap_3 PHY_4278 ();
 sky130_fd_sc_hd__decap_3 PHY_4279 ();
 sky130_fd_sc_hd__decap_3 PHY_4280 ();
 sky130_fd_sc_hd__decap_3 PHY_4281 ();
 sky130_fd_sc_hd__decap_3 PHY_4282 ();
 sky130_fd_sc_hd__decap_3 PHY_4283 ();
 sky130_fd_sc_hd__decap_3 PHY_4284 ();
 sky130_fd_sc_hd__decap_3 PHY_4285 ();
 sky130_fd_sc_hd__decap_3 PHY_4286 ();
 sky130_fd_sc_hd__decap_3 PHY_4287 ();
 sky130_fd_sc_hd__decap_3 PHY_4288 ();
 sky130_fd_sc_hd__decap_3 PHY_4289 ();
 sky130_fd_sc_hd__decap_3 PHY_4290 ();
 sky130_fd_sc_hd__decap_3 PHY_4291 ();
 sky130_fd_sc_hd__decap_3 PHY_4292 ();
 sky130_fd_sc_hd__decap_3 PHY_4293 ();
 sky130_fd_sc_hd__decap_3 PHY_4294 ();
 sky130_fd_sc_hd__decap_3 PHY_4295 ();
 sky130_fd_sc_hd__decap_3 PHY_4296 ();
 sky130_fd_sc_hd__decap_3 PHY_4297 ();
 sky130_fd_sc_hd__decap_3 PHY_4298 ();
 sky130_fd_sc_hd__decap_3 PHY_4299 ();
 sky130_fd_sc_hd__decap_3 PHY_4300 ();
 sky130_fd_sc_hd__decap_3 PHY_4301 ();
 sky130_fd_sc_hd__decap_3 PHY_4302 ();
 sky130_fd_sc_hd__decap_3 PHY_4303 ();
 sky130_fd_sc_hd__decap_3 PHY_4304 ();
 sky130_fd_sc_hd__decap_3 PHY_4305 ();
 sky130_fd_sc_hd__decap_3 PHY_4306 ();
 sky130_fd_sc_hd__decap_3 PHY_4307 ();
 sky130_fd_sc_hd__decap_3 PHY_4308 ();
 sky130_fd_sc_hd__decap_3 PHY_4309 ();
 sky130_fd_sc_hd__decap_3 PHY_4310 ();
 sky130_fd_sc_hd__decap_3 PHY_4311 ();
 sky130_fd_sc_hd__decap_3 PHY_4312 ();
 sky130_fd_sc_hd__decap_3 PHY_4313 ();
 sky130_fd_sc_hd__decap_3 PHY_4314 ();
 sky130_fd_sc_hd__decap_3 PHY_4315 ();
 sky130_fd_sc_hd__decap_3 PHY_4316 ();
 sky130_fd_sc_hd__decap_3 PHY_4317 ();
 sky130_fd_sc_hd__decap_3 PHY_4318 ();
 sky130_fd_sc_hd__decap_3 PHY_4319 ();
 sky130_fd_sc_hd__decap_3 PHY_4320 ();
 sky130_fd_sc_hd__decap_3 PHY_4321 ();
 sky130_fd_sc_hd__decap_3 PHY_4322 ();
 sky130_fd_sc_hd__decap_3 PHY_4323 ();
 sky130_fd_sc_hd__decap_3 PHY_4324 ();
 sky130_fd_sc_hd__decap_3 PHY_4325 ();
 sky130_fd_sc_hd__decap_3 PHY_4326 ();
 sky130_fd_sc_hd__decap_3 PHY_4327 ();
 sky130_fd_sc_hd__decap_3 PHY_4328 ();
 sky130_fd_sc_hd__decap_3 PHY_4329 ();
 sky130_fd_sc_hd__decap_3 PHY_4330 ();
 sky130_fd_sc_hd__decap_3 PHY_4331 ();
 sky130_fd_sc_hd__decap_3 PHY_4332 ();
 sky130_fd_sc_hd__decap_3 PHY_4333 ();
 sky130_fd_sc_hd__decap_3 PHY_4334 ();
 sky130_fd_sc_hd__decap_3 PHY_4335 ();
 sky130_fd_sc_hd__decap_3 PHY_4336 ();
 sky130_fd_sc_hd__decap_3 PHY_4337 ();
 sky130_fd_sc_hd__decap_3 PHY_4338 ();
 sky130_fd_sc_hd__decap_3 PHY_4339 ();
 sky130_fd_sc_hd__decap_3 PHY_4340 ();
 sky130_fd_sc_hd__decap_3 PHY_4341 ();
 sky130_fd_sc_hd__decap_3 PHY_4342 ();
 sky130_fd_sc_hd__decap_3 PHY_4343 ();
 sky130_fd_sc_hd__decap_3 PHY_4344 ();
 sky130_fd_sc_hd__decap_3 PHY_4345 ();
 sky130_fd_sc_hd__decap_3 PHY_4346 ();
 sky130_fd_sc_hd__decap_3 PHY_4347 ();
 sky130_fd_sc_hd__decap_3 PHY_4348 ();
 sky130_fd_sc_hd__decap_3 PHY_4349 ();
 sky130_fd_sc_hd__decap_3 PHY_4350 ();
 sky130_fd_sc_hd__decap_3 PHY_4351 ();
 sky130_fd_sc_hd__decap_3 PHY_4352 ();
 sky130_fd_sc_hd__decap_3 PHY_4353 ();
 sky130_fd_sc_hd__decap_3 PHY_4354 ();
 sky130_fd_sc_hd__decap_3 PHY_4355 ();
 sky130_fd_sc_hd__decap_3 PHY_4356 ();
 sky130_fd_sc_hd__decap_3 PHY_4357 ();
 sky130_fd_sc_hd__decap_3 PHY_4358 ();
 sky130_fd_sc_hd__decap_3 PHY_4359 ();
 sky130_fd_sc_hd__decap_3 PHY_4360 ();
 sky130_fd_sc_hd__decap_3 PHY_4361 ();
 sky130_fd_sc_hd__decap_3 PHY_4362 ();
 sky130_fd_sc_hd__decap_3 PHY_4363 ();
 sky130_fd_sc_hd__decap_3 PHY_4364 ();
 sky130_fd_sc_hd__decap_3 PHY_4365 ();
 sky130_fd_sc_hd__decap_3 PHY_4366 ();
 sky130_fd_sc_hd__decap_3 PHY_4367 ();
 sky130_fd_sc_hd__decap_3 PHY_4368 ();
 sky130_fd_sc_hd__decap_3 PHY_4369 ();
 sky130_fd_sc_hd__decap_3 PHY_4370 ();
 sky130_fd_sc_hd__decap_3 PHY_4371 ();
 sky130_fd_sc_hd__decap_3 PHY_4372 ();
 sky130_fd_sc_hd__decap_3 PHY_4373 ();
 sky130_fd_sc_hd__decap_3 PHY_4374 ();
 sky130_fd_sc_hd__decap_3 PHY_4375 ();
 sky130_fd_sc_hd__decap_3 PHY_4376 ();
 sky130_fd_sc_hd__decap_3 PHY_4377 ();
 sky130_fd_sc_hd__decap_3 PHY_4378 ();
 sky130_fd_sc_hd__decap_3 PHY_4379 ();
 sky130_fd_sc_hd__decap_3 PHY_4380 ();
 sky130_fd_sc_hd__decap_3 PHY_4381 ();
 sky130_fd_sc_hd__decap_3 PHY_4382 ();
 sky130_fd_sc_hd__decap_3 PHY_4383 ();
 sky130_fd_sc_hd__decap_3 PHY_4384 ();
 sky130_fd_sc_hd__decap_3 PHY_4385 ();
 sky130_fd_sc_hd__decap_3 PHY_4386 ();
 sky130_fd_sc_hd__decap_3 PHY_4387 ();
 sky130_fd_sc_hd__decap_3 PHY_4388 ();
 sky130_fd_sc_hd__decap_3 PHY_4389 ();
 sky130_fd_sc_hd__decap_3 PHY_4390 ();
 sky130_fd_sc_hd__decap_3 PHY_4391 ();
 sky130_fd_sc_hd__decap_3 PHY_4392 ();
 sky130_fd_sc_hd__decap_3 PHY_4393 ();
 sky130_fd_sc_hd__decap_3 PHY_4394 ();
 sky130_fd_sc_hd__decap_3 PHY_4395 ();
 sky130_fd_sc_hd__decap_3 PHY_4396 ();
 sky130_fd_sc_hd__decap_3 PHY_4397 ();
 sky130_fd_sc_hd__decap_3 PHY_4398 ();
 sky130_fd_sc_hd__decap_3 PHY_4399 ();
 sky130_fd_sc_hd__decap_3 PHY_4400 ();
 sky130_fd_sc_hd__decap_3 PHY_4401 ();
 sky130_fd_sc_hd__decap_3 PHY_4402 ();
 sky130_fd_sc_hd__decap_3 PHY_4403 ();
 sky130_fd_sc_hd__decap_3 PHY_4404 ();
 sky130_fd_sc_hd__decap_3 PHY_4405 ();
 sky130_fd_sc_hd__decap_3 PHY_4406 ();
 sky130_fd_sc_hd__decap_3 PHY_4407 ();
 sky130_fd_sc_hd__decap_3 PHY_4408 ();
 sky130_fd_sc_hd__decap_3 PHY_4409 ();
 sky130_fd_sc_hd__decap_3 PHY_4410 ();
 sky130_fd_sc_hd__decap_3 PHY_4411 ();
 sky130_fd_sc_hd__decap_3 PHY_4412 ();
 sky130_fd_sc_hd__decap_3 PHY_4413 ();
 sky130_fd_sc_hd__decap_3 PHY_4414 ();
 sky130_fd_sc_hd__decap_3 PHY_4415 ();
 sky130_fd_sc_hd__decap_3 PHY_4416 ();
 sky130_fd_sc_hd__decap_3 PHY_4417 ();
 sky130_fd_sc_hd__decap_3 PHY_4418 ();
 sky130_fd_sc_hd__decap_3 PHY_4419 ();
 sky130_fd_sc_hd__decap_3 PHY_4420 ();
 sky130_fd_sc_hd__decap_3 PHY_4421 ();
 sky130_fd_sc_hd__decap_3 PHY_4422 ();
 sky130_fd_sc_hd__decap_3 PHY_4423 ();
 sky130_fd_sc_hd__decap_3 PHY_4424 ();
 sky130_fd_sc_hd__decap_3 PHY_4425 ();
 sky130_fd_sc_hd__decap_3 PHY_4426 ();
 sky130_fd_sc_hd__decap_3 PHY_4427 ();
 sky130_fd_sc_hd__decap_3 PHY_4428 ();
 sky130_fd_sc_hd__decap_3 PHY_4429 ();
 sky130_fd_sc_hd__decap_3 PHY_4430 ();
 sky130_fd_sc_hd__decap_3 PHY_4431 ();
 sky130_fd_sc_hd__decap_3 PHY_4432 ();
 sky130_fd_sc_hd__decap_3 PHY_4433 ();
 sky130_fd_sc_hd__decap_3 PHY_4434 ();
 sky130_fd_sc_hd__decap_3 PHY_4435 ();
 sky130_fd_sc_hd__decap_3 PHY_4436 ();
 sky130_fd_sc_hd__decap_3 PHY_4437 ();
 sky130_fd_sc_hd__decap_3 PHY_4438 ();
 sky130_fd_sc_hd__decap_3 PHY_4439 ();
 sky130_fd_sc_hd__decap_3 PHY_4440 ();
 sky130_fd_sc_hd__decap_3 PHY_4441 ();
 sky130_fd_sc_hd__decap_3 PHY_4442 ();
 sky130_fd_sc_hd__decap_3 PHY_4443 ();
 sky130_fd_sc_hd__decap_3 PHY_4444 ();
 sky130_fd_sc_hd__decap_3 PHY_4445 ();
 sky130_fd_sc_hd__decap_3 PHY_4446 ();
 sky130_fd_sc_hd__decap_3 PHY_4447 ();
 sky130_fd_sc_hd__decap_3 PHY_4448 ();
 sky130_fd_sc_hd__decap_3 PHY_4449 ();
 sky130_fd_sc_hd__decap_3 PHY_4450 ();
 sky130_fd_sc_hd__decap_3 PHY_4451 ();
 sky130_fd_sc_hd__decap_3 PHY_4452 ();
 sky130_fd_sc_hd__decap_3 PHY_4453 ();
 sky130_fd_sc_hd__decap_3 PHY_4454 ();
 sky130_fd_sc_hd__decap_3 PHY_4455 ();
 sky130_fd_sc_hd__decap_3 PHY_4456 ();
 sky130_fd_sc_hd__decap_3 PHY_4457 ();
 sky130_fd_sc_hd__decap_3 PHY_4458 ();
 sky130_fd_sc_hd__decap_3 PHY_4459 ();
 sky130_fd_sc_hd__decap_3 PHY_4460 ();
 sky130_fd_sc_hd__decap_3 PHY_4461 ();
 sky130_fd_sc_hd__decap_3 PHY_4462 ();
 sky130_fd_sc_hd__decap_3 PHY_4463 ();
 sky130_fd_sc_hd__decap_3 PHY_4464 ();
 sky130_fd_sc_hd__decap_3 PHY_4465 ();
 sky130_fd_sc_hd__decap_3 PHY_4466 ();
 sky130_fd_sc_hd__decap_3 PHY_4467 ();
 sky130_fd_sc_hd__decap_3 PHY_4468 ();
 sky130_fd_sc_hd__decap_3 PHY_4469 ();
 sky130_fd_sc_hd__decap_3 PHY_4470 ();
 sky130_fd_sc_hd__decap_3 PHY_4471 ();
 sky130_fd_sc_hd__decap_3 PHY_4472 ();
 sky130_fd_sc_hd__decap_3 PHY_4473 ();
 sky130_fd_sc_hd__decap_3 PHY_4474 ();
 sky130_fd_sc_hd__decap_3 PHY_4475 ();
 sky130_fd_sc_hd__decap_3 PHY_4476 ();
 sky130_fd_sc_hd__decap_3 PHY_4477 ();
 sky130_fd_sc_hd__decap_3 PHY_4478 ();
 sky130_fd_sc_hd__decap_3 PHY_4479 ();
 sky130_fd_sc_hd__decap_3 PHY_4480 ();
 sky130_fd_sc_hd__decap_3 PHY_4481 ();
 sky130_fd_sc_hd__decap_3 PHY_4482 ();
 sky130_fd_sc_hd__decap_3 PHY_4483 ();
 sky130_fd_sc_hd__decap_3 PHY_4484 ();
 sky130_fd_sc_hd__decap_3 PHY_4485 ();
 sky130_fd_sc_hd__decap_3 PHY_4486 ();
 sky130_fd_sc_hd__decap_3 PHY_4487 ();
 sky130_fd_sc_hd__decap_3 PHY_4488 ();
 sky130_fd_sc_hd__decap_3 PHY_4489 ();
 sky130_fd_sc_hd__decap_3 PHY_4490 ();
 sky130_fd_sc_hd__decap_3 PHY_4491 ();
 sky130_fd_sc_hd__decap_3 PHY_4492 ();
 sky130_fd_sc_hd__decap_3 PHY_4493 ();
 sky130_fd_sc_hd__decap_3 PHY_4494 ();
 sky130_fd_sc_hd__decap_3 PHY_4495 ();
 sky130_fd_sc_hd__decap_3 PHY_4496 ();
 sky130_fd_sc_hd__decap_3 PHY_4497 ();
 sky130_fd_sc_hd__decap_3 PHY_4498 ();
 sky130_fd_sc_hd__decap_3 PHY_4499 ();
 sky130_fd_sc_hd__decap_3 PHY_4500 ();
 sky130_fd_sc_hd__decap_3 PHY_4501 ();
 sky130_fd_sc_hd__decap_3 PHY_4502 ();
 sky130_fd_sc_hd__decap_3 PHY_4503 ();
 sky130_fd_sc_hd__decap_3 PHY_4504 ();
 sky130_fd_sc_hd__decap_3 PHY_4505 ();
 sky130_fd_sc_hd__decap_3 PHY_4506 ();
 sky130_fd_sc_hd__decap_3 PHY_4507 ();
 sky130_fd_sc_hd__decap_3 PHY_4508 ();
 sky130_fd_sc_hd__decap_3 PHY_4509 ();
 sky130_fd_sc_hd__decap_3 PHY_4510 ();
 sky130_fd_sc_hd__decap_3 PHY_4511 ();
 sky130_fd_sc_hd__decap_3 PHY_4512 ();
 sky130_fd_sc_hd__decap_3 PHY_4513 ();
 sky130_fd_sc_hd__decap_3 PHY_4514 ();
 sky130_fd_sc_hd__decap_3 PHY_4515 ();
 sky130_fd_sc_hd__decap_3 PHY_4516 ();
 sky130_fd_sc_hd__decap_3 PHY_4517 ();
 sky130_fd_sc_hd__decap_3 PHY_4518 ();
 sky130_fd_sc_hd__decap_3 PHY_4519 ();
 sky130_fd_sc_hd__decap_3 PHY_4520 ();
 sky130_fd_sc_hd__decap_3 PHY_4521 ();
 sky130_fd_sc_hd__decap_3 PHY_4522 ();
 sky130_fd_sc_hd__decap_3 PHY_4523 ();
 sky130_fd_sc_hd__decap_3 PHY_4524 ();
 sky130_fd_sc_hd__decap_3 PHY_4525 ();
 sky130_fd_sc_hd__decap_3 PHY_4526 ();
 sky130_fd_sc_hd__decap_3 PHY_4527 ();
 sky130_fd_sc_hd__decap_3 PHY_4528 ();
 sky130_fd_sc_hd__decap_3 PHY_4529 ();
 sky130_fd_sc_hd__decap_3 PHY_4530 ();
 sky130_fd_sc_hd__decap_3 PHY_4531 ();
 sky130_fd_sc_hd__decap_3 PHY_4532 ();
 sky130_fd_sc_hd__decap_3 PHY_4533 ();
 sky130_fd_sc_hd__decap_3 PHY_4534 ();
 sky130_fd_sc_hd__decap_3 PHY_4535 ();
 sky130_fd_sc_hd__decap_3 PHY_4536 ();
 sky130_fd_sc_hd__decap_3 PHY_4537 ();
 sky130_fd_sc_hd__decap_3 PHY_4538 ();
 sky130_fd_sc_hd__decap_3 PHY_4539 ();
 sky130_fd_sc_hd__decap_3 PHY_4540 ();
 sky130_fd_sc_hd__decap_3 PHY_4541 ();
 sky130_fd_sc_hd__decap_3 PHY_4542 ();
 sky130_fd_sc_hd__decap_3 PHY_4543 ();
 sky130_fd_sc_hd__decap_3 PHY_4544 ();
 sky130_fd_sc_hd__decap_3 PHY_4545 ();
 sky130_fd_sc_hd__decap_3 PHY_4546 ();
 sky130_fd_sc_hd__decap_3 PHY_4547 ();
 sky130_fd_sc_hd__decap_3 PHY_4548 ();
 sky130_fd_sc_hd__decap_3 PHY_4549 ();
 sky130_fd_sc_hd__decap_3 PHY_4550 ();
 sky130_fd_sc_hd__decap_3 PHY_4551 ();
 sky130_fd_sc_hd__decap_3 PHY_4552 ();
 sky130_fd_sc_hd__decap_3 PHY_4553 ();
 sky130_fd_sc_hd__decap_3 PHY_4554 ();
 sky130_fd_sc_hd__decap_3 PHY_4555 ();
 sky130_fd_sc_hd__decap_3 PHY_4556 ();
 sky130_fd_sc_hd__decap_3 PHY_4557 ();
 sky130_fd_sc_hd__decap_3 PHY_4558 ();
 sky130_fd_sc_hd__decap_3 PHY_4559 ();
 sky130_fd_sc_hd__decap_3 PHY_4560 ();
 sky130_fd_sc_hd__decap_3 PHY_4561 ();
 sky130_fd_sc_hd__decap_3 PHY_4562 ();
 sky130_fd_sc_hd__decap_3 PHY_4563 ();
 sky130_fd_sc_hd__decap_3 PHY_4564 ();
 sky130_fd_sc_hd__decap_3 PHY_4565 ();
 sky130_fd_sc_hd__decap_3 PHY_4566 ();
 sky130_fd_sc_hd__decap_3 PHY_4567 ();
 sky130_fd_sc_hd__decap_3 PHY_4568 ();
 sky130_fd_sc_hd__decap_3 PHY_4569 ();
 sky130_fd_sc_hd__decap_3 PHY_4570 ();
 sky130_fd_sc_hd__decap_3 PHY_4571 ();
 sky130_fd_sc_hd__decap_3 PHY_4572 ();
 sky130_fd_sc_hd__decap_3 PHY_4573 ();
 sky130_fd_sc_hd__decap_3 PHY_4574 ();
 sky130_fd_sc_hd__decap_3 PHY_4575 ();
 sky130_fd_sc_hd__decap_3 PHY_4576 ();
 sky130_fd_sc_hd__decap_3 PHY_4577 ();
 sky130_fd_sc_hd__decap_3 PHY_4578 ();
 sky130_fd_sc_hd__decap_3 PHY_4579 ();
 sky130_fd_sc_hd__decap_3 PHY_4580 ();
 sky130_fd_sc_hd__decap_3 PHY_4581 ();
 sky130_fd_sc_hd__decap_3 PHY_4582 ();
 sky130_fd_sc_hd__decap_3 PHY_4583 ();
 sky130_fd_sc_hd__decap_3 PHY_4584 ();
 sky130_fd_sc_hd__decap_3 PHY_4585 ();
 sky130_fd_sc_hd__decap_3 PHY_4586 ();
 sky130_fd_sc_hd__decap_3 PHY_4587 ();
 sky130_fd_sc_hd__decap_3 PHY_4588 ();
 sky130_fd_sc_hd__decap_3 PHY_4589 ();
 sky130_fd_sc_hd__decap_3 PHY_4590 ();
 sky130_fd_sc_hd__decap_3 PHY_4591 ();
 sky130_fd_sc_hd__decap_3 PHY_4592 ();
 sky130_fd_sc_hd__decap_3 PHY_4593 ();
 sky130_fd_sc_hd__decap_3 PHY_4594 ();
 sky130_fd_sc_hd__decap_3 PHY_4595 ();
 sky130_fd_sc_hd__decap_3 PHY_4596 ();
 sky130_fd_sc_hd__decap_3 PHY_4597 ();
 sky130_fd_sc_hd__decap_3 PHY_4598 ();
 sky130_fd_sc_hd__decap_3 PHY_4599 ();
 sky130_fd_sc_hd__decap_3 PHY_4600 ();
 sky130_fd_sc_hd__decap_3 PHY_4601 ();
 sky130_fd_sc_hd__decap_3 PHY_4602 ();
 sky130_fd_sc_hd__decap_3 PHY_4603 ();
 sky130_fd_sc_hd__decap_3 PHY_4604 ();
 sky130_fd_sc_hd__decap_3 PHY_4605 ();
 sky130_fd_sc_hd__decap_3 PHY_4606 ();
 sky130_fd_sc_hd__decap_3 PHY_4607 ();
 sky130_fd_sc_hd__decap_3 PHY_4608 ();
 sky130_fd_sc_hd__decap_3 PHY_4609 ();
 sky130_fd_sc_hd__decap_3 PHY_4610 ();
 sky130_fd_sc_hd__decap_3 PHY_4611 ();
 sky130_fd_sc_hd__decap_3 PHY_4612 ();
 sky130_fd_sc_hd__decap_3 PHY_4613 ();
 sky130_fd_sc_hd__decap_3 PHY_4614 ();
 sky130_fd_sc_hd__decap_3 PHY_4615 ();
 sky130_fd_sc_hd__decap_3 PHY_4616 ();
 sky130_fd_sc_hd__decap_3 PHY_4617 ();
 sky130_fd_sc_hd__decap_3 PHY_4618 ();
 sky130_fd_sc_hd__decap_3 PHY_4619 ();
 sky130_fd_sc_hd__decap_3 PHY_4620 ();
 sky130_fd_sc_hd__decap_3 PHY_4621 ();
 sky130_fd_sc_hd__decap_3 PHY_4622 ();
 sky130_fd_sc_hd__decap_3 PHY_4623 ();
 sky130_fd_sc_hd__decap_3 PHY_4624 ();
 sky130_fd_sc_hd__decap_3 PHY_4625 ();
 sky130_fd_sc_hd__decap_3 PHY_4626 ();
 sky130_fd_sc_hd__decap_3 PHY_4627 ();
 sky130_fd_sc_hd__decap_3 PHY_4628 ();
 sky130_fd_sc_hd__decap_3 PHY_4629 ();
 sky130_fd_sc_hd__decap_3 PHY_4630 ();
 sky130_fd_sc_hd__decap_3 PHY_4631 ();
 sky130_fd_sc_hd__decap_3 PHY_4632 ();
 sky130_fd_sc_hd__decap_3 PHY_4633 ();
 sky130_fd_sc_hd__decap_3 PHY_4634 ();
 sky130_fd_sc_hd__decap_3 PHY_4635 ();
 sky130_fd_sc_hd__decap_3 PHY_4636 ();
 sky130_fd_sc_hd__decap_3 PHY_4637 ();
 sky130_fd_sc_hd__decap_3 PHY_4638 ();
 sky130_fd_sc_hd__decap_3 PHY_4639 ();
 sky130_fd_sc_hd__decap_3 PHY_4640 ();
 sky130_fd_sc_hd__decap_3 PHY_4641 ();
 sky130_fd_sc_hd__decap_3 PHY_4642 ();
 sky130_fd_sc_hd__decap_3 PHY_4643 ();
 sky130_fd_sc_hd__decap_3 PHY_4644 ();
 sky130_fd_sc_hd__decap_3 PHY_4645 ();
 sky130_fd_sc_hd__decap_3 PHY_4646 ();
 sky130_fd_sc_hd__decap_3 PHY_4647 ();
 sky130_fd_sc_hd__decap_3 PHY_4648 ();
 sky130_fd_sc_hd__decap_3 PHY_4649 ();
 sky130_fd_sc_hd__decap_3 PHY_4650 ();
 sky130_fd_sc_hd__decap_3 PHY_4651 ();
 sky130_fd_sc_hd__decap_3 PHY_4652 ();
 sky130_fd_sc_hd__decap_3 PHY_4653 ();
 sky130_fd_sc_hd__decap_3 PHY_4654 ();
 sky130_fd_sc_hd__decap_3 PHY_4655 ();
 sky130_fd_sc_hd__decap_3 PHY_4656 ();
 sky130_fd_sc_hd__decap_3 PHY_4657 ();
 sky130_fd_sc_hd__decap_3 PHY_4658 ();
 sky130_fd_sc_hd__decap_3 PHY_4659 ();
 sky130_fd_sc_hd__decap_3 PHY_4660 ();
 sky130_fd_sc_hd__decap_3 PHY_4661 ();
 sky130_fd_sc_hd__decap_3 PHY_4662 ();
 sky130_fd_sc_hd__decap_3 PHY_4663 ();
 sky130_fd_sc_hd__decap_3 PHY_4664 ();
 sky130_fd_sc_hd__decap_3 PHY_4665 ();
 sky130_fd_sc_hd__decap_3 PHY_4666 ();
 sky130_fd_sc_hd__decap_3 PHY_4667 ();
 sky130_fd_sc_hd__decap_3 PHY_4668 ();
 sky130_fd_sc_hd__decap_3 PHY_4669 ();
 sky130_fd_sc_hd__decap_3 PHY_4670 ();
 sky130_fd_sc_hd__decap_3 PHY_4671 ();
 sky130_fd_sc_hd__decap_3 PHY_4672 ();
 sky130_fd_sc_hd__decap_3 PHY_4673 ();
 sky130_fd_sc_hd__decap_3 PHY_4674 ();
 sky130_fd_sc_hd__decap_3 PHY_4675 ();
 sky130_fd_sc_hd__decap_3 PHY_4676 ();
 sky130_fd_sc_hd__decap_3 PHY_4677 ();
 sky130_fd_sc_hd__decap_3 PHY_4678 ();
 sky130_fd_sc_hd__decap_3 PHY_4679 ();
 sky130_fd_sc_hd__decap_3 PHY_4680 ();
 sky130_fd_sc_hd__decap_3 PHY_4681 ();
 sky130_fd_sc_hd__decap_3 PHY_4682 ();
 sky130_fd_sc_hd__decap_3 PHY_4683 ();
 sky130_fd_sc_hd__decap_3 PHY_4684 ();
 sky130_fd_sc_hd__decap_3 PHY_4685 ();
 sky130_fd_sc_hd__decap_3 PHY_4686 ();
 sky130_fd_sc_hd__decap_3 PHY_4687 ();
 sky130_fd_sc_hd__decap_3 PHY_4688 ();
 sky130_fd_sc_hd__decap_3 PHY_4689 ();
 sky130_fd_sc_hd__decap_3 PHY_4690 ();
 sky130_fd_sc_hd__decap_3 PHY_4691 ();
 sky130_fd_sc_hd__decap_3 PHY_4692 ();
 sky130_fd_sc_hd__decap_3 PHY_4693 ();
 sky130_fd_sc_hd__decap_3 PHY_4694 ();
 sky130_fd_sc_hd__decap_3 PHY_4695 ();
 sky130_fd_sc_hd__decap_3 PHY_4696 ();
 sky130_fd_sc_hd__decap_3 PHY_4697 ();
 sky130_fd_sc_hd__decap_3 PHY_4698 ();
 sky130_fd_sc_hd__decap_3 PHY_4699 ();
 sky130_fd_sc_hd__decap_3 PHY_4700 ();
 sky130_fd_sc_hd__decap_3 PHY_4701 ();
 sky130_fd_sc_hd__decap_3 PHY_4702 ();
 sky130_fd_sc_hd__decap_3 PHY_4703 ();
 sky130_fd_sc_hd__decap_3 PHY_4704 ();
 sky130_fd_sc_hd__decap_3 PHY_4705 ();
 sky130_fd_sc_hd__decap_3 PHY_4706 ();
 sky130_fd_sc_hd__decap_3 PHY_4707 ();
 sky130_fd_sc_hd__decap_3 PHY_4708 ();
 sky130_fd_sc_hd__decap_3 PHY_4709 ();
 sky130_fd_sc_hd__decap_3 PHY_4710 ();
 sky130_fd_sc_hd__decap_3 PHY_4711 ();
 sky130_fd_sc_hd__decap_3 PHY_4712 ();
 sky130_fd_sc_hd__decap_3 PHY_4713 ();
 sky130_fd_sc_hd__decap_3 PHY_4714 ();
 sky130_fd_sc_hd__decap_3 PHY_4715 ();
 sky130_fd_sc_hd__decap_3 PHY_4716 ();
 sky130_fd_sc_hd__decap_3 PHY_4717 ();
 sky130_fd_sc_hd__decap_3 PHY_4718 ();
 sky130_fd_sc_hd__decap_3 PHY_4719 ();
 sky130_fd_sc_hd__decap_3 PHY_4720 ();
 sky130_fd_sc_hd__decap_3 PHY_4721 ();
 sky130_fd_sc_hd__decap_3 PHY_4722 ();
 sky130_fd_sc_hd__decap_3 PHY_4723 ();
 sky130_fd_sc_hd__decap_3 PHY_4724 ();
 sky130_fd_sc_hd__decap_3 PHY_4725 ();
 sky130_fd_sc_hd__decap_3 PHY_4726 ();
 sky130_fd_sc_hd__decap_3 PHY_4727 ();
 sky130_fd_sc_hd__decap_3 PHY_4728 ();
 sky130_fd_sc_hd__decap_3 PHY_4729 ();
 sky130_fd_sc_hd__decap_3 PHY_4730 ();
 sky130_fd_sc_hd__decap_3 PHY_4731 ();
 sky130_fd_sc_hd__decap_3 PHY_4732 ();
 sky130_fd_sc_hd__decap_3 PHY_4733 ();
 sky130_fd_sc_hd__decap_3 PHY_4734 ();
 sky130_fd_sc_hd__decap_3 PHY_4735 ();
 sky130_fd_sc_hd__decap_3 PHY_4736 ();
 sky130_fd_sc_hd__decap_3 PHY_4737 ();
 sky130_fd_sc_hd__decap_3 PHY_4738 ();
 sky130_fd_sc_hd__decap_3 PHY_4739 ();
 sky130_fd_sc_hd__decap_3 PHY_4740 ();
 sky130_fd_sc_hd__decap_3 PHY_4741 ();
 sky130_fd_sc_hd__decap_3 PHY_4742 ();
 sky130_fd_sc_hd__decap_3 PHY_4743 ();
 sky130_fd_sc_hd__decap_3 PHY_4744 ();
 sky130_fd_sc_hd__decap_3 PHY_4745 ();
 sky130_fd_sc_hd__decap_3 PHY_4746 ();
 sky130_fd_sc_hd__decap_3 PHY_4747 ();
 sky130_fd_sc_hd__decap_3 PHY_4748 ();
 sky130_fd_sc_hd__decap_3 PHY_4749 ();
 sky130_fd_sc_hd__decap_3 PHY_4750 ();
 sky130_fd_sc_hd__decap_3 PHY_4751 ();
 sky130_fd_sc_hd__decap_3 PHY_4752 ();
 sky130_fd_sc_hd__decap_3 PHY_4753 ();
 sky130_fd_sc_hd__decap_3 PHY_4754 ();
 sky130_fd_sc_hd__decap_3 PHY_4755 ();
 sky130_fd_sc_hd__decap_3 PHY_4756 ();
 sky130_fd_sc_hd__decap_3 PHY_4757 ();
 sky130_fd_sc_hd__decap_3 PHY_4758 ();
 sky130_fd_sc_hd__decap_3 PHY_4759 ();
 sky130_fd_sc_hd__decap_3 PHY_4760 ();
 sky130_fd_sc_hd__decap_3 PHY_4761 ();
 sky130_fd_sc_hd__decap_3 PHY_4762 ();
 sky130_fd_sc_hd__decap_3 PHY_4763 ();
 sky130_fd_sc_hd__decap_3 PHY_4764 ();
 sky130_fd_sc_hd__decap_3 PHY_4765 ();
 sky130_fd_sc_hd__decap_3 PHY_4766 ();
 sky130_fd_sc_hd__decap_3 PHY_4767 ();
 sky130_fd_sc_hd__decap_3 PHY_4768 ();
 sky130_fd_sc_hd__decap_3 PHY_4769 ();
 sky130_fd_sc_hd__decap_3 PHY_4770 ();
 sky130_fd_sc_hd__decap_3 PHY_4771 ();
 sky130_fd_sc_hd__decap_3 PHY_4772 ();
 sky130_fd_sc_hd__decap_3 PHY_4773 ();
 sky130_fd_sc_hd__decap_3 PHY_4774 ();
 sky130_fd_sc_hd__decap_3 PHY_4775 ();
 sky130_fd_sc_hd__decap_3 PHY_4776 ();
 sky130_fd_sc_hd__decap_3 PHY_4777 ();
 sky130_fd_sc_hd__decap_3 PHY_4778 ();
 sky130_fd_sc_hd__decap_3 PHY_4779 ();
 sky130_fd_sc_hd__decap_3 PHY_4780 ();
 sky130_fd_sc_hd__decap_3 PHY_4781 ();
 sky130_fd_sc_hd__decap_3 PHY_4782 ();
 sky130_fd_sc_hd__decap_3 PHY_4783 ();
 sky130_fd_sc_hd__decap_3 PHY_4784 ();
 sky130_fd_sc_hd__decap_3 PHY_4785 ();
 sky130_fd_sc_hd__decap_3 PHY_4786 ();
 sky130_fd_sc_hd__decap_3 PHY_4787 ();
 sky130_fd_sc_hd__decap_3 PHY_4788 ();
 sky130_fd_sc_hd__decap_3 PHY_4789 ();
 sky130_fd_sc_hd__decap_3 PHY_4790 ();
 sky130_fd_sc_hd__decap_3 PHY_4791 ();
 sky130_fd_sc_hd__decap_3 PHY_4792 ();
 sky130_fd_sc_hd__decap_3 PHY_4793 ();
 sky130_fd_sc_hd__decap_3 PHY_4794 ();
 sky130_fd_sc_hd__decap_3 PHY_4795 ();
 sky130_fd_sc_hd__decap_3 PHY_4796 ();
 sky130_fd_sc_hd__decap_3 PHY_4797 ();
 sky130_fd_sc_hd__decap_3 PHY_4798 ();
 sky130_fd_sc_hd__decap_3 PHY_4799 ();
 sky130_fd_sc_hd__decap_3 PHY_4800 ();
 sky130_fd_sc_hd__decap_3 PHY_4801 ();
 sky130_fd_sc_hd__decap_3 PHY_4802 ();
 sky130_fd_sc_hd__decap_3 PHY_4803 ();
 sky130_fd_sc_hd__decap_3 PHY_4804 ();
 sky130_fd_sc_hd__decap_3 PHY_4805 ();
 sky130_fd_sc_hd__decap_3 PHY_4806 ();
 sky130_fd_sc_hd__decap_3 PHY_4807 ();
 sky130_fd_sc_hd__decap_3 PHY_4808 ();
 sky130_fd_sc_hd__decap_3 PHY_4809 ();
 sky130_fd_sc_hd__decap_3 PHY_4810 ();
 sky130_fd_sc_hd__decap_3 PHY_4811 ();
 sky130_fd_sc_hd__decap_3 PHY_4812 ();
 sky130_fd_sc_hd__decap_3 PHY_4813 ();
 sky130_fd_sc_hd__decap_3 PHY_4814 ();
 sky130_fd_sc_hd__decap_3 PHY_4815 ();
 sky130_fd_sc_hd__decap_3 PHY_4816 ();
 sky130_fd_sc_hd__decap_3 PHY_4817 ();
 sky130_fd_sc_hd__decap_3 PHY_4818 ();
 sky130_fd_sc_hd__decap_3 PHY_4819 ();
 sky130_fd_sc_hd__decap_3 PHY_4820 ();
 sky130_fd_sc_hd__decap_3 PHY_4821 ();
 sky130_fd_sc_hd__decap_3 PHY_4822 ();
 sky130_fd_sc_hd__decap_3 PHY_4823 ();
 sky130_fd_sc_hd__decap_3 PHY_4824 ();
 sky130_fd_sc_hd__decap_3 PHY_4825 ();
 sky130_fd_sc_hd__decap_3 PHY_4826 ();
 sky130_fd_sc_hd__decap_3 PHY_4827 ();
 sky130_fd_sc_hd__decap_3 PHY_4828 ();
 sky130_fd_sc_hd__decap_3 PHY_4829 ();
 sky130_fd_sc_hd__decap_3 PHY_4830 ();
 sky130_fd_sc_hd__decap_3 PHY_4831 ();
 sky130_fd_sc_hd__decap_3 PHY_4832 ();
 sky130_fd_sc_hd__decap_3 PHY_4833 ();
 sky130_fd_sc_hd__decap_3 PHY_4834 ();
 sky130_fd_sc_hd__decap_3 PHY_4835 ();
 sky130_fd_sc_hd__decap_3 PHY_4836 ();
 sky130_fd_sc_hd__decap_3 PHY_4837 ();
 sky130_fd_sc_hd__decap_3 PHY_4838 ();
 sky130_fd_sc_hd__decap_3 PHY_4839 ();
 sky130_fd_sc_hd__decap_3 PHY_4840 ();
 sky130_fd_sc_hd__decap_3 PHY_4841 ();
 sky130_fd_sc_hd__decap_3 PHY_4842 ();
 sky130_fd_sc_hd__decap_3 PHY_4843 ();
 sky130_fd_sc_hd__decap_3 PHY_4844 ();
 sky130_fd_sc_hd__decap_3 PHY_4845 ();
 sky130_fd_sc_hd__decap_3 PHY_4846 ();
 sky130_fd_sc_hd__decap_3 PHY_4847 ();
 sky130_fd_sc_hd__decap_3 PHY_4848 ();
 sky130_fd_sc_hd__decap_3 PHY_4849 ();
 sky130_fd_sc_hd__decap_3 PHY_4850 ();
 sky130_fd_sc_hd__decap_3 PHY_4851 ();
 sky130_fd_sc_hd__decap_3 PHY_4852 ();
 sky130_fd_sc_hd__decap_3 PHY_4853 ();
 sky130_fd_sc_hd__decap_3 PHY_4854 ();
 sky130_fd_sc_hd__decap_3 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17888 ();
endmodule
