VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 462.820 BY 460.880 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.450 414.855 384.730 418.855 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.030 44.120 395.310 48.120 ;
    END
  END carry_out
  PIN cb_east_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 50.960 413.495 51.560 ;
    END
  END cb_east_in[0]
  PIN cb_east_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 64.560 413.495 65.160 ;
    END
  END cb_east_in[1]
  PIN cb_east_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 78.160 413.495 78.760 ;
    END
  END cb_east_in[2]
  PIN cb_east_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 92.440 413.495 93.040 ;
    END
  END cb_east_in[3]
  PIN cb_east_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 106.040 413.495 106.640 ;
    END
  END cb_east_in[4]
  PIN cb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 120.320 413.495 120.920 ;
    END
  END cb_east_out[0]
  PIN cb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 133.920 413.495 134.520 ;
    END
  END cb_east_out[1]
  PIN cb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 147.520 413.495 148.120 ;
    END
  END cb_east_out[2]
  PIN cb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 161.800 413.495 162.400 ;
    END
  END cb_east_out[3]
  PIN cb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 175.400 413.495 176.000 ;
    END
  END cb_east_out[4]
  PIN cb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 189.680 413.495 190.280 ;
    END
  END cb_east_out[5]
  PIN cb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 203.280 413.495 203.880 ;
    END
  END cb_east_out[6]
  PIN cb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 216.880 413.495 217.480 ;
    END
  END cb_east_out[7]
  PIN cb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 231.160 413.495 231.760 ;
    END
  END cb_east_out[8]
  PIN cb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 409.495 244.760 413.495 245.360 ;
    END
  END cb_east_out[9]
  PIN cb_north_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.090 414.855 55.370 418.855 ;
    END
  END cb_north_in[0]
  PIN cb_north_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.130 414.855 66.410 418.855 ;
    END
  END cb_north_in[1]
  PIN cb_north_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.630 414.855 77.910 418.855 ;
    END
  END cb_north_in[2]
  PIN cb_north_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.130 414.855 89.410 418.855 ;
    END
  END cb_north_in[3]
  PIN cb_north_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.170 414.855 100.450 418.855 ;
    END
  END cb_north_in[4]
  PIN cb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.670 414.855 111.950 418.855 ;
    END
  END cb_north_out[0]
  PIN cb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.170 414.855 123.450 418.855 ;
    END
  END cb_north_out[1]
  PIN cb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.670 414.855 134.950 418.855 ;
    END
  END cb_north_out[2]
  PIN cb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.710 414.855 145.990 418.855 ;
    END
  END cb_north_out[3]
  PIN cb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.210 414.855 157.490 418.855 ;
    END
  END cb_north_out[4]
  PIN cb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.710 414.855 168.990 418.855 ;
    END
  END cb_north_out[5]
  PIN cb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 179.750 414.855 180.030 418.855 ;
    END
  END cb_north_out[6]
  PIN cb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.250 414.855 191.530 418.855 ;
    END
  END cb_north_out[7]
  PIN cb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.750 414.855 203.030 418.855 ;
    END
  END cb_north_out[8]
  PIN cb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.250 414.855 214.530 418.855 ;
    END
  END cb_north_out[9]
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 395.950 414.855 396.230 418.855 ;
    END
  END cen
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.090 44.120 55.370 48.120 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.590 44.120 66.870 48.120 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.550 44.120 78.830 48.120 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.050 44.120 90.330 48.120 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.010 44.120 102.290 48.120 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.510 44.120 113.790 48.120 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.470 44.120 125.750 48.120 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.970 44.120 137.250 48.120 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.930 44.120 149.210 48.120 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.430 44.120 160.710 48.120 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.390 44.120 172.670 48.120 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.890 44.120 184.170 48.120 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.850 44.120 196.130 48.120 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 207.350 44.120 207.630 48.120 ;
    END
  END clb_south_out[3]
  PIN clb_south_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.310 44.120 219.590 48.120 ;
    END
  END clb_south_out[4]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 50.960 53.480 51.560 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 64.560 53.480 65.160 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 78.160 53.480 78.760 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 92.440 53.480 93.040 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 106.040 53.480 106.640 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 120.320 53.480 120.920 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 133.920 53.480 134.520 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 147.520 53.480 148.120 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 161.800 53.480 162.400 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 175.400 53.480 176.000 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 189.680 53.480 190.280 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 203.280 53.480 203.880 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 216.880 53.480 217.480 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 231.160 53.480 231.760 ;
    END
  END clb_west_out[3]
  PIN clb_west_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 244.760 53.480 245.360 ;
    END
  END clb_west_out[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.990 44.120 407.270 48.120 ;
    END
  END clk
  PIN east_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 314.120 413.495 314.720 ;
    END
  END east_double[0]
  PIN east_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 328.400 413.495 329.000 ;
    END
  END east_double[1]
  PIN east_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 342.000 413.495 342.600 ;
    END
  END east_double[2]
  PIN east_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 355.600 413.495 356.200 ;
    END
  END east_double[3]
  PIN east_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 369.880 413.495 370.480 ;
    END
  END east_double[4]
  PIN east_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 383.480 413.495 384.080 ;
    END
  END east_double[5]
  PIN east_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 397.760 413.495 398.360 ;
    END
  END east_double[6]
  PIN east_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 411.360 413.495 411.960 ;
    END
  END east_double[7]
  PIN east_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 259.040 413.495 259.640 ;
    END
  END east_single[0]
  PIN east_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 272.640 413.495 273.240 ;
    END
  END east_single[1]
  PIN east_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 286.240 413.495 286.840 ;
    END
  END east_single[2]
  PIN east_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 409.495 300.520 413.495 301.120 ;
    END
  END east_single[3]
  PIN north_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 270.830 414.855 271.110 418.855 ;
    END
  END north_double[0]
  PIN north_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 282.330 414.855 282.610 418.855 ;
    END
  END north_double[1]
  PIN north_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 293.830 414.855 294.110 418.855 ;
    END
  END north_double[2]
  PIN north_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 304.870 414.855 305.150 418.855 ;
    END
  END north_double[3]
  PIN north_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 316.370 414.855 316.650 418.855 ;
    END
  END north_double[4]
  PIN north_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 327.870 414.855 328.150 418.855 ;
    END
  END north_double[5]
  PIN north_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 338.910 414.855 339.190 418.855 ;
    END
  END north_double[6]
  PIN north_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 350.410 414.855 350.690 418.855 ;
    END
  END north_double[7]
  PIN north_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 225.290 414.855 225.570 418.855 ;
    END
  END north_single[0]
  PIN north_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 236.790 414.855 237.070 418.855 ;
    END
  END north_single[1]
  PIN north_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 248.290 414.855 248.570 418.855 ;
    END
  END north_single[2]
  PIN north_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 259.330 414.855 259.610 418.855 ;
    END
  END north_single[3]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.450 414.855 407.730 418.855 ;
    END
  END rst
  PIN set_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.530 44.120 383.810 48.120 ;
    END
  END set_in_hard
  PIN set_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.410 414.855 373.690 418.855 ;
    END
  END set_out_hard
  PIN shift_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.570 44.120 371.850 48.120 ;
    END
  END shift_in_hard
  PIN shift_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.910 414.855 362.190 418.855 ;
    END
  END shift_out_hard
  PIN south_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 277.730 44.120 278.010 48.120 ;
    END
  END south_double[0]
  PIN south_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 289.690 44.120 289.970 48.120 ;
    END
  END south_double[1]
  PIN south_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 301.190 44.120 301.470 48.120 ;
    END
  END south_double[2]
  PIN south_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 313.150 44.120 313.430 48.120 ;
    END
  END south_double[3]
  PIN south_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 324.650 44.120 324.930 48.120 ;
    END
  END south_double[4]
  PIN south_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 336.610 44.120 336.890 48.120 ;
    END
  END south_double[5]
  PIN south_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 348.110 44.120 348.390 48.120 ;
    END
  END south_double[6]
  PIN south_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 360.070 44.120 360.350 48.120 ;
    END
  END south_double[7]
  PIN south_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 230.810 44.120 231.090 48.120 ;
    END
  END south_single[0]
  PIN south_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 242.770 44.120 243.050 48.120 ;
    END
  END south_single[1]
  PIN south_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 254.270 44.120 254.550 48.120 ;
    END
  END south_single[2]
  PIN south_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 266.230 44.120 266.510 48.120 ;
    END
  END south_single[3]
  PIN west_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 314.120 53.480 314.720 ;
    END
  END west_double[0]
  PIN west_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 328.400 53.480 329.000 ;
    END
  END west_double[1]
  PIN west_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 342.000 53.480 342.600 ;
    END
  END west_double[2]
  PIN west_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 355.600 53.480 356.200 ;
    END
  END west_double[3]
  PIN west_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 369.880 53.480 370.480 ;
    END
  END west_double[4]
  PIN west_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 383.480 53.480 384.080 ;
    END
  END west_double[5]
  PIN west_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 397.760 53.480 398.360 ;
    END
  END west_double[6]
  PIN west_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 411.360 53.480 411.960 ;
    END
  END west_double[7]
  PIN west_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 259.040 53.480 259.640 ;
    END
  END west_single[0]
  PIN west_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 272.640 53.480 273.240 ;
    END
  END west_single[1]
  PIN west_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 286.240 53.480 286.840 ;
    END
  END west_single[2]
  PIN west_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 300.520 53.480 301.120 ;
    END
  END west_single[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 437.820 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 462.820 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 52.365 408.595 405.965 ;
      LAYER met1 ;
        RECT 55.000 50.280 408.670 410.260 ;
      LAYER met2 ;
        RECT 55.650 414.575 65.850 414.855 ;
        RECT 66.690 414.575 77.350 414.855 ;
        RECT 78.190 414.575 88.850 414.855 ;
        RECT 89.690 414.575 99.890 414.855 ;
        RECT 100.730 414.575 111.390 414.855 ;
        RECT 112.230 414.575 122.890 414.855 ;
        RECT 123.730 414.575 134.390 414.855 ;
        RECT 135.230 414.575 145.430 414.855 ;
        RECT 146.270 414.575 156.930 414.855 ;
        RECT 157.770 414.575 168.430 414.855 ;
        RECT 169.270 414.575 179.470 414.855 ;
        RECT 180.310 414.575 190.970 414.855 ;
        RECT 191.810 414.575 202.470 414.855 ;
        RECT 203.310 414.575 213.970 414.855 ;
        RECT 214.810 414.575 225.010 414.855 ;
        RECT 225.850 414.575 236.510 414.855 ;
        RECT 237.350 414.575 248.010 414.855 ;
        RECT 248.850 414.575 259.050 414.855 ;
        RECT 259.890 414.575 270.550 414.855 ;
        RECT 271.390 414.575 282.050 414.855 ;
        RECT 282.890 414.575 293.550 414.855 ;
        RECT 294.390 414.575 304.590 414.855 ;
        RECT 305.430 414.575 316.090 414.855 ;
        RECT 316.930 414.575 327.590 414.855 ;
        RECT 328.430 414.575 338.630 414.855 ;
        RECT 339.470 414.575 350.130 414.855 ;
        RECT 350.970 414.575 361.630 414.855 ;
        RECT 362.470 414.575 373.130 414.855 ;
        RECT 373.970 414.575 384.170 414.855 ;
        RECT 385.010 414.575 395.670 414.855 ;
        RECT 396.510 414.575 407.170 414.855 ;
        RECT 408.010 414.575 409.110 414.855 ;
        RECT 55.100 48.400 409.110 414.575 ;
        RECT 55.650 48.120 66.310 48.400 ;
        RECT 67.150 48.120 78.270 48.400 ;
        RECT 79.110 48.120 89.770 48.400 ;
        RECT 90.610 48.120 101.730 48.400 ;
        RECT 102.570 48.120 113.230 48.400 ;
        RECT 114.070 48.120 125.190 48.400 ;
        RECT 126.030 48.120 136.690 48.400 ;
        RECT 137.530 48.120 148.650 48.400 ;
        RECT 149.490 48.120 160.150 48.400 ;
        RECT 160.990 48.120 172.110 48.400 ;
        RECT 172.950 48.120 183.610 48.400 ;
        RECT 184.450 48.120 195.570 48.400 ;
        RECT 196.410 48.120 207.070 48.400 ;
        RECT 207.910 48.120 219.030 48.400 ;
        RECT 219.870 48.120 230.530 48.400 ;
        RECT 231.370 48.120 242.490 48.400 ;
        RECT 243.330 48.120 253.990 48.400 ;
        RECT 254.830 48.120 265.950 48.400 ;
        RECT 266.790 48.120 277.450 48.400 ;
        RECT 278.290 48.120 289.410 48.400 ;
        RECT 290.250 48.120 300.910 48.400 ;
        RECT 301.750 48.120 312.870 48.400 ;
        RECT 313.710 48.120 324.370 48.400 ;
        RECT 325.210 48.120 336.330 48.400 ;
        RECT 337.170 48.120 347.830 48.400 ;
        RECT 348.670 48.120 359.790 48.400 ;
        RECT 360.630 48.120 371.290 48.400 ;
        RECT 372.130 48.120 383.250 48.400 ;
        RECT 384.090 48.120 394.750 48.400 ;
        RECT 395.590 48.120 406.710 48.400 ;
        RECT 407.550 48.120 409.110 48.400 ;
      LAYER met3 ;
        RECT 53.880 410.960 409.095 411.825 ;
        RECT 53.480 398.760 409.495 410.960 ;
        RECT 53.880 397.360 409.095 398.760 ;
        RECT 53.480 384.480 409.495 397.360 ;
        RECT 53.880 383.080 409.095 384.480 ;
        RECT 53.480 370.880 409.495 383.080 ;
        RECT 53.880 369.480 409.095 370.880 ;
        RECT 53.480 356.600 409.495 369.480 ;
        RECT 53.880 355.200 409.095 356.600 ;
        RECT 53.480 343.000 409.495 355.200 ;
        RECT 53.880 341.600 409.095 343.000 ;
        RECT 53.480 329.400 409.495 341.600 ;
        RECT 53.880 328.000 409.095 329.400 ;
        RECT 53.480 315.120 409.495 328.000 ;
        RECT 53.880 313.720 409.095 315.120 ;
        RECT 53.480 301.520 409.495 313.720 ;
        RECT 53.880 300.120 409.095 301.520 ;
        RECT 53.480 287.240 409.495 300.120 ;
        RECT 53.880 285.840 409.095 287.240 ;
        RECT 53.480 273.640 409.495 285.840 ;
        RECT 53.880 272.240 409.095 273.640 ;
        RECT 53.480 260.040 409.495 272.240 ;
        RECT 53.880 258.640 409.095 260.040 ;
        RECT 53.480 245.760 409.495 258.640 ;
        RECT 53.880 244.360 409.095 245.760 ;
        RECT 53.480 232.160 409.495 244.360 ;
        RECT 53.880 230.760 409.095 232.160 ;
        RECT 53.480 217.880 409.495 230.760 ;
        RECT 53.880 216.480 409.095 217.880 ;
        RECT 53.480 204.280 409.495 216.480 ;
        RECT 53.880 202.880 409.095 204.280 ;
        RECT 53.480 190.680 409.495 202.880 ;
        RECT 53.880 189.280 409.095 190.680 ;
        RECT 53.480 176.400 409.495 189.280 ;
        RECT 53.880 175.000 409.095 176.400 ;
        RECT 53.480 162.800 409.495 175.000 ;
        RECT 53.880 161.400 409.095 162.800 ;
        RECT 53.480 148.520 409.495 161.400 ;
        RECT 53.880 147.120 409.095 148.520 ;
        RECT 53.480 134.920 409.495 147.120 ;
        RECT 53.880 133.520 409.095 134.920 ;
        RECT 53.480 121.320 409.495 133.520 ;
        RECT 53.880 119.920 409.095 121.320 ;
        RECT 53.480 107.040 409.495 119.920 ;
        RECT 53.880 105.640 409.095 107.040 ;
        RECT 53.480 93.440 409.495 105.640 ;
        RECT 53.880 92.040 409.095 93.440 ;
        RECT 53.480 79.160 409.495 92.040 ;
        RECT 53.880 77.760 409.095 79.160 ;
        RECT 53.480 65.560 409.495 77.760 ;
        RECT 53.880 64.160 409.095 65.560 ;
        RECT 53.480 51.960 409.495 64.160 ;
        RECT 53.880 51.095 409.095 51.960 ;
      LAYER met4 ;
        RECT 0.000 0.000 462.820 460.880 ;
      LAYER met5 ;
        RECT 0.000 70.610 462.820 460.880 ;
  END
END clb_tile
END LIBRARY

