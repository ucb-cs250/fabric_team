VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 243.260 BY 253.980 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 249.980 226.230 253.980 ;
    END
  END COUT
  PIN cb_e_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 2.080 243.260 2.680 ;
    END
  END cb_e_clb1_input[0]
  PIN cb_e_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 6.840 243.260 7.440 ;
    END
  END cb_e_clb1_input[1]
  PIN cb_e_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 12.280 243.260 12.880 ;
    END
  END cb_e_clb1_input[2]
  PIN cb_e_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 17.720 243.260 18.320 ;
    END
  END cb_e_clb1_input[3]
  PIN cb_e_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 23.160 243.260 23.760 ;
    END
  END cb_e_clb1_input[4]
  PIN cb_e_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 28.600 243.260 29.200 ;
    END
  END cb_e_clb1_input[5]
  PIN cb_e_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 34.040 243.260 34.640 ;
    END
  END cb_e_clb1_input[6]
  PIN cb_e_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 39.480 243.260 40.080 ;
    END
  END cb_e_clb1_input[7]
  PIN cb_e_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 44.920 243.260 45.520 ;
    END
  END cb_e_clb1_input[8]
  PIN cb_e_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 50.360 243.260 50.960 ;
    END
  END cb_e_clb1_input[9]
  PIN cb_e_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 55.800 243.260 56.400 ;
    END
  END cb_e_clb1_output[0]
  PIN cb_e_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 61.240 243.260 61.840 ;
    END
  END cb_e_clb1_output[1]
  PIN cb_e_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 66.680 243.260 67.280 ;
    END
  END cb_e_clb1_output[2]
  PIN cb_e_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 72.120 243.260 72.720 ;
    END
  END cb_e_clb1_output[3]
  PIN cb_e_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END cb_e_single1_in[0]
  PIN cb_e_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END cb_e_single1_in[10]
  PIN cb_e_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END cb_e_single1_in[11]
  PIN cb_e_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END cb_e_single1_in[12]
  PIN cb_e_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END cb_e_single1_in[13]
  PIN cb_e_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END cb_e_single1_in[14]
  PIN cb_e_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cb_e_single1_in[15]
  PIN cb_e_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END cb_e_single1_in[1]
  PIN cb_e_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END cb_e_single1_in[2]
  PIN cb_e_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END cb_e_single1_in[3]
  PIN cb_e_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END cb_e_single1_in[4]
  PIN cb_e_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END cb_e_single1_in[5]
  PIN cb_e_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END cb_e_single1_in[6]
  PIN cb_e_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END cb_e_single1_in[7]
  PIN cb_e_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END cb_e_single1_in[8]
  PIN cb_e_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END cb_e_single1_in[9]
  PIN cb_e_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cb_e_single1_out[0]
  PIN cb_e_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END cb_e_single1_out[10]
  PIN cb_e_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END cb_e_single1_out[11]
  PIN cb_e_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END cb_e_single1_out[12]
  PIN cb_e_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END cb_e_single1_out[13]
  PIN cb_e_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END cb_e_single1_out[14]
  PIN cb_e_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END cb_e_single1_out[15]
  PIN cb_e_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END cb_e_single1_out[1]
  PIN cb_e_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END cb_e_single1_out[2]
  PIN cb_e_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END cb_e_single1_out[3]
  PIN cb_e_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END cb_e_single1_out[4]
  PIN cb_e_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END cb_e_single1_out[5]
  PIN cb_e_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END cb_e_single1_out[6]
  PIN cb_e_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END cb_e_single1_out[7]
  PIN cb_e_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END cb_e_single1_out[8]
  PIN cb_e_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END cb_e_single1_out[9]
  PIN cb_n_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 249.980 2.670 253.980 ;
    END
  END cb_n_clb1_input[0]
  PIN cb_n_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 249.980 7.270 253.980 ;
    END
  END cb_n_clb1_input[1]
  PIN cb_n_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 249.980 12.330 253.980 ;
    END
  END cb_n_clb1_input[2]
  PIN cb_n_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 249.980 16.930 253.980 ;
    END
  END cb_n_clb1_input[3]
  PIN cb_n_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 249.980 21.990 253.980 ;
    END
  END cb_n_clb1_input[4]
  PIN cb_n_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 249.980 26.590 253.980 ;
    END
  END cb_n_clb1_input[5]
  PIN cb_n_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 249.980 31.650 253.980 ;
    END
  END cb_n_clb1_input[6]
  PIN cb_n_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 249.980 36.710 253.980 ;
    END
  END cb_n_clb1_input[7]
  PIN cb_n_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 249.980 41.310 253.980 ;
    END
  END cb_n_clb1_input[8]
  PIN cb_n_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 249.980 46.370 253.980 ;
    END
  END cb_n_clb1_input[9]
  PIN cb_n_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 249.980 50.970 253.980 ;
    END
  END cb_n_clb1_output[0]
  PIN cb_n_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 249.980 56.030 253.980 ;
    END
  END cb_n_clb1_output[1]
  PIN cb_n_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 249.980 60.630 253.980 ;
    END
  END cb_n_clb1_output[2]
  PIN cb_n_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 249.980 65.690 253.980 ;
    END
  END cb_n_clb1_output[3]
  PIN cb_n_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END cb_n_single1_in[0]
  PIN cb_n_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END cb_n_single1_in[10]
  PIN cb_n_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END cb_n_single1_in[11]
  PIN cb_n_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END cb_n_single1_in[12]
  PIN cb_n_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END cb_n_single1_in[13]
  PIN cb_n_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END cb_n_single1_in[14]
  PIN cb_n_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END cb_n_single1_in[15]
  PIN cb_n_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END cb_n_single1_in[1]
  PIN cb_n_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END cb_n_single1_in[2]
  PIN cb_n_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END cb_n_single1_in[3]
  PIN cb_n_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END cb_n_single1_in[4]
  PIN cb_n_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END cb_n_single1_in[5]
  PIN cb_n_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END cb_n_single1_in[6]
  PIN cb_n_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END cb_n_single1_in[7]
  PIN cb_n_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END cb_n_single1_in[8]
  PIN cb_n_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END cb_n_single1_in[9]
  PIN cb_n_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END cb_n_single1_out[0]
  PIN cb_n_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END cb_n_single1_out[10]
  PIN cb_n_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END cb_n_single1_out[11]
  PIN cb_n_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END cb_n_single1_out[12]
  PIN cb_n_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END cb_n_single1_out[13]
  PIN cb_n_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END cb_n_single1_out[14]
  PIN cb_n_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END cb_n_single1_out[15]
  PIN cb_n_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END cb_n_single1_out[1]
  PIN cb_n_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END cb_n_single1_out[2]
  PIN cb_n_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END cb_n_single1_out[3]
  PIN cb_n_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END cb_n_single1_out[4]
  PIN cb_n_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END cb_n_single1_out[5]
  PIN cb_n_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END cb_n_single1_out[6]
  PIN cb_n_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END cb_n_single1_out[7]
  PIN cb_n_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END cb_n_single1_out[8]
  PIN cb_n_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END cb_n_single1_out[9]
  PIN cfg_bit_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END cfg_bit_in
  PIN cfg_bit_in_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END cfg_bit_in_valid
  PIN cfg_bit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 249.980 235.890 253.980 ;
    END
  END cfg_bit_out
  PIN cfg_bit_out_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 249.980 240.950 253.980 ;
    END
  END cfg_bit_out_valid
  PIN cfg_in_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END cfg_in_start
  PIN cfg_out_start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 249.980 231.290 253.980 ;
    END
  END cfg_out_start
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END clb_south_out[3]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END clb_west_out[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 250.960 243.260 251.560 ;
    END
  END clk
  PIN crst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END crst
  PIN sb_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 77.560 243.260 78.160 ;
    END
  END sb_east_in[0]
  PIN sb_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 131.280 243.260 131.880 ;
    END
  END sb_east_in[10]
  PIN sb_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 136.720 243.260 137.320 ;
    END
  END sb_east_in[11]
  PIN sb_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 142.160 243.260 142.760 ;
    END
  END sb_east_in[12]
  PIN sb_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 147.600 243.260 148.200 ;
    END
  END sb_east_in[13]
  PIN sb_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 153.040 243.260 153.640 ;
    END
  END sb_east_in[14]
  PIN sb_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 158.480 243.260 159.080 ;
    END
  END sb_east_in[15]
  PIN sb_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 83.000 243.260 83.600 ;
    END
  END sb_east_in[1]
  PIN sb_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 88.440 243.260 89.040 ;
    END
  END sb_east_in[2]
  PIN sb_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 93.880 243.260 94.480 ;
    END
  END sb_east_in[3]
  PIN sb_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 99.320 243.260 99.920 ;
    END
  END sb_east_in[4]
  PIN sb_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 104.760 243.260 105.360 ;
    END
  END sb_east_in[5]
  PIN sb_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 110.200 243.260 110.800 ;
    END
  END sb_east_in[6]
  PIN sb_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 115.640 243.260 116.240 ;
    END
  END sb_east_in[7]
  PIN sb_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 121.080 243.260 121.680 ;
    END
  END sb_east_in[8]
  PIN sb_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 126.520 243.260 127.120 ;
    END
  END sb_east_in[9]
  PIN sb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 163.920 243.260 164.520 ;
    END
  END sb_east_out[0]
  PIN sb_east_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 218.320 243.260 218.920 ;
    END
  END sb_east_out[10]
  PIN sb_east_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 223.760 243.260 224.360 ;
    END
  END sb_east_out[11]
  PIN sb_east_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 229.200 243.260 229.800 ;
    END
  END sb_east_out[12]
  PIN sb_east_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 234.640 243.260 235.240 ;
    END
  END sb_east_out[13]
  PIN sb_east_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 240.080 243.260 240.680 ;
    END
  END sb_east_out[14]
  PIN sb_east_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 245.520 243.260 246.120 ;
    END
  END sb_east_out[15]
  PIN sb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 169.360 243.260 169.960 ;
    END
  END sb_east_out[1]
  PIN sb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 174.800 243.260 175.400 ;
    END
  END sb_east_out[2]
  PIN sb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 180.240 243.260 180.840 ;
    END
  END sb_east_out[3]
  PIN sb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 185.680 243.260 186.280 ;
    END
  END sb_east_out[4]
  PIN sb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 191.120 243.260 191.720 ;
    END
  END sb_east_out[5]
  PIN sb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 196.560 243.260 197.160 ;
    END
  END sb_east_out[6]
  PIN sb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 202.000 243.260 202.600 ;
    END
  END sb_east_out[7]
  PIN sb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 207.440 243.260 208.040 ;
    END
  END sb_east_out[8]
  PIN sb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.260 212.880 243.260 213.480 ;
    END
  END sb_east_out[9]
  PIN sb_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 249.980 70.750 253.980 ;
    END
  END sb_north_in[0]
  PIN sb_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 249.980 119.050 253.980 ;
    END
  END sb_north_in[10]
  PIN sb_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 249.980 124.110 253.980 ;
    END
  END sb_north_in[11]
  PIN sb_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 249.980 129.170 253.980 ;
    END
  END sb_north_in[12]
  PIN sb_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 249.980 133.770 253.980 ;
    END
  END sb_north_in[13]
  PIN sb_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 249.980 138.830 253.980 ;
    END
  END sb_north_in[14]
  PIN sb_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 249.980 143.430 253.980 ;
    END
  END sb_north_in[15]
  PIN sb_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 249.980 75.350 253.980 ;
    END
  END sb_north_in[1]
  PIN sb_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 249.980 80.410 253.980 ;
    END
  END sb_north_in[2]
  PIN sb_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 249.980 85.010 253.980 ;
    END
  END sb_north_in[3]
  PIN sb_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 249.980 90.070 253.980 ;
    END
  END sb_north_in[4]
  PIN sb_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 249.980 95.130 253.980 ;
    END
  END sb_north_in[5]
  PIN sb_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 249.980 99.730 253.980 ;
    END
  END sb_north_in[6]
  PIN sb_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 249.980 104.790 253.980 ;
    END
  END sb_north_in[7]
  PIN sb_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 249.980 109.390 253.980 ;
    END
  END sb_north_in[8]
  PIN sb_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 249.980 114.450 253.980 ;
    END
  END sb_north_in[9]
  PIN sb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 249.980 148.490 253.980 ;
    END
  END sb_north_out[0]
  PIN sb_north_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 249.980 197.250 253.980 ;
    END
  END sb_north_out[10]
  PIN sb_north_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 249.980 201.850 253.980 ;
    END
  END sb_north_out[11]
  PIN sb_north_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 249.980 206.910 253.980 ;
    END
  END sb_north_out[12]
  PIN sb_north_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 249.980 211.510 253.980 ;
    END
  END sb_north_out[13]
  PIN sb_north_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 249.980 216.570 253.980 ;
    END
  END sb_north_out[14]
  PIN sb_north_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 249.980 221.630 253.980 ;
    END
  END sb_north_out[15]
  PIN sb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 249.980 153.090 253.980 ;
    END
  END sb_north_out[1]
  PIN sb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 249.980 158.150 253.980 ;
    END
  END sb_north_out[2]
  PIN sb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 249.980 163.210 253.980 ;
    END
  END sb_north_out[3]
  PIN sb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 249.980 167.810 253.980 ;
    END
  END sb_north_out[4]
  PIN sb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 249.980 172.870 253.980 ;
    END
  END sb_north_out[5]
  PIN sb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 249.980 177.470 253.980 ;
    END
  END sb_north_out[6]
  PIN sb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 249.980 182.530 253.980 ;
    END
  END sb_north_out[7]
  PIN sb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 249.980 187.590 253.980 ;
    END
  END sb_north_out[8]
  PIN sb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 249.980 192.190 253.980 ;
    END
  END sb_north_out[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 242.320 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 242.320 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 242.320 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 7.565 237.360 242.165 ;
      LAYER met1 ;
        RECT 2.370 6.160 240.970 242.320 ;
      LAYER met2 ;
        RECT 2.950 249.700 6.710 251.445 ;
        RECT 7.550 249.700 11.770 251.445 ;
        RECT 12.610 249.700 16.370 251.445 ;
        RECT 17.210 249.700 21.430 251.445 ;
        RECT 22.270 249.700 26.030 251.445 ;
        RECT 26.870 249.700 31.090 251.445 ;
        RECT 31.930 249.700 36.150 251.445 ;
        RECT 36.990 249.700 40.750 251.445 ;
        RECT 41.590 249.700 45.810 251.445 ;
        RECT 46.650 249.700 50.410 251.445 ;
        RECT 51.250 249.700 55.470 251.445 ;
        RECT 56.310 249.700 60.070 251.445 ;
        RECT 60.910 249.700 65.130 251.445 ;
        RECT 65.970 249.700 70.190 251.445 ;
        RECT 71.030 249.700 74.790 251.445 ;
        RECT 75.630 249.700 79.850 251.445 ;
        RECT 80.690 249.700 84.450 251.445 ;
        RECT 85.290 249.700 89.510 251.445 ;
        RECT 90.350 249.700 94.570 251.445 ;
        RECT 95.410 249.700 99.170 251.445 ;
        RECT 100.010 249.700 104.230 251.445 ;
        RECT 105.070 249.700 108.830 251.445 ;
        RECT 109.670 249.700 113.890 251.445 ;
        RECT 114.730 249.700 118.490 251.445 ;
        RECT 119.330 249.700 123.550 251.445 ;
        RECT 124.390 249.700 128.610 251.445 ;
        RECT 129.450 249.700 133.210 251.445 ;
        RECT 134.050 249.700 138.270 251.445 ;
        RECT 139.110 249.700 142.870 251.445 ;
        RECT 143.710 249.700 147.930 251.445 ;
        RECT 148.770 249.700 152.530 251.445 ;
        RECT 153.370 249.700 157.590 251.445 ;
        RECT 158.430 249.700 162.650 251.445 ;
        RECT 163.490 249.700 167.250 251.445 ;
        RECT 168.090 249.700 172.310 251.445 ;
        RECT 173.150 249.700 176.910 251.445 ;
        RECT 177.750 249.700 181.970 251.445 ;
        RECT 182.810 249.700 187.030 251.445 ;
        RECT 187.870 249.700 191.630 251.445 ;
        RECT 192.470 249.700 196.690 251.445 ;
        RECT 197.530 249.700 201.290 251.445 ;
        RECT 202.130 249.700 206.350 251.445 ;
        RECT 207.190 249.700 210.950 251.445 ;
        RECT 211.790 249.700 216.010 251.445 ;
        RECT 216.850 249.700 221.070 251.445 ;
        RECT 221.910 249.700 225.670 251.445 ;
        RECT 226.510 249.700 230.730 251.445 ;
        RECT 231.570 249.700 235.330 251.445 ;
        RECT 236.170 249.700 240.390 251.445 ;
        RECT 2.400 4.280 240.940 249.700 ;
        RECT 2.950 2.195 6.710 4.280 ;
        RECT 7.550 2.195 11.310 4.280 ;
        RECT 12.150 2.195 16.370 4.280 ;
        RECT 17.210 2.195 20.970 4.280 ;
        RECT 21.810 2.195 25.570 4.280 ;
        RECT 26.410 2.195 30.630 4.280 ;
        RECT 31.470 2.195 35.230 4.280 ;
        RECT 36.070 2.195 39.830 4.280 ;
        RECT 40.670 2.195 44.890 4.280 ;
        RECT 45.730 2.195 49.490 4.280 ;
        RECT 50.330 2.195 54.550 4.280 ;
        RECT 55.390 2.195 59.150 4.280 ;
        RECT 59.990 2.195 63.750 4.280 ;
        RECT 64.590 2.195 68.810 4.280 ;
        RECT 69.650 2.195 73.410 4.280 ;
        RECT 74.250 2.195 78.010 4.280 ;
        RECT 78.850 2.195 83.070 4.280 ;
        RECT 83.910 2.195 87.670 4.280 ;
        RECT 88.510 2.195 92.730 4.280 ;
        RECT 93.570 2.195 97.330 4.280 ;
        RECT 98.170 2.195 101.930 4.280 ;
        RECT 102.770 2.195 106.990 4.280 ;
        RECT 107.830 2.195 111.590 4.280 ;
        RECT 112.430 2.195 116.190 4.280 ;
        RECT 117.030 2.195 121.250 4.280 ;
        RECT 122.090 2.195 125.850 4.280 ;
        RECT 126.690 2.195 130.910 4.280 ;
        RECT 131.750 2.195 135.510 4.280 ;
        RECT 136.350 2.195 140.110 4.280 ;
        RECT 140.950 2.195 145.170 4.280 ;
        RECT 146.010 2.195 149.770 4.280 ;
        RECT 150.610 2.195 154.370 4.280 ;
        RECT 155.210 2.195 159.430 4.280 ;
        RECT 160.270 2.195 164.030 4.280 ;
        RECT 164.870 2.195 169.090 4.280 ;
        RECT 169.930 2.195 173.690 4.280 ;
        RECT 174.530 2.195 178.290 4.280 ;
        RECT 179.130 2.195 183.350 4.280 ;
        RECT 184.190 2.195 187.950 4.280 ;
        RECT 188.790 2.195 192.550 4.280 ;
        RECT 193.390 2.195 197.610 4.280 ;
        RECT 198.450 2.195 202.210 4.280 ;
        RECT 203.050 2.195 207.270 4.280 ;
        RECT 208.110 2.195 211.870 4.280 ;
        RECT 212.710 2.195 216.470 4.280 ;
        RECT 217.310 2.195 221.530 4.280 ;
        RECT 222.370 2.195 226.130 4.280 ;
        RECT 226.970 2.195 230.730 4.280 ;
        RECT 231.570 2.195 235.790 4.280 ;
        RECT 236.630 2.195 240.390 4.280 ;
      LAYER met3 ;
        RECT 4.400 250.560 238.860 251.425 ;
        RECT 4.000 246.520 239.260 250.560 ;
        RECT 4.400 245.120 238.860 246.520 ;
        RECT 4.000 241.080 239.260 245.120 ;
        RECT 4.400 239.680 238.860 241.080 ;
        RECT 4.000 235.640 239.260 239.680 ;
        RECT 4.400 234.240 238.860 235.640 ;
        RECT 4.000 230.200 239.260 234.240 ;
        RECT 4.400 228.800 238.860 230.200 ;
        RECT 4.000 224.760 239.260 228.800 ;
        RECT 4.400 223.360 238.860 224.760 ;
        RECT 4.000 219.320 239.260 223.360 ;
        RECT 4.400 217.920 238.860 219.320 ;
        RECT 4.000 213.880 239.260 217.920 ;
        RECT 4.000 213.200 238.860 213.880 ;
        RECT 4.400 212.480 238.860 213.200 ;
        RECT 4.400 211.800 239.260 212.480 ;
        RECT 4.000 208.440 239.260 211.800 ;
        RECT 4.000 207.760 238.860 208.440 ;
        RECT 4.400 207.040 238.860 207.760 ;
        RECT 4.400 206.360 239.260 207.040 ;
        RECT 4.000 203.000 239.260 206.360 ;
        RECT 4.000 202.320 238.860 203.000 ;
        RECT 4.400 201.600 238.860 202.320 ;
        RECT 4.400 200.920 239.260 201.600 ;
        RECT 4.000 197.560 239.260 200.920 ;
        RECT 4.000 196.880 238.860 197.560 ;
        RECT 4.400 196.160 238.860 196.880 ;
        RECT 4.400 195.480 239.260 196.160 ;
        RECT 4.000 192.120 239.260 195.480 ;
        RECT 4.000 191.440 238.860 192.120 ;
        RECT 4.400 190.720 238.860 191.440 ;
        RECT 4.400 190.040 239.260 190.720 ;
        RECT 4.000 186.680 239.260 190.040 ;
        RECT 4.000 186.000 238.860 186.680 ;
        RECT 4.400 185.280 238.860 186.000 ;
        RECT 4.400 184.600 239.260 185.280 ;
        RECT 4.000 181.240 239.260 184.600 ;
        RECT 4.000 180.560 238.860 181.240 ;
        RECT 4.400 179.840 238.860 180.560 ;
        RECT 4.400 179.160 239.260 179.840 ;
        RECT 4.000 175.800 239.260 179.160 ;
        RECT 4.000 175.120 238.860 175.800 ;
        RECT 4.400 174.400 238.860 175.120 ;
        RECT 4.400 173.720 239.260 174.400 ;
        RECT 4.000 170.360 239.260 173.720 ;
        RECT 4.000 169.000 238.860 170.360 ;
        RECT 4.400 168.960 238.860 169.000 ;
        RECT 4.400 167.600 239.260 168.960 ;
        RECT 4.000 164.920 239.260 167.600 ;
        RECT 4.000 163.560 238.860 164.920 ;
        RECT 4.400 163.520 238.860 163.560 ;
        RECT 4.400 162.160 239.260 163.520 ;
        RECT 4.000 159.480 239.260 162.160 ;
        RECT 4.000 158.120 238.860 159.480 ;
        RECT 4.400 158.080 238.860 158.120 ;
        RECT 4.400 156.720 239.260 158.080 ;
        RECT 4.000 154.040 239.260 156.720 ;
        RECT 4.000 152.680 238.860 154.040 ;
        RECT 4.400 152.640 238.860 152.680 ;
        RECT 4.400 151.280 239.260 152.640 ;
        RECT 4.000 148.600 239.260 151.280 ;
        RECT 4.000 147.240 238.860 148.600 ;
        RECT 4.400 147.200 238.860 147.240 ;
        RECT 4.400 145.840 239.260 147.200 ;
        RECT 4.000 143.160 239.260 145.840 ;
        RECT 4.000 141.800 238.860 143.160 ;
        RECT 4.400 141.760 238.860 141.800 ;
        RECT 4.400 140.400 239.260 141.760 ;
        RECT 4.000 137.720 239.260 140.400 ;
        RECT 4.000 136.360 238.860 137.720 ;
        RECT 4.400 136.320 238.860 136.360 ;
        RECT 4.400 134.960 239.260 136.320 ;
        RECT 4.000 132.280 239.260 134.960 ;
        RECT 4.000 130.920 238.860 132.280 ;
        RECT 4.400 130.880 238.860 130.920 ;
        RECT 4.400 129.520 239.260 130.880 ;
        RECT 4.000 127.520 239.260 129.520 ;
        RECT 4.000 126.120 238.860 127.520 ;
        RECT 4.000 124.800 239.260 126.120 ;
        RECT 4.400 123.400 239.260 124.800 ;
        RECT 4.000 122.080 239.260 123.400 ;
        RECT 4.000 120.680 238.860 122.080 ;
        RECT 4.000 119.360 239.260 120.680 ;
        RECT 4.400 117.960 239.260 119.360 ;
        RECT 4.000 116.640 239.260 117.960 ;
        RECT 4.000 115.240 238.860 116.640 ;
        RECT 4.000 113.920 239.260 115.240 ;
        RECT 4.400 112.520 239.260 113.920 ;
        RECT 4.000 111.200 239.260 112.520 ;
        RECT 4.000 109.800 238.860 111.200 ;
        RECT 4.000 108.480 239.260 109.800 ;
        RECT 4.400 107.080 239.260 108.480 ;
        RECT 4.000 105.760 239.260 107.080 ;
        RECT 4.000 104.360 238.860 105.760 ;
        RECT 4.000 103.040 239.260 104.360 ;
        RECT 4.400 101.640 239.260 103.040 ;
        RECT 4.000 100.320 239.260 101.640 ;
        RECT 4.000 98.920 238.860 100.320 ;
        RECT 4.000 97.600 239.260 98.920 ;
        RECT 4.400 96.200 239.260 97.600 ;
        RECT 4.000 94.880 239.260 96.200 ;
        RECT 4.000 93.480 238.860 94.880 ;
        RECT 4.000 92.160 239.260 93.480 ;
        RECT 4.400 90.760 239.260 92.160 ;
        RECT 4.000 89.440 239.260 90.760 ;
        RECT 4.000 88.040 238.860 89.440 ;
        RECT 4.000 86.040 239.260 88.040 ;
        RECT 4.400 84.640 239.260 86.040 ;
        RECT 4.000 84.000 239.260 84.640 ;
        RECT 4.000 82.600 238.860 84.000 ;
        RECT 4.000 80.600 239.260 82.600 ;
        RECT 4.400 79.200 239.260 80.600 ;
        RECT 4.000 78.560 239.260 79.200 ;
        RECT 4.000 77.160 238.860 78.560 ;
        RECT 4.000 75.160 239.260 77.160 ;
        RECT 4.400 73.760 239.260 75.160 ;
        RECT 4.000 73.120 239.260 73.760 ;
        RECT 4.000 71.720 238.860 73.120 ;
        RECT 4.000 69.720 239.260 71.720 ;
        RECT 4.400 68.320 239.260 69.720 ;
        RECT 4.000 67.680 239.260 68.320 ;
        RECT 4.000 66.280 238.860 67.680 ;
        RECT 4.000 64.280 239.260 66.280 ;
        RECT 4.400 62.880 239.260 64.280 ;
        RECT 4.000 62.240 239.260 62.880 ;
        RECT 4.000 60.840 238.860 62.240 ;
        RECT 4.000 58.840 239.260 60.840 ;
        RECT 4.400 57.440 239.260 58.840 ;
        RECT 4.000 56.800 239.260 57.440 ;
        RECT 4.000 55.400 238.860 56.800 ;
        RECT 4.000 53.400 239.260 55.400 ;
        RECT 4.400 52.000 239.260 53.400 ;
        RECT 4.000 51.360 239.260 52.000 ;
        RECT 4.000 49.960 238.860 51.360 ;
        RECT 4.000 47.960 239.260 49.960 ;
        RECT 4.400 46.560 239.260 47.960 ;
        RECT 4.000 45.920 239.260 46.560 ;
        RECT 4.000 44.520 238.860 45.920 ;
        RECT 4.000 41.840 239.260 44.520 ;
        RECT 4.400 40.480 239.260 41.840 ;
        RECT 4.400 40.440 238.860 40.480 ;
        RECT 4.000 39.080 238.860 40.440 ;
        RECT 4.000 36.400 239.260 39.080 ;
        RECT 4.400 35.040 239.260 36.400 ;
        RECT 4.400 35.000 238.860 35.040 ;
        RECT 4.000 33.640 238.860 35.000 ;
        RECT 4.000 30.960 239.260 33.640 ;
        RECT 4.400 29.600 239.260 30.960 ;
        RECT 4.400 29.560 238.860 29.600 ;
        RECT 4.000 28.200 238.860 29.560 ;
        RECT 4.000 25.520 239.260 28.200 ;
        RECT 4.400 24.160 239.260 25.520 ;
        RECT 4.400 24.120 238.860 24.160 ;
        RECT 4.000 22.760 238.860 24.120 ;
        RECT 4.000 20.080 239.260 22.760 ;
        RECT 4.400 18.720 239.260 20.080 ;
        RECT 4.400 18.680 238.860 18.720 ;
        RECT 4.000 17.320 238.860 18.680 ;
        RECT 4.000 14.640 239.260 17.320 ;
        RECT 4.400 13.280 239.260 14.640 ;
        RECT 4.400 13.240 238.860 13.280 ;
        RECT 4.000 11.880 238.860 13.240 ;
        RECT 4.000 9.200 239.260 11.880 ;
        RECT 4.400 7.840 239.260 9.200 ;
        RECT 4.400 7.800 238.860 7.840 ;
        RECT 4.000 6.440 238.860 7.800 ;
        RECT 4.000 3.760 239.260 6.440 ;
        RECT 4.400 3.080 239.260 3.760 ;
        RECT 4.400 2.360 238.860 3.080 ;
        RECT 4.000 2.215 238.860 2.360 ;
      LAYER met4 ;
        RECT 13.175 12.415 20.640 239.865 ;
        RECT 23.040 12.415 97.440 239.865 ;
        RECT 99.840 12.415 174.240 239.865 ;
        RECT 176.640 12.415 231.545 239.865 ;
  END
END clb_tile
END LIBRARY

