VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block
  CLASS BLOCK ;
  FOREIGN baked_connection_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 242.560 BY 253.280 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 6.840 242.560 7.440 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 21.120 242.560 21.720 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 36.080 242.560 36.680 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 51.040 242.560 51.640 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 66.000 242.560 66.600 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 80.960 242.560 81.560 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 95.920 242.560 96.520 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 110.880 242.560 111.480 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 125.840 242.560 126.440 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 140.120 242.560 140.720 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 155.080 242.560 155.680 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 238.560 170.040 242.560 170.640 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 185.000 242.560 185.600 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 199.960 242.560 200.560 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 214.920 242.560 215.520 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 229.880 242.560 230.480 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 244.840 242.560 245.440 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.150 249.280 189.430 253.280 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 249.280 67.990 253.280 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 249.280 83.170 253.280 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 249.280 98.350 253.280 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 249.280 113.530 253.280 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 128.430 249.280 128.710 253.280 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 249.280 143.890 253.280 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 249.280 159.070 253.280 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 249.280 174.250 253.280 ;
    END
  END double1[7]
  PIN global[-1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END global[-1]
  PIN global[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 204.330 249.280 204.610 253.280 ;
    END
  END global[0]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.510 249.280 219.790 253.280 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.690 249.280 234.970 253.280 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 249.280 7.730 253.280 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 249.280 22.450 253.280 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 249.280 37.630 253.280 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 249.280 52.810 253.280 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 242.320 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 242.320 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 236.900 242.165 ;
      LAYER met1 ;
        RECT 5.520 10.640 236.900 242.320 ;
      LAYER met2 ;
        RECT 7.000 249.000 7.170 249.280 ;
        RECT 8.010 249.000 21.890 249.280 ;
        RECT 22.730 249.000 37.070 249.280 ;
        RECT 37.910 249.000 52.250 249.280 ;
        RECT 53.090 249.000 67.430 249.280 ;
        RECT 68.270 249.000 82.610 249.280 ;
        RECT 83.450 249.000 97.790 249.280 ;
        RECT 98.630 249.000 112.970 249.280 ;
        RECT 113.810 249.000 128.150 249.280 ;
        RECT 128.990 249.000 143.330 249.280 ;
        RECT 144.170 249.000 158.510 249.280 ;
        RECT 159.350 249.000 173.690 249.280 ;
        RECT 174.530 249.000 188.870 249.280 ;
        RECT 189.710 249.000 204.050 249.280 ;
        RECT 204.890 249.000 219.230 249.280 ;
        RECT 220.070 249.000 234.410 249.280 ;
        RECT 7.000 4.280 234.960 249.000 ;
        RECT 7.000 4.000 7.170 4.280 ;
        RECT 8.010 4.000 21.890 4.280 ;
        RECT 22.730 4.000 37.070 4.280 ;
        RECT 37.910 4.000 52.250 4.280 ;
        RECT 53.090 4.000 67.430 4.280 ;
        RECT 68.270 4.000 82.610 4.280 ;
        RECT 83.450 4.000 97.790 4.280 ;
        RECT 98.630 4.000 112.970 4.280 ;
        RECT 113.810 4.000 128.150 4.280 ;
        RECT 128.990 4.000 143.330 4.280 ;
        RECT 144.170 4.000 158.510 4.280 ;
        RECT 159.350 4.000 173.690 4.280 ;
        RECT 174.530 4.000 188.870 4.280 ;
        RECT 189.710 4.000 204.050 4.280 ;
        RECT 204.890 4.000 219.230 4.280 ;
        RECT 220.070 4.000 234.410 4.280 ;
      LAYER met3 ;
        RECT 4.400 244.440 238.160 245.305 ;
        RECT 4.000 230.880 238.560 244.440 ;
        RECT 4.400 229.480 238.160 230.880 ;
        RECT 4.000 215.920 238.560 229.480 ;
        RECT 4.400 214.520 238.160 215.920 ;
        RECT 4.000 200.960 238.560 214.520 ;
        RECT 4.400 199.560 238.160 200.960 ;
        RECT 4.000 186.000 238.560 199.560 ;
        RECT 4.400 184.600 238.160 186.000 ;
        RECT 4.000 171.040 238.560 184.600 ;
        RECT 4.400 169.640 238.160 171.040 ;
        RECT 4.000 156.080 238.560 169.640 ;
        RECT 4.400 154.680 238.160 156.080 ;
        RECT 4.000 141.120 238.560 154.680 ;
        RECT 4.400 139.720 238.160 141.120 ;
        RECT 4.000 126.840 238.560 139.720 ;
        RECT 4.400 125.440 238.160 126.840 ;
        RECT 4.000 111.880 238.560 125.440 ;
        RECT 4.400 110.480 238.160 111.880 ;
        RECT 4.000 96.920 238.560 110.480 ;
        RECT 4.400 95.520 238.160 96.920 ;
        RECT 4.000 81.960 238.560 95.520 ;
        RECT 4.400 80.560 238.160 81.960 ;
        RECT 4.000 67.000 238.560 80.560 ;
        RECT 4.400 65.600 238.160 67.000 ;
        RECT 4.000 52.040 238.560 65.600 ;
        RECT 4.400 50.640 238.160 52.040 ;
        RECT 4.000 37.080 238.560 50.640 ;
        RECT 4.400 35.680 238.160 37.080 ;
        RECT 4.000 22.120 238.560 35.680 ;
        RECT 4.400 20.720 238.160 22.120 ;
        RECT 4.000 7.840 238.560 20.720 ;
        RECT 4.400 6.975 238.160 7.840 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 242.320 ;
  END
END baked_connection_block
END LIBRARY

