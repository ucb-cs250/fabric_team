magic
tech sky130A
magscale 1 2
timestamp 1623787548
<< locali >>
rect 7573 11067 7607 11237
rect 489 3723 523 4233
rect 673 3587 707 5117
rect 765 3179 799 9333
rect 857 3383 891 9469
rect 6193 7735 6227 7973
rect 8861 7939 8895 8041
rect 8585 7191 8619 7293
rect 7113 6103 7147 6341
rect 765 3145 891 3179
rect 673 1819 707 3009
rect 765 1887 799 3077
rect 857 2091 891 3145
rect 949 1955 983 5729
rect 3433 5627 3467 5729
rect 9781 2839 9815 3145
<< viali >>
rect 4169 12937 4203 12971
rect 6193 12937 6227 12971
rect 7757 12937 7791 12971
rect 7941 12937 7975 12971
rect 9873 12937 9907 12971
rect 11345 12937 11379 12971
rect 8585 12869 8619 12903
rect 11069 12869 11103 12903
rect 3341 12801 3375 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 1961 12733 1995 12767
rect 2513 12733 2547 12767
rect 2789 12733 2823 12767
rect 3065 12733 3099 12767
rect 3525 12733 3559 12767
rect 4353 12733 4387 12767
rect 4629 12733 4663 12767
rect 4997 12733 5031 12767
rect 5549 12733 5583 12767
rect 5641 12733 5675 12767
rect 6101 12733 6135 12767
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 7205 12733 7239 12767
rect 8133 12733 8167 12767
rect 8493 12733 8527 12767
rect 8585 12733 8619 12767
rect 8769 12733 8803 12767
rect 9045 12733 9079 12767
rect 9321 12733 9355 12767
rect 9781 12733 9815 12767
rect 10057 12733 10091 12767
rect 10517 12733 10551 12767
rect 10885 12733 10919 12767
rect 11713 12733 11747 12767
rect 2329 12665 2363 12699
rect 7665 12665 7699 12699
rect 8309 12665 8343 12699
rect 11253 12665 11287 12699
rect 1777 12597 1811 12631
rect 2145 12597 2179 12631
rect 2697 12597 2731 12631
rect 2973 12597 3007 12631
rect 4905 12597 4939 12631
rect 5365 12597 5399 12631
rect 6561 12597 6595 12631
rect 8861 12597 8895 12631
rect 9413 12597 9447 12631
rect 10333 12597 10367 12631
rect 11529 12597 11563 12631
rect 5273 12393 5307 12427
rect 8217 12393 8251 12427
rect 8493 12393 8527 12427
rect 9137 12393 9171 12427
rect 3709 12325 3743 12359
rect 4160 12325 4194 12359
rect 9965 12325 9999 12359
rect 10394 12325 10428 12359
rect 1676 12257 1710 12291
rect 2881 12257 2915 12291
rect 3525 12257 3559 12291
rect 5365 12257 5399 12291
rect 5632 12257 5666 12291
rect 6837 12257 6871 12291
rect 7093 12257 7127 12291
rect 8585 12257 8619 12291
rect 8769 12257 8803 12291
rect 9321 12257 9355 12291
rect 9873 12257 9907 12291
rect 10057 12257 10091 12291
rect 11621 12257 11655 12291
rect 1409 12189 1443 12223
rect 3893 12189 3927 12223
rect 9597 12189 9631 12223
rect 10149 12189 10183 12223
rect 6745 12121 6779 12155
rect 2789 12053 2823 12087
rect 8309 12053 8343 12087
rect 9505 12053 9539 12087
rect 11529 12053 11563 12087
rect 4537 11849 4571 11883
rect 5089 11849 5123 11883
rect 6653 11849 6687 11883
rect 9137 11849 9171 11883
rect 9413 11849 9447 11883
rect 10149 11849 10183 11883
rect 10241 11849 10275 11883
rect 11253 11849 11287 11883
rect 1685 11781 1719 11815
rect 7205 11781 7239 11815
rect 2145 11713 2179 11747
rect 2329 11713 2363 11747
rect 4997 11713 5031 11747
rect 5181 11713 5215 11747
rect 6745 11713 6779 11747
rect 10333 11713 10367 11747
rect 1409 11645 1443 11679
rect 2053 11645 2087 11679
rect 2513 11645 2547 11679
rect 4169 11645 4203 11679
rect 4445 11645 4479 11679
rect 4905 11645 4939 11679
rect 5273 11645 5307 11679
rect 5733 11645 5767 11679
rect 6009 11645 6043 11679
rect 6285 11645 6319 11679
rect 6469 11645 6503 11679
rect 6561 11645 6595 11679
rect 6837 11645 6871 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 8024 11645 8058 11679
rect 9321 11645 9355 11679
rect 9689 11645 9723 11679
rect 9965 11645 9999 11679
rect 10057 11645 10091 11679
rect 10425 11645 10459 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 11161 11645 11195 11679
rect 11437 11645 11471 11679
rect 2780 11577 2814 11611
rect 5365 11577 5399 11611
rect 6929 11577 6963 11611
rect 10517 11577 10551 11611
rect 1501 11509 1535 11543
rect 3893 11509 3927 11543
rect 3985 11509 4019 11543
rect 5549 11509 5583 11543
rect 5825 11509 5859 11543
rect 6101 11509 6135 11543
rect 7481 11509 7515 11543
rect 10977 11509 11011 11543
rect 1685 11305 1719 11339
rect 2789 11305 2823 11339
rect 3065 11305 3099 11339
rect 5457 11305 5491 11339
rect 7941 11305 7975 11339
rect 10149 11305 10183 11339
rect 1869 11237 1903 11271
rect 4169 11237 4203 11271
rect 6346 11237 6380 11271
rect 7573 11237 7607 11271
rect 7849 11237 7883 11271
rect 8493 11237 8527 11271
rect 8709 11237 8743 11271
rect 9965 11237 9999 11271
rect 1409 11169 1443 11203
rect 1777 11169 1811 11203
rect 2145 11169 2179 11203
rect 2329 11169 2363 11203
rect 2513 11169 2547 11203
rect 2881 11169 2915 11203
rect 3341 11169 3375 11203
rect 3525 11169 3559 11203
rect 3893 11169 3927 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 5089 11169 5123 11203
rect 5181 11169 5215 11203
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6101 11169 6135 11203
rect 1685 11101 1719 11135
rect 2237 11101 2271 11135
rect 2789 11101 2823 11135
rect 3433 11101 3467 11135
rect 4169 11101 4203 11135
rect 8125 11169 8159 11203
rect 9137 11169 9171 11203
rect 9689 11169 9723 11203
rect 9873 11169 9907 11203
rect 10609 11169 10643 11203
rect 10698 11169 10732 11203
rect 10793 11169 10827 11203
rect 10977 11169 11011 11203
rect 11069 11169 11103 11203
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 9781 11101 9815 11135
rect 10149 11101 10183 11135
rect 11161 11101 11195 11135
rect 3985 11033 4019 11067
rect 4261 11033 4295 11067
rect 7481 11033 7515 11067
rect 7573 11033 7607 11067
rect 8217 11033 8251 11067
rect 9321 11033 9355 11067
rect 1501 10965 1535 10999
rect 2605 10965 2639 10999
rect 4537 10965 4571 10999
rect 4905 10965 4939 10999
rect 5273 10965 5307 10999
rect 5917 10965 5951 10999
rect 8677 10965 8711 10999
rect 8861 10965 8895 10999
rect 10333 10965 10367 10999
rect 11345 10965 11379 10999
rect 1409 10761 1443 10795
rect 5549 10761 5583 10795
rect 5825 10761 5859 10795
rect 6561 10761 6595 10795
rect 8861 10761 8895 10795
rect 9505 10761 9539 10795
rect 11529 10761 11563 10795
rect 2605 10693 2639 10727
rect 7205 10693 7239 10727
rect 2053 10625 2087 10659
rect 3617 10625 3651 10659
rect 3709 10625 3743 10659
rect 6285 10625 6319 10659
rect 7297 10625 7331 10659
rect 9781 10625 9815 10659
rect 10149 10625 10183 10659
rect 1777 10557 1811 10591
rect 1869 10557 1903 10591
rect 2329 10557 2363 10591
rect 2513 10557 2547 10591
rect 2789 10557 2823 10591
rect 3065 10557 3099 10591
rect 3985 10557 4019 10591
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 5739 10557 5773 10591
rect 5917 10557 5951 10591
rect 6009 10557 6043 10591
rect 6101 10557 6135 10591
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 6929 10557 6963 10591
rect 7021 10557 7055 10591
rect 7564 10557 7598 10591
rect 9045 10557 9079 10591
rect 9321 10557 9355 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 11897 10557 11931 10591
rect 4252 10489 4286 10523
rect 10416 10489 10450 10523
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 3157 10421 3191 10455
rect 3525 10421 3559 10455
rect 5365 10421 5399 10455
rect 6285 10421 6319 10455
rect 6745 10421 6779 10455
rect 8677 10421 8711 10455
rect 9229 10421 9263 10455
rect 11713 10421 11747 10455
rect 4721 10217 4755 10251
rect 9505 10217 9539 10251
rect 9965 10217 9999 10251
rect 10425 10217 10459 10251
rect 1685 10149 1719 10183
rect 2022 10149 2056 10183
rect 5816 10149 5850 10183
rect 1409 10081 1443 10115
rect 1501 10081 1535 10115
rect 3433 10081 3467 10115
rect 3525 10081 3559 10115
rect 4077 10081 4111 10115
rect 4353 10081 4387 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 7113 10081 7147 10115
rect 7481 10081 7515 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 8059 10081 8093 10115
rect 8493 10081 8527 10115
rect 8769 10081 8803 10115
rect 8953 10081 8987 10115
rect 9137 10081 9171 10115
rect 9781 10081 9815 10115
rect 10241 10081 10275 10115
rect 10425 10081 10459 10115
rect 10609 10081 10643 10115
rect 10876 10081 10910 10115
rect 1685 10013 1719 10047
rect 1777 10013 1811 10047
rect 7389 10013 7423 10047
rect 3157 9945 3191 9979
rect 3893 9945 3927 9979
rect 3249 9877 3283 9911
rect 3617 9877 3651 9911
rect 4169 9877 4203 9911
rect 4905 9877 4939 9911
rect 5181 9877 5215 9911
rect 6929 9877 6963 9911
rect 7205 9877 7239 9911
rect 7297 9877 7331 9911
rect 7849 9877 7883 9911
rect 8769 9877 8803 9911
rect 9505 9877 9539 9911
rect 9689 9877 9723 9911
rect 11989 9877 12023 9911
rect 3249 9673 3283 9707
rect 4445 9673 4479 9707
rect 5733 9673 5767 9707
rect 6929 9673 6963 9707
rect 8769 9673 8803 9707
rect 10609 9673 10643 9707
rect 10793 9673 10827 9707
rect 1961 9605 1995 9639
rect 2881 9605 2915 9639
rect 3433 9605 3467 9639
rect 4353 9605 4387 9639
rect 5365 9605 5399 9639
rect 8493 9605 8527 9639
rect 2513 9537 2547 9571
rect 3985 9537 4019 9571
rect 4537 9537 4571 9571
rect 4813 9537 4847 9571
rect 857 9469 891 9503
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 3157 9469 3191 9503
rect 4261 9469 4295 9503
rect 4721 9469 4755 9503
rect 4905 9469 4939 9503
rect 5181 9469 5215 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 5825 9469 5859 9503
rect 6009 9469 6043 9503
rect 6201 9469 6235 9503
rect 6469 9469 6503 9503
rect 6837 9469 6871 9503
rect 7113 9469 7147 9503
rect 7380 9469 7414 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 9689 9469 9723 9503
rect 10885 9469 10919 9503
rect 11529 9469 11563 9503
rect 11897 9469 11931 9503
rect 765 9333 799 9367
rect 673 5117 707 5151
rect 489 4233 523 4267
rect 489 3689 523 3723
rect 673 3553 707 3587
rect 3801 9401 3835 9435
rect 3893 9401 3927 9435
rect 6101 9401 6135 9435
rect 9965 9401 9999 9435
rect 10149 9401 10183 9435
rect 10333 9401 10367 9435
rect 10425 9401 10459 9435
rect 10641 9401 10675 9435
rect 1409 9333 1443 9367
rect 1685 9333 1719 9367
rect 2421 9333 2455 9367
rect 4997 9333 5031 9367
rect 2789 9129 2823 9163
rect 3617 9129 3651 9163
rect 6561 9129 6595 9163
rect 6653 9129 6687 9163
rect 8401 9129 8435 9163
rect 9137 9129 9171 9163
rect 9597 9129 9631 9163
rect 3508 9061 3542 9095
rect 4160 9061 4194 9095
rect 5825 9061 5859 9095
rect 9965 9061 9999 9095
rect 10333 9061 10367 9095
rect 10425 9061 10459 9095
rect 10641 9061 10675 9095
rect 10977 9061 11011 9095
rect 1409 8993 1443 9027
rect 1676 8993 1710 9027
rect 3065 8993 3099 9027
rect 3341 8993 3375 9027
rect 5733 8993 5767 9027
rect 7021 8993 7055 9027
rect 7196 8993 7230 9027
rect 7297 8993 7331 9027
rect 7573 8993 7607 9027
rect 8033 8993 8067 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 8677 8993 8711 9027
rect 9505 8993 9539 9027
rect 10149 8993 10183 9027
rect 10885 8993 10919 9027
rect 11069 8993 11103 9027
rect 3893 8925 3927 8959
rect 6009 8925 6043 8959
rect 6837 8925 6871 8959
rect 8861 8925 8895 8959
rect 9781 8925 9815 8959
rect 5365 8857 5399 8891
rect 7113 8857 7147 8891
rect 11621 8857 11655 8891
rect 2881 8789 2915 8823
rect 3157 8789 3191 8823
rect 5273 8789 5307 8823
rect 6193 8789 6227 8823
rect 10609 8789 10643 8823
rect 10793 8789 10827 8823
rect 11345 8789 11379 8823
rect 11897 8789 11931 8823
rect 1409 8585 1443 8619
rect 1869 8585 1903 8619
rect 4261 8585 4295 8619
rect 8401 8585 8435 8619
rect 8953 8585 8987 8619
rect 9413 8585 9447 8619
rect 11253 8585 11287 8619
rect 1777 8517 1811 8551
rect 6101 8517 6135 8551
rect 1961 8449 1995 8483
rect 2421 8449 2455 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5641 8449 5675 8483
rect 6929 8449 6963 8483
rect 10149 8449 10183 8483
rect 1593 8381 1627 8415
rect 1685 8381 1719 8415
rect 2237 8381 2271 8415
rect 2329 8381 2363 8415
rect 2513 8381 2547 8415
rect 2605 8381 2639 8415
rect 2881 8381 2915 8415
rect 4905 8381 4939 8415
rect 5365 8381 5399 8415
rect 5457 8381 5491 8415
rect 6653 8381 6687 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 8493 8381 8527 8415
rect 8861 8381 8895 8415
rect 9229 8381 9263 8415
rect 9781 8381 9815 8415
rect 9873 8381 9907 8415
rect 11897 8381 11931 8415
rect 3126 8313 3160 8347
rect 5917 8313 5951 8347
rect 6929 8313 6963 8347
rect 7266 8313 7300 8347
rect 2053 8245 2087 8279
rect 4537 8245 4571 8279
rect 5641 8245 5675 8279
rect 1961 8041 1995 8075
rect 2513 8041 2547 8075
rect 3065 8041 3099 8075
rect 4537 8041 4571 8075
rect 6377 8041 6411 8075
rect 8401 8041 8435 8075
rect 8861 8041 8895 8075
rect 2053 7973 2087 8007
rect 3985 7973 4019 8007
rect 4988 7973 5022 8007
rect 6193 7973 6227 8007
rect 2421 7905 2455 7939
rect 2789 7905 2823 7939
rect 2881 7905 2915 7939
rect 3249 7905 3283 7939
rect 3433 7905 3467 7939
rect 3525 7905 3559 7939
rect 4445 7905 4479 7939
rect 2145 7837 2179 7871
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 4721 7837 4755 7871
rect 1593 7769 1627 7803
rect 10600 7973 10634 8007
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 7021 7905 7055 7939
rect 7665 7905 7699 7939
rect 7941 7905 7975 7939
rect 8861 7905 8895 7939
rect 9137 7905 9171 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 6653 7837 6687 7871
rect 7205 7837 7239 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10241 7837 10275 7871
rect 10333 7837 10367 7871
rect 9229 7769 9263 7803
rect 4077 7701 4111 7735
rect 6101 7701 6135 7735
rect 6193 7701 6227 7735
rect 7113 7701 7147 7735
rect 8033 7701 8067 7735
rect 9321 7701 9355 7735
rect 9965 7701 9999 7735
rect 11713 7701 11747 7735
rect 11989 7701 12023 7735
rect 2053 7497 2087 7531
rect 2697 7497 2731 7531
rect 3985 7497 4019 7531
rect 5181 7497 5215 7531
rect 6193 7497 6227 7531
rect 8401 7497 8435 7531
rect 10057 7497 10091 7531
rect 10425 7497 10459 7531
rect 3525 7429 3559 7463
rect 3617 7429 3651 7463
rect 7941 7429 7975 7463
rect 10333 7429 10367 7463
rect 3709 7361 3743 7395
rect 5365 7361 5399 7395
rect 5825 7361 5859 7395
rect 8677 7361 8711 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 11345 7361 11379 7395
rect 1501 7293 1535 7327
rect 1777 7293 1811 7327
rect 2237 7293 2271 7327
rect 2513 7293 2547 7327
rect 2605 7293 2639 7327
rect 3249 7293 3283 7327
rect 3433 7293 3467 7327
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 4813 7293 4847 7327
rect 5089 7293 5123 7327
rect 5457 7293 5491 7327
rect 5733 7293 5767 7327
rect 5925 7293 5959 7327
rect 8309 7293 8343 7327
rect 8493 7293 8527 7327
rect 8585 7293 8619 7327
rect 8944 7293 8978 7327
rect 10241 7293 10275 7327
rect 10609 7293 10643 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 11897 7293 11931 7327
rect 3893 7225 3927 7259
rect 6101 7225 6135 7259
rect 6469 7225 6503 7259
rect 10701 7225 10735 7259
rect 2329 7157 2363 7191
rect 3065 7157 3099 7191
rect 5365 7157 5399 7191
rect 8585 7157 8619 7191
rect 3249 6953 3283 6987
rect 6745 6953 6779 6987
rect 8861 6953 8895 6987
rect 9229 6953 9263 6987
rect 9781 6953 9815 6987
rect 9873 6953 9907 6987
rect 10609 6953 10643 6987
rect 10701 6953 10735 6987
rect 7104 6885 7138 6919
rect 8677 6885 8711 6919
rect 1409 6817 1443 6851
rect 1676 6817 1710 6851
rect 3341 6817 3375 6851
rect 3893 6817 3927 6851
rect 4160 6817 4194 6851
rect 5365 6817 5399 6851
rect 5632 6817 5666 6851
rect 8493 6817 8527 6851
rect 8769 6817 8803 6851
rect 9137 6817 9171 6851
rect 11069 6817 11103 6851
rect 3433 6749 3467 6783
rect 6837 6749 6871 6783
rect 9965 6749 9999 6783
rect 10793 6749 10827 6783
rect 11529 6749 11563 6783
rect 2881 6681 2915 6715
rect 8217 6681 8251 6715
rect 9413 6681 9447 6715
rect 10241 6681 10275 6715
rect 2789 6613 2823 6647
rect 5273 6613 5307 6647
rect 11161 6613 11195 6647
rect 11805 6613 11839 6647
rect 1593 6409 1627 6443
rect 3709 6409 3743 6443
rect 3985 6409 4019 6443
rect 5917 6409 5951 6443
rect 6561 6409 6595 6443
rect 7205 6409 7239 6443
rect 8217 6409 8251 6443
rect 2697 6341 2731 6375
rect 4997 6341 5031 6375
rect 7113 6341 7147 6375
rect 1685 6273 1719 6307
rect 2329 6273 2363 6307
rect 5457 6273 5491 6307
rect 5641 6273 5675 6307
rect 6745 6273 6779 6307
rect 1409 6205 1443 6239
rect 1501 6205 1535 6239
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 3065 6205 3099 6239
rect 3341 6205 3375 6239
rect 3617 6205 3651 6239
rect 3893 6205 3927 6239
rect 4077 6205 4111 6239
rect 4169 6205 4203 6239
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 5365 6205 5399 6239
rect 5825 6205 5859 6239
rect 6101 6205 6135 6239
rect 6469 6205 6503 6239
rect 6837 6205 6871 6239
rect 6929 6137 6963 6171
rect 7757 6273 7791 6307
rect 8493 6273 8527 6307
rect 10149 6273 10183 6307
rect 7573 6205 7607 6239
rect 8033 6205 8067 6239
rect 11713 6205 11747 6239
rect 11897 6205 11931 6239
rect 8760 6137 8794 6171
rect 10416 6137 10450 6171
rect 1777 6069 1811 6103
rect 2145 6069 2179 6103
rect 2237 6069 2271 6103
rect 6745 6069 6779 6103
rect 7113 6069 7147 6103
rect 7665 6069 7699 6103
rect 9873 6069 9907 6103
rect 11529 6069 11563 6103
rect 11805 6069 11839 6103
rect 1777 5865 1811 5899
rect 2421 5865 2455 5899
rect 3893 5865 3927 5899
rect 5733 5865 5767 5899
rect 7941 5865 7975 5899
rect 8125 5865 8159 5899
rect 10701 5865 10735 5899
rect 4261 5797 4295 5831
rect 5273 5797 5307 5831
rect 6101 5797 6135 5831
rect 6193 5797 6227 5831
rect 6806 5797 6840 5831
rect 8953 5797 8987 5831
rect 11069 5797 11103 5831
rect 857 3349 891 3383
rect 949 5729 983 5763
rect 1593 5729 1627 5763
rect 1685 5729 1719 5763
rect 2973 5729 3007 5763
rect 3065 5729 3099 5763
rect 3433 5729 3467 5763
rect 3525 5729 3559 5763
rect 4721 5729 4755 5763
rect 5089 5729 5123 5763
rect 6561 5729 6595 5763
rect 8033 5729 8067 5763
rect 8217 5729 8251 5763
rect 8401 5729 8435 5763
rect 8585 5729 8619 5763
rect 8677 5729 8711 5763
rect 9137 5729 9171 5763
rect 9597 5729 9631 5763
rect 9781 5729 9815 5763
rect 9873 5729 9907 5763
rect 10425 5729 10459 5763
rect 10885 5729 10919 5763
rect 11897 5729 11931 5763
rect 765 3077 799 3111
rect 673 3009 707 3043
rect 857 2057 891 2091
rect 2513 5661 2547 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 4353 5661 4387 5695
rect 4537 5661 4571 5695
rect 6377 5661 6411 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 9689 5661 9723 5695
rect 10149 5661 10183 5695
rect 10701 5661 10735 5695
rect 1409 5593 1443 5627
rect 3433 5593 3467 5627
rect 10517 5593 10551 5627
rect 11345 5593 11379 5627
rect 2053 5525 2087 5559
rect 3157 5525 3191 5559
rect 5641 5525 5675 5559
rect 8769 5525 8803 5559
rect 9965 5525 9999 5559
rect 10057 5525 10091 5559
rect 11621 5525 11655 5559
rect 2789 5321 2823 5355
rect 4537 5321 4571 5355
rect 6285 5321 6319 5355
rect 8677 5321 8711 5355
rect 9597 5321 9631 5355
rect 11529 5321 11563 5355
rect 2973 5253 3007 5287
rect 5273 5253 5307 5287
rect 7481 5253 7515 5287
rect 7113 5185 7147 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 9137 5185 9171 5219
rect 9321 5185 9355 5219
rect 10149 5185 10183 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 3157 5117 3191 5151
rect 3413 5117 3447 5151
rect 4629 5117 4663 5151
rect 5641 5117 5675 5151
rect 5825 5117 5859 5151
rect 7389 5117 7423 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 8401 5117 8435 5151
rect 9045 5117 9079 5151
rect 9505 5117 9539 5151
rect 10416 5117 10450 5151
rect 11805 5117 11839 5151
rect 1676 5049 1710 5083
rect 5089 5049 5123 5083
rect 5457 5049 5491 5083
rect 7021 5049 7055 5083
rect 9873 5049 9907 5083
rect 11989 5049 12023 5083
rect 4813 4981 4847 5015
rect 5917 4981 5951 5015
rect 6561 4981 6595 5015
rect 6929 4981 6963 5015
rect 7665 4981 7699 5015
rect 8125 4981 8159 5015
rect 9965 4981 9999 5015
rect 2421 4777 2455 4811
rect 4353 4777 4387 4811
rect 8677 4777 8711 4811
rect 9137 4777 9171 4811
rect 10425 4777 10459 4811
rect 10793 4777 10827 4811
rect 2605 4709 2639 4743
rect 4905 4709 4939 4743
rect 6728 4709 6762 4743
rect 7564 4709 7598 4743
rect 9597 4709 9631 4743
rect 10057 4709 10091 4743
rect 11437 4709 11471 4743
rect 1501 4641 1535 4675
rect 1869 4641 1903 4675
rect 2145 4641 2179 4675
rect 2513 4641 2547 4675
rect 2789 4641 2823 4675
rect 2973 4641 3007 4675
rect 3249 4641 3283 4675
rect 3525 4641 3559 4675
rect 3985 4641 4019 4675
rect 4169 4641 4203 4675
rect 4261 4641 4295 4675
rect 4445 4641 4479 4675
rect 5437 4641 5471 4675
rect 7021 4641 7055 4675
rect 7297 4641 7331 4675
rect 8769 4641 8803 4675
rect 9505 4641 9539 4675
rect 11805 4641 11839 4675
rect 2421 4573 2455 4607
rect 2881 4573 2915 4607
rect 5181 4573 5215 4607
rect 9689 4573 9723 4607
rect 10885 4573 10919 4607
rect 10977 4573 11011 4607
rect 4721 4505 4755 4539
rect 6929 4505 6963 4539
rect 11989 4505 12023 4539
rect 1593 4437 1627 4471
rect 2237 4437 2271 4471
rect 4077 4437 4111 4471
rect 4997 4437 5031 4471
rect 6561 4437 6595 4471
rect 7113 4437 7147 4471
rect 8861 4437 8895 4471
rect 10149 4437 10183 4471
rect 11529 4437 11563 4471
rect 2237 4233 2271 4267
rect 3433 4233 3467 4267
rect 5457 4233 5491 4267
rect 5733 4233 5767 4267
rect 6653 4233 6687 4267
rect 7573 4233 7607 4267
rect 6009 4165 6043 4199
rect 9045 4165 9079 4199
rect 2789 4097 2823 4131
rect 3620 4097 3654 4131
rect 6561 4097 6595 4131
rect 6748 4097 6782 4131
rect 7389 4097 7423 4131
rect 8493 4097 8527 4131
rect 9229 4097 9263 4131
rect 11161 4097 11195 4131
rect 1685 4029 1719 4063
rect 2605 4029 2639 4063
rect 2697 4029 2731 4063
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 3341 4029 3375 4063
rect 3709 4029 3743 4063
rect 6285 4029 6319 4063
rect 6469 4029 6503 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7481 4029 7515 4063
rect 7941 4029 7975 4063
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 8953 4029 8987 4063
rect 9321 4029 9355 4063
rect 10977 4029 11011 4063
rect 11345 4029 11379 4063
rect 11805 4029 11839 4063
rect 1501 3961 1535 3995
rect 1869 3961 1903 3995
rect 3617 3961 3651 3995
rect 3954 3961 3988 3995
rect 6929 3961 6963 3995
rect 8309 3961 8343 3995
rect 9229 3961 9263 3995
rect 9566 3961 9600 3995
rect 11529 3961 11563 3995
rect 1961 3893 1995 3927
rect 3157 3893 3191 3927
rect 5089 3893 5123 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 10701 3893 10735 3927
rect 11897 3893 11931 3927
rect 2789 3689 2823 3723
rect 3985 3689 4019 3723
rect 7389 3689 7423 3723
rect 7757 3689 7791 3723
rect 10793 3689 10827 3723
rect 1676 3621 1710 3655
rect 3157 3621 3191 3655
rect 5273 3621 5307 3655
rect 6653 3621 6687 3655
rect 8769 3621 8803 3655
rect 9229 3621 9263 3655
rect 9597 3621 9631 3655
rect 9965 3621 9999 3655
rect 10333 3621 10367 3655
rect 10701 3621 10735 3655
rect 11437 3621 11471 3655
rect 11621 3621 11655 3655
rect 1409 3553 1443 3587
rect 2881 3553 2915 3587
rect 2973 3553 3007 3587
rect 3249 3553 3283 3587
rect 3525 3553 3559 3587
rect 3893 3553 3927 3587
rect 4169 3553 4203 3587
rect 4353 3553 4387 3587
rect 4721 3553 4755 3587
rect 4813 3553 4847 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 5457 3553 5491 3587
rect 5641 3553 5675 3587
rect 6193 3553 6227 3587
rect 6561 3553 6595 3587
rect 8217 3553 8251 3587
rect 11069 3553 11103 3587
rect 11805 3553 11839 3587
rect 3157 3485 3191 3519
rect 5089 3485 5123 3519
rect 5549 3485 5583 3519
rect 6469 3485 6503 3519
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 8493 3485 8527 3519
rect 8953 3485 8987 3519
rect 9413 3485 9447 3519
rect 10517 3485 10551 3519
rect 11253 3485 11287 3519
rect 3617 3417 3651 3451
rect 6101 3417 6135 3451
rect 7021 3417 7055 3451
rect 10149 3417 10183 3451
rect 11989 3417 12023 3451
rect 3341 3349 3375 3383
rect 4261 3349 4295 3383
rect 4997 3349 5031 3383
rect 6285 3349 6319 3383
rect 6377 3349 6411 3383
rect 7297 3349 7331 3383
rect 8309 3349 8343 3383
rect 8401 3349 8435 3383
rect 9689 3349 9723 3383
rect 2697 3145 2731 3179
rect 3893 3145 3927 3179
rect 8953 3145 8987 3179
rect 9781 3145 9815 3179
rect 10149 3145 10183 3179
rect 3617 3077 3651 3111
rect 6469 3077 6503 3111
rect 3249 3009 3283 3043
rect 3801 3009 3835 3043
rect 4445 3009 4479 3043
rect 4813 3009 4847 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 9321 3009 9355 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 2145 2941 2179 2975
rect 2605 2941 2639 2975
rect 3157 2941 3191 2975
rect 3525 2941 3559 2975
rect 5080 2941 5114 2975
rect 6837 2941 6871 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 7840 2941 7874 2975
rect 9137 2941 9171 2975
rect 3065 2873 3099 2907
rect 4261 2873 4295 2907
rect 9505 2873 9539 2907
rect 10609 3077 10643 3111
rect 10977 3009 11011 3043
rect 10057 2941 10091 2975
rect 10793 2941 10827 2975
rect 11989 2941 12023 2975
rect 10408 2873 10442 2907
rect 11161 2873 11195 2907
rect 11805 2873 11839 2907
rect 3801 2805 3835 2839
rect 4353 2805 4387 2839
rect 6193 2805 6227 2839
rect 9597 2805 9631 2839
rect 9781 2805 9815 2839
rect 11253 2805 11287 2839
rect 3341 2601 3375 2635
rect 5365 2601 5399 2635
rect 6285 2601 6319 2635
rect 7941 2601 7975 2635
rect 8953 2601 8987 2635
rect 10149 2601 10183 2635
rect 4160 2533 4194 2567
rect 6806 2533 6840 2567
rect 8401 2533 8435 2567
rect 8493 2533 8527 2567
rect 9321 2533 9355 2567
rect 10701 2533 10735 2567
rect 11069 2533 11103 2567
rect 11437 2533 11471 2567
rect 1593 2465 1627 2499
rect 1961 2465 1995 2499
rect 2145 2465 2179 2499
rect 2697 2465 2731 2499
rect 3433 2465 3467 2499
rect 3893 2465 3927 2499
rect 5733 2465 5767 2499
rect 5825 2465 5859 2499
rect 6193 2465 6227 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 8861 2465 8895 2499
rect 9689 2465 9723 2499
rect 9965 2465 9999 2499
rect 10149 2465 10183 2499
rect 10333 2465 10367 2499
rect 3525 2397 3559 2431
rect 6009 2397 6043 2431
rect 8585 2397 8619 2431
rect 11621 2397 11655 2431
rect 2789 2329 2823 2363
rect 2973 2329 3007 2363
rect 5273 2329 5307 2363
rect 8033 2329 8067 2363
rect 10517 2329 10551 2363
rect 9413 2261 9447 2295
rect 9781 2261 9815 2295
rect 10793 2261 10827 2295
rect 11161 2261 11195 2295
rect 949 1921 983 1955
rect 765 1853 799 1887
rect 673 1785 707 1819
<< metal1 >>
rect 566 13404 572 13456
rect 624 13444 630 13456
rect 9030 13444 9036 13456
rect 624 13416 9036 13444
rect 624 13404 630 13416
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 658 13336 664 13388
rect 716 13376 722 13388
rect 7282 13376 7288 13388
rect 716 13348 7288 13376
rect 716 13336 722 13348
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 1210 13268 1216 13320
rect 1268 13308 1274 13320
rect 6270 13308 6276 13320
rect 1268 13280 6276 13308
rect 1268 13268 1274 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 1118 13200 1124 13252
rect 1176 13240 1182 13252
rect 5534 13240 5540 13252
rect 1176 13212 5540 13240
rect 1176 13200 1182 13212
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 2682 13132 2688 13184
rect 2740 13172 2746 13184
rect 7926 13172 7932 13184
rect 2740 13144 7932 13172
rect 2740 13132 2746 13144
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 1104 13082 12328 13104
rect 1104 13030 2852 13082
rect 2904 13030 2916 13082
rect 2968 13030 2980 13082
rect 3032 13030 3044 13082
rect 3096 13030 6594 13082
rect 6646 13030 6658 13082
rect 6710 13030 6722 13082
rect 6774 13030 6786 13082
rect 6838 13030 10335 13082
rect 10387 13030 10399 13082
rect 10451 13030 10463 13082
rect 10515 13030 10527 13082
rect 10579 13030 12328 13082
rect 1104 13008 12328 13030
rect 934 12928 940 12980
rect 992 12968 998 12980
rect 4157 12971 4215 12977
rect 4157 12968 4169 12971
rect 992 12940 4169 12968
rect 992 12928 998 12940
rect 4157 12937 4169 12940
rect 4203 12937 4215 12971
rect 4157 12931 4215 12937
rect 750 12860 756 12912
rect 808 12900 814 12912
rect 808 12872 3464 12900
rect 808 12860 814 12872
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 1360 12804 3341 12832
rect 1360 12792 1366 12804
rect 2792 12773 2820 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 1949 12767 2007 12773
rect 1949 12764 1961 12767
rect 1780 12736 1961 12764
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1780 12637 1808 12736
rect 1949 12733 1961 12736
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 3053 12767 3111 12773
rect 2823 12736 2857 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3436 12764 3464 12872
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3099 12736 3525 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3513 12733 3525 12736
rect 3559 12733 3571 12767
rect 4172 12764 4200 12931
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5224 12940 6193 12968
rect 5224 12928 5230 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 6972 12940 7757 12968
rect 6972 12928 6978 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7745 12931 7803 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8076 12940 9628 12968
rect 8076 12928 8082 12940
rect 8202 12900 8208 12912
rect 7208 12872 8208 12900
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4580 12804 4721 12832
rect 4580 12792 4586 12804
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 5258 12832 5264 12844
rect 4939 12804 5264 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 6638 12832 6644 12844
rect 5368 12804 6644 12832
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4172 12736 4353 12764
rect 3513 12727 3571 12733
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4614 12764 4620 12776
rect 4575 12736 4620 12764
rect 4341 12727 4399 12733
rect 1854 12656 1860 12708
rect 1912 12696 1918 12708
rect 2317 12699 2375 12705
rect 2317 12696 2329 12699
rect 1912 12668 2329 12696
rect 1912 12656 1918 12668
rect 2317 12665 2329 12668
rect 2363 12696 2375 12699
rect 2516 12696 2544 12727
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5074 12764 5080 12776
rect 5031 12736 5080 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5368 12764 5396 12804
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 7208 12776 7236 12872
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 8573 12903 8631 12909
rect 8573 12900 8585 12903
rect 8352 12872 8585 12900
rect 8352 12860 8358 12872
rect 8573 12869 8585 12872
rect 8619 12869 8631 12903
rect 9600 12900 9628 12940
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9732 12940 9873 12968
rect 9732 12928 9738 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11204 12940 11345 12968
rect 11204 12928 11210 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 11057 12903 11115 12909
rect 9600 12872 10548 12900
rect 8573 12863 8631 12869
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 10520 12832 10548 12872
rect 11057 12869 11069 12903
rect 11103 12900 11115 12903
rect 12618 12900 12624 12912
rect 11103 12872 12624 12900
rect 11103 12869 11115 12872
rect 11057 12863 11115 12869
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 7984 12804 9812 12832
rect 7984 12792 7990 12804
rect 5534 12764 5540 12776
rect 5224 12736 5396 12764
rect 5495 12736 5540 12764
rect 5224 12724 5230 12736
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5684 12736 6101 12764
rect 5684 12724 5690 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6733 12767 6791 12773
rect 6733 12764 6745 12767
rect 6328 12736 6745 12764
rect 6328 12724 6334 12736
rect 6733 12733 6745 12736
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 7190 12764 7196 12776
rect 7103 12736 7196 12764
rect 6825 12727 6883 12733
rect 2363 12668 2544 12696
rect 2363 12665 2375 12668
rect 2317 12659 2375 12665
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3476 12668 5580 12696
rect 3476 12656 3482 12668
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1636 12600 1777 12628
rect 1636 12588 1642 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 1765 12591 1823 12597
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 2096 12600 2145 12628
rect 2096 12588 2102 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2133 12591 2191 12597
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2648 12600 2697 12628
rect 2648 12588 2654 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 2961 12631 3019 12637
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 3234 12628 3240 12640
rect 3007 12600 3240 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4304 12600 4905 12628
rect 4304 12588 4310 12600
rect 4893 12597 4905 12600
rect 4939 12597 4951 12631
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 4893 12591 4951 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 5552 12628 5580 12668
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 6840 12696 6868 12727
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 8121 12767 8179 12773
rect 8121 12764 8133 12767
rect 7340 12736 8133 12764
rect 7340 12724 7346 12736
rect 8121 12733 8133 12736
rect 8167 12733 8179 12767
rect 8121 12727 8179 12733
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8444 12736 8493 12764
rect 8444 12724 8450 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 8754 12764 8760 12776
rect 8715 12736 8760 12764
rect 8573 12727 8631 12733
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 6236 12668 7665 12696
rect 6236 12656 6242 12668
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 8297 12699 8355 12705
rect 8297 12696 8309 12699
rect 8260 12668 8309 12696
rect 8260 12656 8266 12668
rect 8297 12665 8309 12668
rect 8343 12665 8355 12699
rect 8588 12696 8616 12727
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9784 12773 9812 12804
rect 10520 12804 11744 12832
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 9180 12736 9321 12764
rect 9180 12724 9186 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 9769 12727 9827 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10520 12773 10548 12804
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12764 10931 12767
rect 10962 12764 10968 12776
rect 10919 12736 10968 12764
rect 10919 12733 10931 12736
rect 10873 12727 10931 12733
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11716 12773 11744 12804
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 8938 12696 8944 12708
rect 8588 12668 8944 12696
rect 8297 12659 8355 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 11146 12696 11152 12708
rect 10336 12668 11152 12696
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 5552 12600 6561 12628
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 8849 12631 8907 12637
rect 8849 12628 8861 12631
rect 6696 12600 8861 12628
rect 6696 12588 6702 12600
rect 8849 12597 8861 12600
rect 8895 12597 8907 12631
rect 8849 12591 8907 12597
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 10336 12637 10364 12668
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 11606 12696 11612 12708
rect 11287 12668 11612 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 9364 12600 9413 12628
rect 9364 12588 9370 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12597 10379 12631
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 10321 12591 10379 12597
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 1104 12538 12328 12560
rect 1104 12486 4723 12538
rect 4775 12486 4787 12538
rect 4839 12486 4851 12538
rect 4903 12486 4915 12538
rect 4967 12486 8464 12538
rect 8516 12486 8528 12538
rect 8580 12486 8592 12538
rect 8644 12486 8656 12538
rect 8708 12486 12328 12538
rect 1104 12464 12328 12486
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 5132 12396 5273 12424
rect 5132 12384 5138 12396
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 6362 12424 6368 12436
rect 5684 12396 6368 12424
rect 5684 12384 5690 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 8202 12424 8208 12436
rect 6472 12396 7880 12424
rect 8163 12396 8208 12424
rect 3694 12356 3700 12368
rect 3655 12328 3700 12356
rect 3694 12316 3700 12328
rect 3752 12316 3758 12368
rect 4148 12359 4206 12365
rect 4148 12325 4160 12359
rect 4194 12356 4206 12359
rect 4246 12356 4252 12368
rect 4194 12328 4252 12356
rect 4194 12325 4206 12328
rect 4148 12319 4206 12325
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5166 12356 5172 12368
rect 4764 12328 5172 12356
rect 4764 12316 4770 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 6472 12356 6500 12396
rect 7742 12356 7748 12368
rect 5368 12328 6500 12356
rect 6840 12328 7748 12356
rect 1670 12297 1676 12300
rect 1664 12251 1676 12297
rect 1728 12288 1734 12300
rect 1728 12260 1764 12288
rect 1670 12248 1676 12251
rect 1728 12248 1734 12260
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2869 12291 2927 12297
rect 2869 12288 2881 12291
rect 2464 12260 2881 12288
rect 2464 12248 2470 12260
rect 2869 12257 2881 12260
rect 2915 12257 2927 12291
rect 2869 12251 2927 12257
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12288 3571 12291
rect 4430 12288 4436 12300
rect 3559 12260 4436 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2884 12220 2912 12251
rect 4430 12248 4436 12260
rect 4488 12288 4494 12300
rect 4982 12288 4988 12300
rect 4488 12260 4988 12288
rect 4488 12248 4494 12260
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5368 12297 5396 12328
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5620 12291 5678 12297
rect 5620 12257 5632 12291
rect 5666 12288 5678 12291
rect 5902 12288 5908 12300
rect 5666 12260 5908 12288
rect 5666 12257 5678 12260
rect 5620 12251 5678 12257
rect 3694 12220 3700 12232
rect 2884 12192 3700 12220
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2777 12087 2835 12093
rect 2777 12084 2789 12087
rect 2188 12056 2789 12084
rect 2188 12044 2194 12056
rect 2777 12053 2789 12056
rect 2823 12053 2835 12087
rect 2777 12047 2835 12053
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3896 12084 3924 12183
rect 5368 12084 5396 12251
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6840 12297 6868 12328
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 7852 12356 7880 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 8754 12424 8760 12436
rect 8527 12396 8760 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8996 12396 9137 12424
rect 8996 12384 9002 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9214 12384 9220 12436
rect 9272 12424 9278 12436
rect 11606 12424 11612 12436
rect 9272 12396 11612 12424
rect 9272 12384 9278 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 9766 12356 9772 12368
rect 7852 12328 9772 12356
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9953 12359 10011 12365
rect 9953 12325 9965 12359
rect 9999 12356 10011 12359
rect 10382 12359 10440 12365
rect 10382 12356 10394 12359
rect 9999 12328 10394 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 10382 12325 10394 12328
rect 10428 12325 10440 12359
rect 10382 12319 10440 12325
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7081 12291 7139 12297
rect 7081 12288 7093 12291
rect 6972 12260 7093 12288
rect 6972 12248 6978 12260
rect 7081 12257 7093 12260
rect 7127 12257 7139 12291
rect 7081 12251 7139 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 8938 12288 8944 12300
rect 8803 12260 8944 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 8588 12220 8616 12251
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9306 12288 9312 12300
rect 9267 12260 9312 12288
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9858 12288 9864 12300
rect 9819 12260 9864 12288
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 11606 12288 11612 12300
rect 11567 12260 11612 12288
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 9398 12220 9404 12232
rect 8588 12192 9404 12220
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 9582 12220 9588 12232
rect 9543 12192 9588 12220
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 6733 12155 6791 12161
rect 6733 12152 6745 12155
rect 6420 12124 6745 12152
rect 6420 12112 6426 12124
rect 6733 12121 6745 12124
rect 6779 12121 6791 12155
rect 6733 12115 6791 12121
rect 3660 12056 5396 12084
rect 3660 12044 3666 12056
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 8168 12056 8309 12084
rect 8168 12044 8174 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 8297 12047 8355 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 10836 12056 11529 12084
rect 10836 12044 10842 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11517 12047 11575 12053
rect 1104 11994 12328 12016
rect 1104 11942 2852 11994
rect 2904 11942 2916 11994
rect 2968 11942 2980 11994
rect 3032 11942 3044 11994
rect 3096 11942 6594 11994
rect 6646 11942 6658 11994
rect 6710 11942 6722 11994
rect 6774 11942 6786 11994
rect 6838 11942 10335 11994
rect 10387 11942 10399 11994
rect 10451 11942 10463 11994
rect 10515 11942 10527 11994
rect 10579 11942 12328 11994
rect 1104 11920 12328 11942
rect 106 11840 112 11892
rect 164 11880 170 11892
rect 4525 11883 4583 11889
rect 164 11852 4200 11880
rect 164 11840 170 11852
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11781 1731 11815
rect 2406 11812 2412 11824
rect 1673 11775 1731 11781
rect 2332 11784 2412 11812
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1688 11676 1716 11775
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2332 11753 2360 11784
rect 2406 11772 2412 11784
rect 2464 11772 2470 11824
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2424 11716 2636 11744
rect 1443 11648 1716 11676
rect 2041 11679 2099 11685
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2424 11676 2452 11716
rect 2087 11648 2452 11676
rect 2501 11679 2559 11685
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 2608 11676 2636 11716
rect 4172 11685 4200 11852
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 4614 11880 4620 11892
rect 4571 11852 4620 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5902 11880 5908 11892
rect 5123 11852 5908 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 6914 11880 6920 11892
rect 6687 11852 6920 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 9548 11852 10149 11880
rect 9548 11840 9554 11852
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 11238 11880 11244 11892
rect 10284 11852 10329 11880
rect 11199 11852 11244 11880
rect 10284 11840 10290 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 5350 11812 5356 11824
rect 4264 11784 5356 11812
rect 4157 11679 4215 11685
rect 2608 11648 4108 11676
rect 2501 11639 2559 11645
rect 2516 11608 2544 11639
rect 2774 11617 2780 11620
rect 1412 11580 2544 11608
rect 1412 11552 1440 11580
rect 1394 11500 1400 11552
rect 1452 11500 1458 11552
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 2038 11540 2044 11552
rect 1535 11512 2044 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2516 11540 2544 11580
rect 2768 11571 2780 11617
rect 2832 11608 2838 11620
rect 3602 11608 3608 11620
rect 2832 11580 2868 11608
rect 2976 11580 3608 11608
rect 2774 11568 2780 11571
rect 2832 11568 2838 11580
rect 2976 11540 3004 11580
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 4080 11608 4108 11648
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4264 11608 4292 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 7193 11815 7251 11821
rect 7193 11812 7205 11815
rect 5500 11784 7205 11812
rect 5500 11772 5506 11784
rect 7193 11781 7205 11784
rect 7239 11781 7251 11815
rect 7193 11775 7251 11781
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 9508 11812 9536 11840
rect 8996 11784 9536 11812
rect 9692 11784 10640 11812
rect 8996 11772 9002 11784
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4580 11716 4997 11744
rect 4580 11704 4586 11716
rect 4985 11713 4997 11716
rect 5031 11744 5043 11747
rect 5074 11744 5080 11756
rect 5031 11716 5080 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5534 11744 5540 11756
rect 5215 11716 5540 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 5868 11716 6316 11744
rect 5868 11704 5874 11716
rect 4430 11676 4436 11688
rect 4391 11648 4436 11676
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11676 5319 11679
rect 5718 11676 5724 11688
rect 5307 11648 5488 11676
rect 5679 11648 5724 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 4080 11580 4292 11608
rect 4908 11608 4936 11639
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 4908 11580 5365 11608
rect 5353 11577 5365 11580
rect 5399 11577 5411 11611
rect 5460 11608 5488 11648
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 5994 11676 6000 11688
rect 5955 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6288 11685 6316 11716
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6420 11716 6745 11744
rect 6420 11704 6426 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 9692 11688 9720 11784
rect 10321 11747 10379 11753
rect 9968 11716 10180 11744
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 6457 11679 6515 11685
rect 6457 11645 6469 11679
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 5626 11608 5632 11620
rect 5460 11580 5632 11608
rect 5353 11571 5411 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6472 11608 6500 11639
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 6825 11679 6883 11685
rect 6604 11648 6649 11676
rect 6604 11636 6610 11648
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7190 11676 7196 11688
rect 6871 11648 7196 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7650 11676 7656 11688
rect 7611 11648 7656 11676
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 8012 11679 8070 11685
rect 7800 11648 7893 11676
rect 7800 11636 7806 11648
rect 8012 11645 8024 11679
rect 8058 11676 8070 11679
rect 8294 11676 8300 11688
rect 8058 11648 8300 11676
rect 8058 11645 8070 11648
rect 8012 11639 8070 11645
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9180 11648 9321 11676
rect 9180 11636 9186 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9968 11685 9996 11716
rect 9953 11679 10011 11685
rect 9732 11648 9825 11676
rect 9732 11636 9738 11648
rect 9953 11645 9965 11679
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10152 11676 10180 11716
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10502 11744 10508 11756
rect 10367 11716 10508 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10612 11744 10640 11784
rect 10778 11744 10784 11756
rect 10612 11716 10784 11744
rect 10410 11676 10416 11688
rect 10152 11648 10416 11676
rect 10045 11639 10103 11645
rect 6917 11611 6975 11617
rect 6917 11608 6929 11611
rect 5736 11580 6408 11608
rect 6472 11580 6929 11608
rect 2516 11512 3004 11540
rect 3326 11500 3332 11552
rect 3384 11540 3390 11552
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3384 11512 3893 11540
rect 3384 11500 3390 11512
rect 3881 11509 3893 11512
rect 3927 11509 3939 11543
rect 3881 11503 3939 11509
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5537 11543 5595 11549
rect 4028 11512 4073 11540
rect 4028 11500 4034 11512
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 5736 11540 5764 11580
rect 5583 11512 5764 11540
rect 5813 11543 5871 11549
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 5902 11540 5908 11552
rect 5859 11512 5908 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6086 11540 6092 11552
rect 6047 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6380 11540 6408 11580
rect 6917 11577 6929 11580
rect 6963 11577 6975 11611
rect 7760 11608 7788 11636
rect 8202 11608 8208 11620
rect 7760 11580 8208 11608
rect 6917 11571 6975 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 10060 11608 10088 11639
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10612 11685 10640 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11645 10747 11679
rect 11146 11676 11152 11688
rect 11107 11648 11152 11676
rect 10689 11639 10747 11645
rect 10505 11611 10563 11617
rect 10505 11608 10517 11611
rect 9640 11580 10517 11608
rect 9640 11568 9646 11580
rect 10505 11577 10517 11580
rect 10551 11577 10563 11611
rect 10505 11571 10563 11577
rect 7282 11540 7288 11552
rect 6380 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7558 11540 7564 11552
rect 7515 11512 7564 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10704 11540 10732 11639
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 11514 11676 11520 11688
rect 11471 11648 11520 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 10962 11540 10968 11552
rect 10008 11512 10732 11540
rect 10923 11512 10968 11540
rect 10008 11500 10014 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 1104 11450 12328 11472
rect 1104 11398 4723 11450
rect 4775 11398 4787 11450
rect 4839 11398 4851 11450
rect 4903 11398 4915 11450
rect 4967 11398 8464 11450
rect 8516 11398 8528 11450
rect 8580 11398 8592 11450
rect 8644 11398 8656 11450
rect 8708 11398 12328 11450
rect 1104 11376 12328 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2280 11308 2636 11336
rect 2280 11296 2286 11308
rect 1857 11271 1915 11277
rect 1857 11268 1869 11271
rect 1412 11240 1869 11268
rect 1412 11209 1440 11240
rect 1857 11237 1869 11240
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 2608 11268 2636 11308
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3050 11336 3056 11348
rect 2832 11308 2877 11336
rect 3011 11308 3056 11336
rect 2832 11296 2838 11308
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 5626 11336 5632 11348
rect 5491 11308 5632 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6178 11336 6184 11348
rect 5828 11308 6184 11336
rect 4157 11271 4215 11277
rect 2096 11240 2544 11268
rect 2608 11240 2774 11268
rect 2096 11228 2102 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1397 11163 1455 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2130 11200 2136 11212
rect 2091 11172 2136 11200
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2516 11209 2544 11240
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11169 2375 11203
rect 2317 11163 2375 11169
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11169 2559 11203
rect 2746 11200 2774 11240
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 4246 11268 4252 11280
rect 4203 11240 4252 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2746 11172 2881 11200
rect 2501 11163 2559 11169
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 3326 11200 3332 11212
rect 3287 11172 3332 11200
rect 2869 11163 2927 11169
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1719 11104 2237 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2332 11132 2360 11163
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11169 3571 11203
rect 3878 11200 3884 11212
rect 3839 11172 3884 11200
rect 3513 11163 3571 11169
rect 2777 11135 2835 11141
rect 2332 11104 2544 11132
rect 2225 11095 2283 11101
rect 2516 11076 2544 11104
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 3421 11135 3479 11141
rect 3421 11132 3433 11135
rect 2823 11104 3433 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 3421 11101 3433 11104
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 566 11024 572 11076
rect 624 11064 630 11076
rect 842 11064 848 11076
rect 624 11036 848 11064
rect 624 11024 630 11036
rect 842 11024 848 11036
rect 900 11024 906 11076
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 3528 11064 3556 11163
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4522 11200 4528 11212
rect 4479 11172 4528 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 4154 11132 4160 11144
rect 4115 11104 4160 11132
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4724 11132 4752 11163
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 4856 11172 5089 11200
rect 4856 11160 4862 11172
rect 5077 11169 5089 11172
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5258 11200 5264 11212
rect 5215 11172 5264 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5442 11200 5448 11212
rect 5399 11172 5448 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5828 11209 5856 11308
rect 6178 11296 6184 11308
rect 6236 11336 6242 11348
rect 6236 11308 6500 11336
rect 6236 11296 6242 11308
rect 6270 11228 6276 11280
rect 6328 11277 6334 11280
rect 6328 11271 6392 11277
rect 6328 11237 6346 11271
rect 6380 11237 6392 11271
rect 6472 11268 6500 11308
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 7926 11336 7932 11348
rect 6604 11308 7932 11336
rect 6604 11296 6610 11308
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 9674 11296 9680 11348
rect 9732 11296 9738 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 10100 11308 10149 11336
rect 10100 11296 10106 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10376 11308 11100 11336
rect 10376 11296 10382 11308
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 6472 11240 7573 11268
rect 6328 11231 6392 11237
rect 7561 11237 7573 11240
rect 7607 11237 7619 11271
rect 7561 11231 7619 11237
rect 7837 11271 7895 11277
rect 7837 11237 7849 11271
rect 7883 11268 7895 11271
rect 8294 11268 8300 11280
rect 7883 11240 8300 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 6328 11228 6334 11231
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 8478 11268 8484 11280
rect 8439 11240 8484 11268
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8697 11271 8755 11277
rect 8697 11237 8709 11271
rect 8743 11268 8755 11271
rect 8938 11268 8944 11280
rect 8743 11240 8944 11268
rect 8743 11237 8755 11240
rect 8697 11231 8755 11237
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6914 11200 6920 11212
rect 6135 11172 6920 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 8110 11200 8116 11212
rect 8071 11172 8116 11200
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9692 11209 9720 11296
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 10410 11268 10416 11280
rect 9999 11240 10416 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 10560 11240 10824 11268
rect 10560 11228 10566 11240
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 9088 11172 9137 11200
rect 9088 11160 9094 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11200 9919 11203
rect 10318 11200 10324 11212
rect 9907 11172 10324 11200
rect 9907 11169 9919 11172
rect 9861 11163 9919 11169
rect 9766 11132 9772 11144
rect 4396 11104 4752 11132
rect 9727 11104 9772 11132
rect 4396 11092 4402 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9876 11076 9904 11163
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10520 11200 10548 11228
rect 10796 11209 10824 11240
rect 10419 11172 10548 11200
rect 10597 11203 10655 11209
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 2556 11036 3556 11064
rect 3973 11067 4031 11073
rect 2556 11024 2562 11036
rect 3973 11033 3985 11067
rect 4019 11033 4031 11067
rect 3973 11027 4031 11033
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 4430 11064 4436 11076
rect 4295 11036 4436 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10996 1550 11008
rect 2593 10999 2651 11005
rect 2593 10996 2605 10999
rect 1544 10968 2605 10996
rect 1544 10956 1550 10968
rect 2593 10965 2605 10968
rect 2639 10996 2651 10999
rect 3988 10996 4016 11027
rect 4430 11024 4436 11036
rect 4488 11024 4494 11076
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7515 11036 7573 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 7561 11027 7619 11033
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 9309 11067 9367 11073
rect 8251 11036 9076 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 4062 10996 4068 11008
rect 2639 10968 4068 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4525 10999 4583 11005
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 4798 10996 4804 11008
rect 4571 10968 4804 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 4948 10968 4993 10996
rect 4948 10956 4954 10968
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 5261 10999 5319 11005
rect 5261 10996 5273 10999
rect 5224 10968 5273 10996
rect 5224 10956 5230 10968
rect 5261 10965 5273 10968
rect 5307 10965 5319 10999
rect 5261 10959 5319 10965
rect 5905 10999 5963 11005
rect 5905 10965 5917 10999
rect 5951 10996 5963 10999
rect 5994 10996 6000 11008
rect 5951 10968 6000 10996
rect 5951 10965 5963 10968
rect 5905 10959 5963 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 8680 11005 8708 11036
rect 8665 10999 8723 11005
rect 8665 10965 8677 10999
rect 8711 10965 8723 10999
rect 8846 10996 8852 11008
rect 8807 10968 8852 10996
rect 8665 10959 8723 10965
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9048 10996 9076 11036
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9858 11064 9864 11076
rect 9355 11036 9864 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 10419 11064 10447 11172
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 10686 11203 10744 11209
rect 10686 11169 10698 11203
rect 10732 11169 10744 11203
rect 10686 11163 10744 11169
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 10100 11036 10447 11064
rect 10612 11064 10640 11163
rect 10704 11132 10732 11163
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11072 11209 11100 11308
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10928 11172 10977 11200
rect 10928 11160 10934 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11238 11200 11244 11212
rect 11199 11172 11244 11200
rect 11057 11163 11115 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11514 11200 11520 11212
rect 11475 11172 11520 11200
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 10704 11104 11161 11132
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 10686 11064 10692 11076
rect 10612 11036 10692 11064
rect 10100 11024 10106 11036
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 10060 10996 10088 11024
rect 9048 10968 10088 10996
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10996 10379 10999
rect 10778 10996 10784 11008
rect 10367 10968 10784 10996
rect 10367 10965 10379 10968
rect 10321 10959 10379 10965
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11330 10996 11336 11008
rect 11291 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 1104 10906 12328 10928
rect 1104 10854 2852 10906
rect 2904 10854 2916 10906
rect 2968 10854 2980 10906
rect 3032 10854 3044 10906
rect 3096 10854 6594 10906
rect 6646 10854 6658 10906
rect 6710 10854 6722 10906
rect 6774 10854 6786 10906
rect 6838 10854 10335 10906
rect 10387 10854 10399 10906
rect 10451 10854 10463 10906
rect 10515 10854 10527 10906
rect 10579 10854 12328 10906
rect 1104 10832 12328 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 1762 10792 1768 10804
rect 1443 10764 1768 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 3418 10792 3424 10804
rect 1872 10764 3424 10792
rect 1872 10656 1900 10764
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 5534 10792 5540 10804
rect 3568 10764 4936 10792
rect 5495 10764 5540 10792
rect 3568 10752 3574 10764
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 2774 10724 2780 10736
rect 2639 10696 2780 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 3786 10724 3792 10736
rect 3292 10696 3792 10724
rect 3292 10684 3298 10696
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 4908 10724 4936 10764
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5859 10764 6132 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 4908 10696 5488 10724
rect 1780 10628 1900 10656
rect 2041 10659 2099 10665
rect 1780 10597 1808 10628
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2222 10656 2228 10668
rect 2087 10628 2228 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2222 10616 2228 10628
rect 2280 10656 2286 10668
rect 2406 10656 2412 10668
rect 2280 10628 2412 10656
rect 2280 10616 2286 10628
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3384 10628 3617 10656
rect 3384 10616 3390 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 3752 10628 3797 10656
rect 3752 10616 3758 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2317 10591 2375 10597
rect 2317 10588 2329 10591
rect 1903 10560 2329 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2317 10557 2329 10560
rect 2363 10557 2375 10591
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2317 10551 2375 10557
rect 2332 10520 2360 10551
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2774 10588 2780 10600
rect 2735 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 5460 10597 5488 10696
rect 5994 10684 6000 10736
rect 6052 10684 6058 10736
rect 6104 10724 6132 10764
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6420 10764 6561 10792
rect 6420 10752 6426 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8202 10792 8208 10804
rect 7064 10764 8208 10792
rect 7064 10752 7070 10764
rect 7193 10727 7251 10733
rect 7193 10724 7205 10727
rect 6104 10696 6224 10724
rect 5644 10628 5948 10656
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 5445 10591 5503 10597
rect 4019 10560 5396 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 2958 10520 2964 10532
rect 2332 10492 2964 10520
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 3068 10520 3096 10551
rect 3326 10520 3332 10532
rect 3068 10492 3332 10520
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 3602 10520 3608 10532
rect 3436 10492 3608 10520
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2866 10452 2872 10464
rect 2827 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3234 10412 3240 10464
rect 3292 10452 3298 10464
rect 3436 10452 3464 10492
rect 3602 10480 3608 10492
rect 3660 10520 3666 10532
rect 3988 10520 4016 10551
rect 4237 10520 4243 10532
rect 3660 10492 4016 10520
rect 4198 10492 4243 10520
rect 3660 10480 3666 10492
rect 4237 10480 4243 10492
rect 4295 10480 4301 10532
rect 5368 10520 5396 10560
rect 5445 10557 5457 10591
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5644 10597 5672 10628
rect 5920 10597 5948 10628
rect 6012 10597 6040 10684
rect 6196 10656 6224 10696
rect 6656 10696 7205 10724
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 6196 10628 6285 10656
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 6656 10600 6684 10696
rect 7193 10693 7205 10696
rect 7239 10693 7251 10727
rect 7193 10687 7251 10693
rect 7300 10665 7328 10764
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8536 10764 8861 10792
rect 8536 10752 8542 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 10870 10792 10876 10804
rect 9539 10764 10876 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11296 10764 11529 10792
rect 11296 10752 11302 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 8220 10724 8248 10752
rect 9674 10724 9680 10736
rect 8220 10696 9680 10724
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 9858 10684 9864 10736
rect 9916 10684 9922 10736
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 7285 10619 7343 10625
rect 9048 10628 9781 10656
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5592 10560 5641 10588
rect 5592 10548 5598 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5727 10591 5785 10597
rect 5727 10557 5739 10591
rect 5773 10557 5785 10591
rect 5727 10551 5785 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6178 10588 6184 10600
rect 6135 10560 6184 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 5368 10492 5580 10520
rect 5552 10464 5580 10492
rect 3292 10424 3464 10452
rect 3513 10455 3571 10461
rect 3292 10412 3298 10424
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3970 10452 3976 10464
rect 3559 10424 3976 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 4672 10424 5365 10452
rect 4672 10412 4678 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 5736 10452 5764 10551
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10557 6515 10591
rect 6638 10588 6644 10600
rect 6599 10560 6644 10588
rect 6457 10551 6515 10557
rect 6472 10520 6500 10551
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6914 10588 6920 10600
rect 6875 10560 6920 10588
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7552 10591 7610 10597
rect 7552 10557 7564 10591
rect 7598 10588 7610 10591
rect 8846 10588 8852 10600
rect 7598 10560 8852 10588
rect 7598 10557 7610 10560
rect 7552 10551 7610 10557
rect 6196 10492 6500 10520
rect 6196 10464 6224 10492
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 7024 10520 7052 10551
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9048 10597 9076 10628
rect 9769 10625 9781 10628
rect 9815 10656 9827 10659
rect 9876 10656 9904 10684
rect 9815 10628 9904 10656
rect 10137 10659 10195 10665
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10183 10628 10272 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10244 10600 10272 10628
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9355 10560 9689 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9677 10557 9689 10560
rect 9723 10588 9735 10591
rect 9861 10591 9919 10597
rect 9723 10560 9812 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9784 10532 9812 10560
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 9999 10560 10088 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 8294 10520 8300 10532
rect 6604 10492 6960 10520
rect 7024 10492 8300 10520
rect 6604 10480 6610 10492
rect 5994 10452 6000 10464
rect 5736 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6178 10412 6184 10464
rect 6236 10412 6242 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6362 10452 6368 10464
rect 6319 10424 6368 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6730 10452 6736 10464
rect 6691 10424 6736 10452
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 6932 10452 6960 10492
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 9582 10520 9588 10532
rect 8588 10492 9588 10520
rect 8588 10452 8616 10492
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 9766 10480 9772 10532
rect 9824 10480 9830 10532
rect 6932 10424 8616 10452
rect 8665 10455 8723 10461
rect 8665 10421 8677 10455
rect 8711 10452 8723 10455
rect 9030 10452 9036 10464
rect 8711 10424 9036 10452
rect 8711 10421 8723 10424
rect 8665 10415 8723 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9217 10455 9275 10461
rect 9217 10421 9229 10455
rect 9263 10452 9275 10455
rect 9674 10452 9680 10464
rect 9263 10424 9680 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 9674 10412 9680 10424
rect 9732 10452 9738 10464
rect 9876 10452 9904 10551
rect 9732 10424 9904 10452
rect 10060 10452 10088 10560
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10336 10560 10907 10588
rect 10336 10452 10364 10560
rect 10404 10523 10462 10529
rect 10404 10489 10416 10523
rect 10450 10520 10462 10523
rect 10778 10520 10784 10532
rect 10450 10492 10784 10520
rect 10450 10489 10462 10492
rect 10404 10483 10462 10489
rect 10778 10480 10784 10492
rect 10836 10480 10842 10532
rect 10879 10520 10907 10560
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11204 10560 11897 10588
rect 11204 10548 11210 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 11238 10520 11244 10532
rect 10879 10492 11244 10520
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 10060 10424 10364 10452
rect 9732 10412 9738 10424
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 10560 10424 11713 10452
rect 10560 10412 10566 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 1104 10362 12328 10384
rect 1104 10310 4723 10362
rect 4775 10310 4787 10362
rect 4839 10310 4851 10362
rect 4903 10310 4915 10362
rect 4967 10310 8464 10362
rect 8516 10310 8528 10362
rect 8580 10310 8592 10362
rect 8644 10310 8656 10362
rect 8708 10310 12328 10362
rect 1104 10288 12328 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 2924 10220 3648 10248
rect 2924 10208 2930 10220
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 2010 10183 2068 10189
rect 2010 10180 2022 10183
rect 1719 10152 2022 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 2010 10149 2022 10152
rect 2056 10149 2068 10183
rect 2010 10143 2068 10149
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 3200 10152 3556 10180
rect 3200 10140 3206 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 2406 10112 2412 10124
rect 1544 10084 1589 10112
rect 1688 10084 2412 10112
rect 1544 10072 1550 10084
rect 1688 10053 1716 10084
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 3418 10112 3424 10124
rect 3379 10084 3424 10112
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 3528 10121 3556 10152
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10081 3571 10115
rect 3620 10112 3648 10220
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4212 10220 4721 10248
rect 4212 10208 4218 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9766 10248 9772 10260
rect 9539 10220 9772 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9766 10208 9772 10220
rect 9824 10248 9830 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9824 10220 9965 10248
rect 9824 10208 9830 10220
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 9953 10211 10011 10217
rect 10413 10251 10471 10257
rect 10413 10217 10425 10251
rect 10459 10248 10471 10251
rect 10686 10248 10692 10260
rect 10459 10220 10692 10248
rect 10459 10217 10471 10220
rect 10413 10211 10471 10217
rect 4890 10180 4896 10192
rect 4172 10152 4896 10180
rect 4172 10124 4200 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 5810 10189 5816 10192
rect 5804 10143 5816 10189
rect 5868 10180 5874 10192
rect 5868 10152 5904 10180
rect 5810 10140 5816 10143
rect 5868 10140 5874 10152
rect 7834 10140 7840 10192
rect 7892 10180 7898 10192
rect 9858 10180 9864 10192
rect 7892 10152 7972 10180
rect 7892 10140 7898 10152
rect 3878 10112 3884 10124
rect 3620 10084 3884 10112
rect 3513 10075 3571 10081
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 4080 10044 4108 10075
rect 4154 10072 4160 10124
rect 4212 10072 4218 10124
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10112 4399 10115
rect 4430 10112 4436 10124
rect 4387 10084 4436 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 4614 10112 4620 10124
rect 4575 10084 4620 10112
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4764 10084 4813 10112
rect 4764 10072 4770 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5353 10115 5411 10121
rect 5132 10084 5177 10112
rect 5132 10072 5138 10084
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5353 10075 5411 10081
rect 1820 10016 1865 10044
rect 2884 10016 4108 10044
rect 1820 10004 1826 10016
rect 1486 9868 1492 9920
rect 1544 9908 1550 9920
rect 2884 9908 2912 10016
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5368 10044 5396 10075
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7098 10112 7104 10124
rect 7059 10084 7104 10112
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 7944 10121 7972 10152
rect 8772 10152 9168 10180
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7745 10115 7803 10121
rect 7515 10084 7696 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 4948 10016 5396 10044
rect 7377 10047 7435 10053
rect 4948 10004 4954 10016
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7423 10016 7604 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3145 9979 3203 9985
rect 3145 9976 3157 9979
rect 3016 9948 3157 9976
rect 3016 9936 3022 9948
rect 3145 9945 3157 9948
rect 3191 9945 3203 9979
rect 3145 9939 3203 9945
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4246 9976 4252 9988
rect 3927 9948 4252 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 1544 9880 2912 9908
rect 3237 9911 3295 9917
rect 1544 9868 1550 9880
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3510 9908 3516 9920
rect 3283 9880 3516 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 3970 9908 3976 9920
rect 3651 9880 3976 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9908 4215 9911
rect 4706 9908 4712 9920
rect 4203 9880 4712 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 4893 9911 4951 9917
rect 4893 9877 4905 9911
rect 4939 9908 4951 9911
rect 5074 9908 5080 9920
rect 4939 9880 5080 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5534 9908 5540 9920
rect 5215 9880 5540 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7190 9908 7196 9920
rect 7151 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7374 9908 7380 9920
rect 7331 9880 7380 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7576 9908 7604 10016
rect 7668 9976 7696 10084
rect 7745 10081 7757 10115
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8047 10115 8105 10121
rect 8047 10081 8059 10115
rect 8093 10112 8105 10115
rect 8202 10112 8208 10124
rect 8093 10084 8208 10112
rect 8093 10081 8105 10084
rect 8047 10075 8105 10081
rect 7760 10044 7788 10075
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8772 10121 8800 10152
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10081 8815 10115
rect 8938 10112 8944 10124
rect 8899 10084 8944 10112
rect 8757 10075 8815 10081
rect 8386 10044 8392 10056
rect 7760 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8496 10044 8524 10075
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9140 10121 9168 10152
rect 9508 10152 9864 10180
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9398 10112 9404 10124
rect 9171 10084 9404 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 8846 10044 8852 10056
rect 8496 10016 8852 10044
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8662 9976 8668 9988
rect 7668 9948 8668 9976
rect 8662 9936 8668 9948
rect 8720 9936 8726 9988
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7576 9880 7849 9908
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9122 9908 9128 9920
rect 8803 9880 9128 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9508 9917 9536 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9968 10112 9996 10211
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10318 10180 10324 10192
rect 10100 10152 10324 10180
rect 10100 10140 10106 10152
rect 10318 10140 10324 10152
rect 10376 10180 10382 10192
rect 11330 10180 11336 10192
rect 10376 10152 11336 10180
rect 10376 10140 10382 10152
rect 10612 10121 10640 10152
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 10870 10121 10876 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 9968 10084 10241 10112
rect 9769 10075 9827 10081
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 10864 10075 10876 10121
rect 10928 10112 10934 10124
rect 10928 10084 10964 10112
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9877 9551 9911
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9784 9908 9812 10075
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10428 10044 10456 10075
rect 10870 10072 10876 10075
rect 10928 10072 10934 10084
rect 9916 10016 10456 10044
rect 9916 10004 9922 10016
rect 10244 9988 10272 10016
rect 10226 9936 10232 9988
rect 10284 9936 10290 9988
rect 9950 9908 9956 9920
rect 9784 9880 9956 9908
rect 9950 9868 9956 9880
rect 10008 9908 10014 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 10008 9880 11989 9908
rect 10008 9868 10014 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 1104 9818 12328 9840
rect 1104 9766 2852 9818
rect 2904 9766 2916 9818
rect 2968 9766 2980 9818
rect 3032 9766 3044 9818
rect 3096 9766 6594 9818
rect 6646 9766 6658 9818
rect 6710 9766 6722 9818
rect 6774 9766 6786 9818
rect 6838 9766 10335 9818
rect 10387 9766 10399 9818
rect 10451 9766 10463 9818
rect 10515 9766 10527 9818
rect 10579 9766 12328 9818
rect 1104 9744 12328 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 3237 9707 3295 9713
rect 1452 9676 2912 9704
rect 1452 9664 1458 9676
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9636 2007 9639
rect 2774 9636 2780 9648
rect 1995 9608 2780 9636
rect 1995 9605 2007 9608
rect 1949 9599 2007 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2884 9645 2912 9676
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3283 9676 3556 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9605 2927 9639
rect 3418 9636 3424 9648
rect 3379 9608 3424 9636
rect 2869 9599 2927 9605
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 3528 9636 3556 9676
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 4433 9707 4491 9713
rect 4120 9676 4384 9704
rect 4120 9664 4126 9676
rect 4356 9645 4384 9676
rect 4433 9673 4445 9707
rect 4479 9704 4491 9707
rect 4706 9704 4712 9716
rect 4479 9676 4712 9704
rect 4479 9673 4491 9676
rect 4433 9667 4491 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4982 9664 4988 9716
rect 5040 9704 5046 9716
rect 5721 9707 5779 9713
rect 5040 9676 5672 9704
rect 5040 9664 5046 9676
rect 4341 9639 4399 9645
rect 3528 9608 4292 9636
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 1084 9540 1900 9568
rect 1084 9528 1090 9540
rect 1872 9509 1900 9540
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2280 9540 2513 9568
rect 2280 9528 2286 9540
rect 2501 9537 2513 9540
rect 2547 9568 2559 9571
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 2547 9540 3985 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 845 9503 903 9509
rect 845 9469 857 9503
rect 891 9500 903 9503
rect 1581 9503 1639 9509
rect 1581 9500 1593 9503
rect 891 9472 1593 9500
rect 891 9469 903 9472
rect 845 9463 903 9469
rect 1581 9469 1593 9472
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2682 9500 2688 9512
rect 2363 9472 2688 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3145 9503 3203 9509
rect 2832 9472 2877 9500
rect 2832 9460 2838 9472
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3418 9500 3424 9512
rect 3191 9472 3424 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 4264 9509 4292 9608
rect 4341 9605 4353 9639
rect 4387 9605 4399 9639
rect 4341 9599 4399 9605
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9605 5411 9639
rect 5644 9636 5672 9676
rect 5721 9673 5733 9707
rect 5767 9704 5779 9707
rect 5810 9704 5816 9716
rect 5767 9676 5816 9704
rect 5767 9673 5779 9676
rect 5721 9667 5779 9673
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6454 9704 6460 9716
rect 5920 9676 6460 9704
rect 5920 9636 5948 9676
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9704 6975 9707
rect 7098 9704 7104 9716
rect 6963 9676 7104 9704
rect 6963 9673 6975 9676
rect 6917 9667 6975 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 8938 9704 8944 9716
rect 8803 9676 8944 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10284 9676 10609 9704
rect 10284 9664 10290 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 10597 9667 10655 9673
rect 10781 9707 10839 9713
rect 10781 9673 10793 9707
rect 10827 9704 10839 9707
rect 10870 9704 10876 9716
rect 10827 9676 10876 9704
rect 10827 9673 10839 9676
rect 10781 9667 10839 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 5644 9608 5948 9636
rect 5353 9599 5411 9605
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9568 4583 9571
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4571 9540 4813 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 5368 9568 5396 9599
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 6420 9608 7144 9636
rect 6420 9596 6426 9608
rect 6914 9568 6920 9580
rect 5368 9540 5856 9568
rect 4801 9531 4859 9537
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4614 9460 4620 9512
rect 4672 9460 4678 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 3789 9435 3847 9441
rect 3789 9432 3801 9435
rect 1688 9404 3801 9432
rect 1688 9373 1716 9404
rect 3789 9401 3801 9404
rect 3835 9401 3847 9435
rect 3789 9395 3847 9401
rect 3881 9435 3939 9441
rect 3881 9401 3893 9435
rect 3927 9432 3939 9435
rect 4632 9432 4660 9460
rect 3927 9404 4660 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 753 9367 811 9373
rect 753 9333 765 9367
rect 799 9364 811 9367
rect 1397 9367 1455 9373
rect 1397 9364 1409 9367
rect 799 9336 1409 9364
rect 799 9333 811 9336
rect 753 9327 811 9333
rect 1397 9333 1409 9336
rect 1443 9333 1455 9367
rect 1397 9327 1455 9333
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9333 1731 9367
rect 1673 9327 1731 9333
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 2774 9364 2780 9376
rect 2455 9336 2780 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4724 9364 4752 9463
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 4908 9432 4936 9463
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 5132 9472 5181 9500
rect 5132 9460 5138 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5350 9500 5356 9512
rect 5307 9472 5356 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5828 9509 5856 9540
rect 6012 9540 6920 9568
rect 6012 9509 6040 9540
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7116 9568 7144 9608
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8444 9608 8493 9636
rect 8444 9596 8450 9608
rect 8481 9605 8493 9608
rect 8527 9636 8539 9639
rect 9214 9636 9220 9648
rect 8527 9608 9220 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 9950 9568 9956 9580
rect 7116 9540 7236 9568
rect 5629 9503 5687 9509
rect 5500 9472 5545 9500
rect 5500 9460 5506 9472
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 5534 9432 5540 9444
rect 4856 9404 5540 9432
rect 4856 9392 4862 9404
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 5644 9432 5672 9463
rect 6178 9460 6184 9512
rect 6236 9509 6242 9512
rect 6236 9500 6247 9509
rect 6236 9472 6329 9500
rect 6236 9463 6247 9472
rect 6236 9460 6242 9463
rect 6089 9435 6147 9441
rect 6089 9432 6101 9435
rect 5644 9404 6101 9432
rect 6089 9401 6101 9404
rect 6135 9401 6147 9435
rect 6288 9432 6316 9472
rect 6362 9460 6368 9512
rect 6420 9500 6426 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 6420 9472 6469 9500
rect 6420 9460 6426 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6696 9472 6837 9500
rect 6696 9460 6702 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 7098 9500 7104 9512
rect 7059 9472 7104 9500
rect 6825 9463 6883 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7208 9500 7236 9540
rect 8864 9540 9956 9568
rect 7374 9509 7380 9512
rect 7208 9472 7328 9500
rect 7190 9432 7196 9444
rect 6288 9404 7196 9432
rect 6089 9395 6147 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7300 9432 7328 9472
rect 7368 9463 7380 9509
rect 7432 9500 7438 9512
rect 8864 9509 8892 9540
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 8849 9503 8907 9509
rect 7432 9472 7468 9500
rect 7374 9460 7380 9463
rect 7432 9460 7438 9472
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 8849 9463 8907 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9723 9472 10180 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 10152 9444 10180 9472
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10836 9472 10885 9500
rect 10836 9460 10842 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 11514 9500 11520 9512
rect 11475 9472 11520 9500
rect 10873 9463 10931 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 12066 9500 12072 9512
rect 11931 9472 12072 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 7300 9404 9904 9432
rect 4028 9336 4752 9364
rect 4985 9367 5043 9373
rect 4028 9324 4034 9336
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 7650 9364 7656 9376
rect 5031 9336 7656 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 9674 9364 9680 9376
rect 9456 9336 9680 9364
rect 9456 9324 9462 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9876 9364 9904 9404
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10134 9432 10140 9444
rect 10008 9404 10053 9432
rect 10095 9404 10140 9432
rect 10008 9392 10014 9404
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 10686 9441 10692 9444
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9432 10379 9435
rect 10413 9435 10471 9441
rect 10413 9432 10425 9435
rect 10367 9404 10425 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 10413 9401 10425 9404
rect 10459 9401 10471 9435
rect 10413 9395 10471 9401
rect 10629 9435 10692 9441
rect 10629 9401 10641 9435
rect 10675 9401 10692 9435
rect 10629 9395 10692 9401
rect 10686 9392 10692 9395
rect 10744 9392 10750 9444
rect 10870 9364 10876 9376
rect 9876 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 1104 9274 12328 9296
rect 1104 9222 4723 9274
rect 4775 9222 4787 9274
rect 4839 9222 4851 9274
rect 4903 9222 4915 9274
rect 4967 9222 8464 9274
rect 8516 9222 8528 9274
rect 8580 9222 8592 9274
rect 8644 9222 8656 9274
rect 8708 9222 12328 9274
rect 1104 9200 12328 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3605 9163 3663 9169
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4062 9160 4068 9172
rect 3651 9132 4068 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 6144 9132 6561 9160
rect 6144 9120 6150 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 6914 9160 6920 9172
rect 6687 9132 6920 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 8352 9132 8401 9160
rect 8352 9120 8358 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 1762 9092 1768 9104
rect 1412 9064 1768 9092
rect 1412 9033 1440 9064
rect 1762 9052 1768 9064
rect 1820 9052 1826 9104
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 3234 9092 3240 9104
rect 2556 9064 3240 9092
rect 2556 9052 2562 9064
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 3496 9095 3554 9101
rect 3496 9061 3508 9095
rect 3542 9092 3554 9095
rect 3970 9092 3976 9104
rect 3542 9064 3976 9092
rect 3542 9061 3554 9064
rect 3496 9055 3554 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4148 9095 4206 9101
rect 4148 9061 4160 9095
rect 4194 9092 4206 9095
rect 4614 9092 4620 9104
rect 4194 9064 4620 9092
rect 4194 9061 4206 9064
rect 4148 9055 4206 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 4798 9052 4804 9104
rect 4856 9092 4862 9104
rect 5813 9095 5871 9101
rect 5813 9092 5825 9095
rect 4856 9064 5825 9092
rect 4856 9052 4862 9064
rect 5813 9061 5825 9064
rect 5859 9061 5871 9095
rect 5813 9055 5871 9061
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 9140 9092 9168 9123
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 9585 9163 9643 9169
rect 9585 9160 9597 9163
rect 9456 9132 9597 9160
rect 9456 9120 9462 9132
rect 9585 9129 9597 9132
rect 9631 9129 9643 9163
rect 9585 9123 9643 9129
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 6328 9064 7411 9092
rect 9140 9064 9965 9092
rect 6328 9052 6334 9064
rect 1670 9033 1676 9036
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1664 8987 1676 9033
rect 1728 9024 1734 9036
rect 1728 8996 1764 9024
rect 1670 8984 1676 8987
rect 1728 8984 1734 8996
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2280 8996 3065 9024
rect 2280 8984 2286 8996
rect 3053 8993 3065 8996
rect 3099 8993 3111 9027
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 3053 8987 3111 8993
rect 3140 8996 3341 9024
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 3140 8956 3168 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 3329 8987 3387 8993
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 4764 8996 5733 9024
rect 4764 8984 4770 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7190 9033 7196 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6972 8996 7021 9024
rect 6972 8984 6978 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7184 9024 7196 9033
rect 7151 8996 7196 9024
rect 7009 8987 7067 8993
rect 7184 8987 7196 8996
rect 7190 8984 7196 8987
rect 7248 8984 7254 9036
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 2464 8928 3168 8956
rect 2464 8916 2470 8928
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3881 8959 3939 8965
rect 3881 8956 3893 8959
rect 3292 8928 3893 8956
rect 3292 8916 3298 8928
rect 3881 8925 3893 8928
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2556 8792 2881 8820
rect 2556 8780 2562 8792
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3326 8820 3332 8832
rect 3191 8792 3332 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3896 8820 3924 8919
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5132 8928 6009 8956
rect 5132 8916 5138 8928
rect 5997 8925 6009 8928
rect 6043 8956 6055 8959
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6043 8928 6837 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 6638 8888 6644 8900
rect 5399 8860 6644 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 6638 8848 6644 8860
rect 6696 8848 6702 8900
rect 4062 8820 4068 8832
rect 3896 8792 4068 8820
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 4856 8792 5273 8820
rect 4856 8780 4862 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 6270 8820 6276 8832
rect 6227 8792 6276 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6840 8820 6868 8919
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 6972 8860 7113 8888
rect 6972 8848 6978 8860
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7300 8888 7328 8987
rect 7248 8860 7328 8888
rect 7383 8888 7411 9064
rect 9953 9061 9965 9064
rect 9999 9092 10011 9095
rect 10321 9095 10379 9101
rect 9999 9064 10272 9092
rect 9999 9061 10011 9064
rect 9953 9055 10011 9061
rect 7558 9024 7564 9036
rect 7519 8996 7564 9024
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8662 9024 8668 9036
rect 8623 8996 8668 9024
rect 8481 8987 8539 8993
rect 8496 8956 8524 8987
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 8938 8984 8944 9036
rect 8996 9024 9002 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8996 8996 9505 9024
rect 8996 8984 9002 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 10134 9024 10140 9036
rect 9493 8987 9551 8993
rect 9600 8996 10140 9024
rect 8849 8959 8907 8965
rect 8849 8956 8861 8959
rect 8496 8928 8861 8956
rect 8849 8925 8861 8928
rect 8895 8956 8907 8959
rect 9214 8956 9220 8968
rect 8895 8928 9220 8956
rect 8895 8925 8907 8928
rect 8849 8919 8907 8925
rect 9214 8916 9220 8928
rect 9272 8956 9278 8968
rect 9600 8956 9628 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10244 9024 10272 9064
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 10413 9095 10471 9101
rect 10413 9092 10425 9095
rect 10367 9064 10425 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 10413 9061 10425 9064
rect 10459 9061 10471 9095
rect 10413 9055 10471 9061
rect 10629 9095 10687 9101
rect 10629 9061 10641 9095
rect 10675 9092 10687 9095
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 10675 9064 10977 9092
rect 10675 9061 10687 9064
rect 10629 9055 10687 9061
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 10965 9055 11023 9061
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10244 8996 10885 9024
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11146 9024 11152 9036
rect 11103 8996 11152 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 9272 8928 9628 8956
rect 9769 8959 9827 8965
rect 9272 8916 9278 8928
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 11238 8956 11244 8968
rect 9815 8928 11244 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 9950 8888 9956 8900
rect 7383 8860 9956 8888
rect 7248 8848 7254 8860
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 8662 8820 8668 8832
rect 6840 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8820 8726 8832
rect 9030 8820 9036 8832
rect 8720 8792 9036 8820
rect 8720 8780 8726 8792
rect 9030 8780 9036 8792
rect 9088 8820 9094 8832
rect 10060 8820 10088 8928
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 10192 8860 11621 8888
rect 10192 8848 10198 8860
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 9088 8792 10088 8820
rect 9088 8780 9094 8792
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10284 8792 10609 8820
rect 10284 8780 10290 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 10597 8783 10655 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11330 8820 11336 8832
rect 11291 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11756 8792 11897 8820
rect 11756 8780 11762 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 11885 8783 11943 8789
rect 1104 8730 12328 8752
rect 1104 8678 2852 8730
rect 2904 8678 2916 8730
rect 2968 8678 2980 8730
rect 3032 8678 3044 8730
rect 3096 8678 6594 8730
rect 6646 8678 6658 8730
rect 6710 8678 6722 8730
rect 6774 8678 6786 8730
rect 6838 8678 10335 8730
rect 10387 8678 10399 8730
rect 10451 8678 10463 8730
rect 10515 8678 10527 8730
rect 10579 8678 12328 8730
rect 1104 8656 12328 8678
rect 1394 8616 1400 8628
rect 1355 8588 1400 8616
rect 1394 8576 1400 8588
rect 1452 8576 1458 8628
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1857 8619 1915 8625
rect 1857 8616 1869 8619
rect 1728 8588 1869 8616
rect 1728 8576 1734 8588
rect 1857 8585 1869 8588
rect 1903 8585 1915 8619
rect 1857 8579 1915 8585
rect 2240 8588 2912 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 2240 8548 2268 8588
rect 2884 8560 2912 8588
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 3292 8588 4261 8616
rect 3292 8576 3298 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7190 8616 7196 8628
rect 7064 8588 7196 8616
rect 7064 8576 7070 8588
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 8386 8616 8392 8628
rect 8347 8588 8392 8616
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 8938 8616 8944 8628
rect 8899 8588 8944 8616
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9766 8616 9772 8628
rect 9447 8588 9772 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9766 8576 9772 8588
rect 9824 8616 9830 8628
rect 9824 8588 10824 8616
rect 9824 8576 9830 8588
rect 1811 8520 2268 8548
rect 2516 8520 2774 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 1995 8452 2421 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2409 8449 2421 8452
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 842 8372 848 8424
rect 900 8412 906 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 900 8384 1593 8412
rect 900 8372 906 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 1688 8344 1716 8375
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 2038 8412 2044 8424
rect 1820 8384 2044 8412
rect 1820 8372 1826 8384
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2516 8421 2544 8520
rect 2746 8480 2774 8520
rect 2866 8508 2872 8560
rect 2924 8508 2930 8560
rect 5350 8548 5356 8560
rect 4816 8520 5356 8548
rect 2746 8452 3004 8480
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 2869 8415 2927 8421
rect 2639 8384 2820 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2130 8344 2136 8356
rect 1688 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 2332 8344 2360 8375
rect 2682 8344 2688 8356
rect 2332 8316 2688 8344
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 2038 8276 2044 8288
rect 1999 8248 2044 8276
rect 2038 8236 2044 8248
rect 2096 8236 2102 8288
rect 2792 8276 2820 8384
rect 2869 8381 2881 8415
rect 2915 8381 2927 8415
rect 2976 8412 3004 8452
rect 3418 8412 3424 8424
rect 2976 8384 3424 8412
rect 2869 8375 2927 8381
rect 2884 8344 2912 8375
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4816 8412 4844 8520
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6178 8548 6184 8560
rect 6135 8520 6184 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 6178 8508 6184 8520
rect 6236 8508 6242 8560
rect 10796 8548 10824 8588
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11238 8616 11244 8628
rect 11112 8588 11244 8616
rect 11112 8576 11118 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11146 8548 11152 8560
rect 10796 8520 11152 8548
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 4982 8480 4988 8492
rect 4943 8452 4988 8480
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5629 8483 5687 8489
rect 5132 8452 5177 8480
rect 5132 8440 5138 8452
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 6454 8480 6460 8492
rect 5675 8452 6460 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10778 8480 10784 8492
rect 10183 8452 10784 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4816 8384 4905 8412
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 5350 8412 5356 8424
rect 5311 8384 5356 8412
rect 4893 8375 4951 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5534 8412 5540 8424
rect 5491 8384 5540 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 6638 8412 6644 8424
rect 5592 8384 6500 8412
rect 6599 8384 6644 8412
rect 5592 8372 5598 8384
rect 2958 8344 2964 8356
rect 2884 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3050 8304 3056 8356
rect 3108 8353 3114 8356
rect 3108 8347 3172 8353
rect 3108 8313 3126 8347
rect 3160 8313 3172 8347
rect 3108 8307 3172 8313
rect 3108 8304 3114 8307
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 4028 8316 5917 8344
rect 4028 8304 4034 8316
rect 5460 8288 5488 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 6472 8344 6500 8384
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7098 8412 7104 8424
rect 7055 8384 7104 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 6748 8344 6776 8375
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8481 8415 8539 8421
rect 8481 8412 8493 8415
rect 7800 8384 8493 8412
rect 7800 8372 7806 8384
rect 8481 8381 8493 8384
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 9214 8412 9220 8424
rect 9175 8384 9220 8412
rect 8849 8375 8907 8381
rect 6822 8344 6828 8356
rect 6472 8316 6828 8344
rect 5905 8307 5963 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 6917 8347 6975 8353
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 7254 8347 7312 8353
rect 7254 8344 7266 8347
rect 6963 8316 7266 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 7254 8313 7266 8316
rect 7300 8313 7312 8347
rect 7254 8307 7312 8313
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8864 8344 8892 8375
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9766 8412 9772 8424
rect 9727 8384 9772 8412
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10060 8412 10088 8440
rect 10226 8412 10232 8424
rect 9907 8384 10232 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 11882 8412 11888 8424
rect 11843 8384 11888 8412
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 8352 8316 8892 8344
rect 8352 8304 8358 8316
rect 3878 8276 3884 8288
rect 2792 8248 3884 8276
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 4488 8248 4537 8276
rect 4488 8236 4494 8248
rect 4525 8245 4537 8248
rect 4571 8245 4583 8279
rect 4525 8239 4583 8245
rect 5442 8236 5448 8288
rect 5500 8236 5506 8288
rect 5626 8276 5632 8288
rect 5587 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 1104 8186 12328 8208
rect 1104 8134 4723 8186
rect 4775 8134 4787 8186
rect 4839 8134 4851 8186
rect 4903 8134 4915 8186
rect 4967 8134 8464 8186
rect 8516 8134 8528 8186
rect 8580 8134 8592 8186
rect 8644 8134 8656 8186
rect 8708 8134 12328 8186
rect 1104 8112 12328 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 2188 8044 2513 8072
rect 2188 8032 2194 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 3050 8072 3056 8084
rect 3011 8044 3056 8072
rect 2501 8035 2559 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5350 8072 5356 8084
rect 4571 8044 5356 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6638 8072 6644 8084
rect 6411 8044 6644 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 7340 8044 8401 8072
rect 7340 8032 7346 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8849 8075 8907 8081
rect 8849 8041 8861 8075
rect 8895 8072 8907 8075
rect 9950 8072 9956 8084
rect 8895 8044 9956 8072
rect 8895 8041 8907 8044
rect 8849 8035 8907 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 2041 8007 2099 8013
rect 2041 7973 2053 8007
rect 2087 8004 2099 8007
rect 3970 8004 3976 8016
rect 2087 7976 3280 8004
rect 3931 7976 3976 8004
rect 2087 7973 2099 7976
rect 2041 7967 2099 7973
rect 3252 7948 3280 7976
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 4976 8007 5034 8013
rect 4080 7976 4568 8004
rect 2409 7939 2467 7945
rect 2409 7905 2421 7939
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 2130 7868 2136 7880
rect 1820 7840 2136 7868
rect 1820 7828 1826 7840
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 382 7760 388 7812
rect 440 7800 446 7812
rect 1302 7800 1308 7812
rect 440 7772 1308 7800
rect 440 7760 446 7772
rect 1302 7760 1308 7772
rect 1360 7760 1366 7812
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2424 7800 2452 7899
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2740 7908 2789 7936
rect 2740 7896 2746 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3234 7936 3240 7948
rect 2924 7908 2969 7936
rect 3195 7908 3240 7936
rect 2924 7896 2930 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3418 7936 3424 7948
rect 3379 7908 3424 7936
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 3878 7936 3884 7948
rect 3559 7908 3884 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4080 7936 4108 7976
rect 4430 7936 4436 7948
rect 3988 7908 4108 7936
rect 4391 7908 4436 7936
rect 1627 7772 2452 7800
rect 2884 7800 2912 7896
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3099 7840 3341 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3142 7800 3148 7812
rect 2884 7772 3148 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 3988 7800 4016 7908
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4540 7936 4568 7976
rect 4976 7973 4988 8007
rect 5022 8004 5034 8007
rect 5626 8004 5632 8016
rect 5022 7976 5632 8004
rect 5022 7973 5034 7976
rect 4976 7967 5034 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 6178 8004 6184 8016
rect 6091 7976 6184 8004
rect 6178 7964 6184 7976
rect 6236 8004 6242 8016
rect 6236 7976 6776 8004
rect 6236 7964 6242 7976
rect 5994 7936 6000 7948
rect 4540 7908 6000 7936
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6748 7945 6776 7976
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 9398 8004 9404 8016
rect 6880 7976 7052 8004
rect 6880 7964 6886 7976
rect 7024 7945 7052 7976
rect 7668 7976 9404 8004
rect 7668 7945 7696 7976
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 10042 8004 10048 8016
rect 9508 7976 10048 8004
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6380 7908 6561 7936
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4120 7840 4721 7868
rect 4120 7828 4126 7840
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 6380 7868 6408 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8849 7939 8907 7945
rect 8849 7936 8861 7939
rect 7975 7908 8861 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8849 7905 8861 7908
rect 8895 7905 8907 7939
rect 9122 7936 9128 7948
rect 9083 7908 9128 7936
rect 8849 7899 8907 7905
rect 4709 7831 4767 7837
rect 6104 7840 6408 7868
rect 3292 7772 4016 7800
rect 3292 7760 3298 7772
rect 3160 7732 3188 7760
rect 6104 7744 6132 7840
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6512 7840 6653 7868
rect 6512 7828 6518 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6270 7760 6276 7812
rect 6328 7800 6334 7812
rect 6546 7800 6552 7812
rect 6328 7772 6552 7800
rect 6328 7760 6334 7772
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 6932 7800 6960 7899
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9508 7945 9536 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10588 8007 10646 8013
rect 10588 7973 10600 8007
rect 10634 8004 10646 8007
rect 10686 8004 10692 8016
rect 10634 7976 10692 8004
rect 10634 7973 10646 7976
rect 10588 7967 10646 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 11054 7936 11060 7948
rect 9723 7908 11060 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 8352 7840 8493 7868
rect 8352 7828 8358 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9030 7868 9036 7880
rect 8720 7840 9036 7868
rect 8720 7828 8726 7840
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9447 7840 9597 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10008 7840 10241 7868
rect 10008 7828 10014 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10376 7840 10421 7868
rect 10376 7828 10382 7840
rect 8846 7800 8852 7812
rect 6932 7772 8852 7800
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 9217 7803 9275 7809
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 9674 7800 9680 7812
rect 9263 7772 9680 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3160 7704 4077 7732
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 4065 7695 4123 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 6236 7704 6281 7732
rect 6236 7692 6242 7704
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 8021 7735 8079 7741
rect 7156 7704 7201 7732
rect 7156 7692 7162 7704
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 9030 7732 9036 7744
rect 8067 7704 9036 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9953 7735 10011 7741
rect 9364 7704 9409 7732
rect 9364 7692 9370 7704
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10226 7732 10232 7744
rect 9999 7704 10232 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11020 7704 11713 7732
rect 11020 7692 11026 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11974 7732 11980 7744
rect 11935 7704 11980 7732
rect 11701 7695 11759 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 1104 7642 12328 7664
rect 1104 7590 2852 7642
rect 2904 7590 2916 7642
rect 2968 7590 2980 7642
rect 3032 7590 3044 7642
rect 3096 7590 6594 7642
rect 6646 7590 6658 7642
rect 6710 7590 6722 7642
rect 6774 7590 6786 7642
rect 6838 7590 10335 7642
rect 10387 7590 10399 7642
rect 10451 7590 10463 7642
rect 10515 7590 10527 7642
rect 10579 7590 12328 7642
rect 1104 7568 12328 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2314 7528 2320 7540
rect 2087 7500 2320 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2682 7528 2688 7540
rect 2643 7500 2688 7528
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 3234 7528 3240 7540
rect 2976 7500 3240 7528
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1946 7460 1952 7472
rect 1544 7432 1952 7460
rect 1544 7420 1550 7432
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 1486 7324 1492 7336
rect 1447 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7284 1550 7336
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2406 7324 2412 7336
rect 2271 7296 2412 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 2866 7324 2872 7336
rect 2639 7296 2872 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 2516 7256 2544 7287
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 2774 7256 2780 7268
rect 2516 7228 2780 7256
rect 2774 7216 2780 7228
rect 2832 7216 2838 7268
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2976 7188 3004 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3476 7500 3985 7528
rect 3476 7488 3482 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 5074 7528 5080 7540
rect 3973 7491 4031 7497
rect 4724 7500 5080 7528
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3513 7463 3571 7469
rect 3513 7460 3525 7463
rect 3200 7432 3525 7460
rect 3200 7420 3206 7432
rect 3513 7429 3525 7432
rect 3559 7429 3571 7463
rect 3513 7423 3571 7429
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7429 3663 7463
rect 3605 7423 3663 7429
rect 3050 7284 3056 7336
rect 3108 7284 3114 7336
rect 3234 7324 3240 7336
rect 3195 7296 3240 7324
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3620 7324 3648 7423
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3970 7392 3976 7404
rect 3743 7364 3976 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4724 7392 4752 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5534 7528 5540 7540
rect 5215 7500 5540 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5534 7488 5540 7500
rect 5592 7528 5598 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 5592 7500 6193 7528
rect 5592 7488 5598 7500
rect 6181 7497 6193 7500
rect 6227 7528 6239 7531
rect 6454 7528 6460 7540
rect 6227 7500 6460 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 7248 7500 8401 7528
rect 7248 7488 7254 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 8389 7491 8447 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10413 7531 10471 7537
rect 10413 7497 10425 7531
rect 10459 7528 10471 7531
rect 10686 7528 10692 7540
rect 10459 7500 10692 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 6822 7460 6828 7472
rect 4264 7364 4752 7392
rect 4816 7432 6828 7460
rect 4154 7324 4160 7336
rect 3620 7296 4160 7324
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4264 7333 4292 7364
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4706 7324 4712 7336
rect 4571 7296 4712 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4816 7333 4844 7432
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 7926 7460 7932 7472
rect 7887 7432 7932 7460
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10321 7463 10379 7469
rect 10321 7460 10333 7463
rect 9732 7432 10333 7460
rect 9732 7420 9738 7432
rect 10321 7429 10333 7432
rect 10367 7429 10379 7463
rect 10321 7423 10379 7429
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5399 7364 5825 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6178 7392 6184 7404
rect 6052 7364 6184 7392
rect 6052 7352 6058 7364
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 7248 7364 8677 7392
rect 7248 7352 7254 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10505 7395 10563 7401
rect 9916 7364 10364 7392
rect 9916 7352 9922 7364
rect 10336 7336 10364 7364
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 10551 7364 10977 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 12434 7392 12440 7404
rect 11379 7364 12440 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5534 7324 5540 7336
rect 5491 7296 5540 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 3068 7256 3096 7284
rect 3881 7259 3939 7265
rect 3881 7256 3893 7259
rect 3068 7228 3893 7256
rect 3881 7225 3893 7228
rect 3927 7225 3939 7259
rect 5092 7256 5120 7287
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 5913 7327 5971 7333
rect 5913 7293 5925 7327
rect 5959 7293 5971 7327
rect 8294 7324 8300 7336
rect 8255 7296 8300 7324
rect 5913 7287 5971 7293
rect 5644 7256 5672 7284
rect 5092 7228 5672 7256
rect 3881 7219 3939 7225
rect 2363 7160 3004 7188
rect 3053 7191 3111 7197
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 5258 7188 5264 7200
rect 3099 7160 5264 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5626 7188 5632 7200
rect 5399 7160 5632 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5736 7188 5764 7287
rect 5920 7256 5948 7287
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8527 7296 8585 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8932 7327 8990 7333
rect 8932 7293 8944 7327
rect 8978 7324 8990 7327
rect 9306 7324 9312 7336
rect 8978 7296 9312 7324
rect 8978 7293 8990 7296
rect 8932 7287 8990 7293
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 5994 7256 6000 7268
rect 5920 7228 6000 7256
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6178 7256 6184 7268
rect 6135 7228 6184 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 6457 7259 6515 7265
rect 6457 7225 6469 7259
rect 6503 7256 6515 7259
rect 6914 7256 6920 7268
rect 6503 7228 6920 7256
rect 6503 7225 6515 7228
rect 6457 7219 6515 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 8662 7256 8668 7268
rect 7432 7228 8668 7256
rect 7432 7216 7438 7228
rect 8662 7216 8668 7228
rect 8720 7256 8726 7268
rect 9858 7256 9864 7268
rect 8720 7228 9864 7256
rect 8720 7216 8726 7228
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10244 7256 10272 7287
rect 10318 7284 10324 7336
rect 10376 7284 10382 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10597 7327 10655 7333
rect 10597 7324 10609 7327
rect 10468 7296 10609 7324
rect 10468 7284 10474 7296
rect 10597 7293 10609 7296
rect 10643 7293 10655 7327
rect 10870 7324 10876 7336
rect 10831 7296 10876 7324
rect 10597 7287 10655 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11238 7324 11244 7336
rect 11112 7296 11244 7324
rect 11112 7284 11118 7296
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11480 7296 11897 7324
rect 11480 7284 11486 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 10689 7259 10747 7265
rect 10689 7256 10701 7259
rect 10244 7228 10701 7256
rect 10689 7225 10701 7228
rect 10735 7225 10747 7259
rect 10689 7219 10747 7225
rect 6270 7188 6276 7200
rect 5736 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7188 6334 7200
rect 6638 7188 6644 7200
rect 6328 7160 6644 7188
rect 6328 7148 6334 7160
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8168 7160 8585 7188
rect 8168 7148 8174 7160
rect 8573 7157 8585 7160
rect 8619 7188 8631 7191
rect 11072 7188 11100 7284
rect 8619 7160 11100 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 1104 7098 12328 7120
rect 1104 7046 4723 7098
rect 4775 7046 4787 7098
rect 4839 7046 4851 7098
rect 4903 7046 4915 7098
rect 4967 7046 8464 7098
rect 8516 7046 8528 7098
rect 8580 7046 8592 7098
rect 8644 7046 8656 7098
rect 8708 7046 12328 7098
rect 1104 7024 12328 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3237 6987 3295 6993
rect 3237 6984 3249 6987
rect 2648 6956 3249 6984
rect 2648 6944 2654 6956
rect 3237 6953 3249 6956
rect 3283 6953 3295 6987
rect 3237 6947 3295 6953
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 3936 6956 6592 6984
rect 3936 6944 3942 6956
rect 1412 6888 5304 6916
rect 1412 6857 1440 6888
rect 1670 6857 1676 6860
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6817 1455 6851
rect 1397 6811 1455 6817
rect 1664 6811 1676 6857
rect 1728 6848 1734 6860
rect 1728 6820 1764 6848
rect 1670 6808 1676 6811
rect 1728 6808 1734 6820
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 3896 6857 3924 6888
rect 5276 6860 5304 6888
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 5994 6916 6000 6928
rect 5592 6888 6000 6916
rect 5592 6876 5598 6888
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 6564 6916 6592 6956
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 6733 6987 6791 6993
rect 6733 6984 6745 6987
rect 6696 6956 6745 6984
rect 6696 6944 6702 6956
rect 6733 6953 6745 6956
rect 6779 6953 6791 6987
rect 8846 6984 8852 6996
rect 8807 6956 8852 6984
rect 6733 6947 6791 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 9180 6956 9229 6984
rect 9180 6944 9186 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9217 6947 9275 6953
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 9640 6956 9781 6984
rect 9640 6944 9646 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 10042 6984 10048 6996
rect 9907 6956 10048 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10376 6956 10609 6984
rect 10376 6944 10382 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 10689 6987 10747 6993
rect 10689 6953 10701 6987
rect 10735 6984 10747 6987
rect 10870 6984 10876 6996
rect 10735 6956 10876 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 6914 6916 6920 6928
rect 6564 6888 6920 6916
rect 6914 6876 6920 6888
rect 6972 6876 6978 6928
rect 7098 6925 7104 6928
rect 7092 6916 7104 6925
rect 7059 6888 7104 6916
rect 7092 6879 7104 6888
rect 7098 6876 7104 6879
rect 7156 6876 7162 6928
rect 8665 6919 8723 6925
rect 8665 6885 8677 6919
rect 8711 6916 8723 6919
rect 9674 6916 9680 6928
rect 8711 6888 9680 6916
rect 8711 6885 8723 6888
rect 8665 6879 8723 6885
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 4154 6857 4160 6860
rect 3329 6851 3387 6857
rect 2188 6820 2774 6848
rect 2188 6808 2194 6820
rect 2746 6780 2774 6820
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3881 6851 3939 6857
rect 3375 6820 3556 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 2746 6752 3433 6780
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 2866 6712 2872 6724
rect 2827 6684 2872 6712
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2648 6616 2789 6644
rect 2648 6604 2654 6616
rect 2777 6613 2789 6616
rect 2823 6644 2835 6647
rect 3528 6644 3556 6820
rect 3881 6817 3893 6851
rect 3927 6817 3939 6851
rect 4148 6848 4160 6857
rect 4115 6820 4160 6848
rect 3881 6811 3939 6817
rect 4148 6811 4160 6820
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3896 6780 3924 6811
rect 4154 6808 4160 6811
rect 4212 6808 4218 6860
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5626 6857 5632 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5316 6820 5365 6848
rect 5316 6808 5322 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5620 6848 5632 6857
rect 5587 6820 5632 6848
rect 5353 6811 5411 6817
rect 5620 6811 5632 6820
rect 5626 6808 5632 6811
rect 5684 6808 5690 6860
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 6236 6820 8493 6848
rect 6236 6808 6242 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6817 8815 6851
rect 8757 6811 8815 6817
rect 3660 6752 3924 6780
rect 6825 6783 6883 6789
rect 3660 6740 3666 6752
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 2823 6616 3556 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 3936 6616 5273 6644
rect 3936 6604 3942 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 6840 6644 6868 6743
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8772 6780 8800 6811
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 9088 6820 9137 6848
rect 9088 6808 9094 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 11057 6851 11115 6857
rect 9125 6811 9183 6817
rect 9968 6820 10824 6848
rect 7892 6752 8800 6780
rect 7892 6740 7898 6752
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9858 6780 9864 6792
rect 9364 6752 9864 6780
rect 9364 6740 9370 6752
rect 9858 6740 9864 6752
rect 9916 6780 9922 6792
rect 9968 6789 9996 6820
rect 9953 6783 10011 6789
rect 9953 6780 9965 6783
rect 9916 6752 9965 6780
rect 9916 6740 9922 6752
rect 9953 6749 9965 6752
rect 9999 6749 10011 6783
rect 10410 6780 10416 6792
rect 9953 6743 10011 6749
rect 10060 6752 10416 6780
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 8294 6712 8300 6724
rect 8251 6684 8300 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 9401 6715 9459 6721
rect 9401 6681 9413 6715
rect 9447 6712 9459 6715
rect 10060 6712 10088 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10796 6789 10824 6820
rect 11057 6817 11069 6851
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 9447 6684 10088 6712
rect 10229 6715 10287 6721
rect 9447 6681 9459 6684
rect 9401 6675 9459 6681
rect 10229 6681 10241 6715
rect 10275 6712 10287 6715
rect 11072 6712 11100 6811
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11204 6752 11529 6780
rect 11204 6740 11210 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 10275 6684 11100 6712
rect 10275 6681 10287 6684
rect 10229 6675 10287 6681
rect 7190 6644 7196 6656
rect 6840 6616 7196 6644
rect 5261 6607 5319 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 10836 6616 11161 6644
rect 10836 6604 10842 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11664 6616 11805 6644
rect 11664 6604 11670 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 1104 6554 12328 6576
rect 1104 6502 2852 6554
rect 2904 6502 2916 6554
rect 2968 6502 2980 6554
rect 3032 6502 3044 6554
rect 3096 6502 6594 6554
rect 6646 6502 6658 6554
rect 6710 6502 6722 6554
rect 6774 6502 6786 6554
rect 6838 6502 10335 6554
rect 10387 6502 10399 6554
rect 10451 6502 10463 6554
rect 10515 6502 10527 6554
rect 10579 6502 12328 6554
rect 1104 6480 12328 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3476 6412 3709 6440
rect 3476 6400 3482 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3970 6440 3976 6452
rect 3931 6412 3976 6440
rect 3697 6403 3755 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 5534 6440 5540 6452
rect 4724 6412 5540 6440
rect 2685 6375 2743 6381
rect 2685 6372 2697 6375
rect 1688 6344 2697 6372
rect 1688 6313 1716 6344
rect 2685 6341 2697 6344
rect 2731 6341 2743 6375
rect 2685 6335 2743 6341
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 2188 6276 2329 6304
rect 2188 6264 2194 6276
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 3142 6304 3148 6316
rect 2317 6267 2375 6273
rect 2792 6276 3148 6304
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6205 1547 6239
rect 2332 6236 2360 6267
rect 2406 6236 2412 6248
rect 2332 6208 2412 6236
rect 1489 6199 1547 6205
rect 1504 6168 1532 6199
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2792 6245 2820 6276
rect 3142 6264 3148 6276
rect 3200 6304 3206 6316
rect 3200 6276 4108 6304
rect 3200 6264 3206 6276
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6205 2835 6239
rect 3050 6236 3056 6248
rect 3011 6208 3056 6236
rect 2777 6199 2835 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6205 3387 6239
rect 3329 6199 3387 6205
rect 3234 6168 3240 6180
rect 1504 6140 3240 6168
rect 3234 6128 3240 6140
rect 3292 6128 3298 6180
rect 3344 6168 3372 6199
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 3476 6208 3617 6236
rect 3476 6196 3482 6208
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3605 6199 3663 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4080 6245 4108 6276
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 4157 6199 4215 6205
rect 3970 6168 3976 6180
rect 3344 6140 3976 6168
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1765 6103 1823 6109
rect 1765 6100 1777 6103
rect 1728 6072 1777 6100
rect 1728 6060 1734 6072
rect 1765 6069 1777 6072
rect 1811 6069 1823 6103
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 1765 6063 1823 6069
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 3878 6100 3884 6112
rect 2271 6072 3884 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4172 6100 4200 6199
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4724 6245 4752 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5868 6412 5917 6440
rect 5868 6400 5874 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6512 6412 6561 6440
rect 6512 6400 6518 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7834 6440 7840 6452
rect 7239 6412 7840 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 8168 6412 8217 6440
rect 8168 6400 8174 6412
rect 8205 6409 8217 6412
rect 8251 6440 8263 6443
rect 8294 6440 8300 6452
rect 8251 6412 8300 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 11054 6440 11060 6452
rect 10152 6412 11060 6440
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6341 5043 6375
rect 6086 6372 6092 6384
rect 4985 6335 5043 6341
rect 5460 6344 6092 6372
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 5000 6168 5028 6335
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5460 6313 5488 6344
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6656 6344 7113 6372
rect 5445 6307 5503 6313
rect 5224 6276 5396 6304
rect 5224 6264 5230 6276
rect 5368 6245 5396 6276
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 6656 6304 6684 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7208 6344 7871 6372
rect 7208 6316 7236 6344
rect 5675 6276 6684 6304
rect 6733 6307 6791 6313
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 6564 6248 6592 6276
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 6779 6276 7144 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6205 5411 6239
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5353 6199 5411 6205
rect 5736 6208 5825 6236
rect 5000 6140 5496 6168
rect 5258 6100 5264 6112
rect 4172 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5468 6100 5496 6140
rect 5736 6100 5764 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6178 6236 6184 6248
rect 6135 6208 6184 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 6472 6168 6500 6199
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6696 6208 6837 6236
rect 6696 6196 6702 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 6472 6140 6929 6168
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 7116 6168 7144 6276
rect 7190 6264 7196 6316
rect 7248 6264 7254 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7432 6276 7757 6304
rect 7432 6264 7438 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7843 6304 7871 6344
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 7843 6276 8493 6304
rect 7745 6267 7803 6273
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7340 6208 7573 6236
rect 7340 6196 7346 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7892 6208 8033 6236
rect 7892 6196 7898 6208
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8496 6236 8524 6267
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10152 6313 10180 6412
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10100 6276 10149 6304
rect 10100 6264 10106 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11296 6276 11928 6304
rect 11296 6264 11302 6276
rect 10060 6236 10088 6264
rect 11900 6245 11928 6276
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 8496 6208 10088 6236
rect 11532 6208 11713 6236
rect 8021 6199 8079 6205
rect 8110 6168 8116 6180
rect 7116 6140 8116 6168
rect 6917 6131 6975 6137
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 8748 6171 8806 6177
rect 8748 6137 8760 6171
rect 8794 6168 8806 6171
rect 8938 6168 8944 6180
rect 8794 6140 8944 6168
rect 8794 6137 8806 6140
rect 8748 6131 8806 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 10404 6171 10462 6177
rect 10404 6137 10416 6171
rect 10450 6168 10462 6171
rect 10686 6168 10692 6180
rect 10450 6140 10692 6168
rect 10450 6137 10462 6140
rect 10404 6131 10462 6137
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 6730 6100 6736 6112
rect 5468 6072 5764 6100
rect 6691 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 7098 6100 7104 6112
rect 7011 6072 7104 6100
rect 7098 6060 7104 6072
rect 7156 6100 7162 6112
rect 7374 6100 7380 6112
rect 7156 6072 7380 6100
rect 7156 6060 7162 6072
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7653 6103 7711 6109
rect 7653 6069 7665 6103
rect 7699 6100 7711 6103
rect 7926 6100 7932 6112
rect 7699 6072 7932 6100
rect 7699 6069 7711 6072
rect 7653 6063 7711 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9861 6103 9919 6109
rect 9861 6100 9873 6103
rect 9640 6072 9873 6100
rect 9640 6060 9646 6072
rect 9861 6069 9873 6072
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11532 6109 11560 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11112 6072 11529 6100
rect 11112 6060 11118 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11517 6063 11575 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 1104 6010 12328 6032
rect 1104 5958 4723 6010
rect 4775 5958 4787 6010
rect 4839 5958 4851 6010
rect 4903 5958 4915 6010
rect 4967 5958 8464 6010
rect 8516 5958 8528 6010
rect 8580 5958 8592 6010
rect 8644 5958 8656 6010
rect 8708 5958 12328 6010
rect 1104 5936 12328 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1452 5868 1777 5896
rect 1452 5856 1458 5868
rect 1765 5865 1777 5868
rect 1811 5865 1823 5899
rect 1765 5859 1823 5865
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 2096 5868 2421 5896
rect 2096 5856 2102 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3476 5868 3893 5896
rect 3476 5856 3482 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 6638 5896 6644 5908
rect 5767 5868 6644 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7926 5896 7932 5908
rect 7887 5868 7932 5896
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8110 5896 8116 5908
rect 8071 5868 8116 5896
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 10686 5896 10692 5908
rect 8588 5868 9720 5896
rect 10647 5868 10692 5896
rect 3234 5828 3240 5840
rect 3068 5800 3240 5828
rect 937 5763 995 5769
rect 937 5729 949 5763
rect 983 5760 995 5763
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 983 5732 1593 5760
rect 983 5729 995 5732
rect 937 5723 995 5729
rect 1581 5729 1593 5732
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 1728 5732 1773 5760
rect 1728 5720 1734 5732
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 2406 5760 2412 5772
rect 2188 5732 2412 5760
rect 2188 5720 2194 5732
rect 2406 5720 2412 5732
rect 2464 5760 2470 5772
rect 2464 5732 2636 5760
rect 2464 5720 2470 5732
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2608 5701 2636 5732
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3068 5769 3096 5800
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 3344 5800 3648 5828
rect 2961 5763 3019 5769
rect 2961 5760 2973 5763
rect 2740 5732 2973 5760
rect 2740 5720 2746 5732
rect 2961 5729 2973 5732
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5729 3111 5763
rect 3344 5760 3372 5800
rect 3053 5723 3111 5729
rect 3160 5732 3372 5760
rect 3421 5763 3479 5769
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3160 5692 3188 5732
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 3513 5763 3571 5769
rect 3513 5760 3525 5763
rect 3467 5732 3525 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 3513 5729 3525 5732
rect 3559 5729 3571 5763
rect 3620 5760 3648 5800
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3844 5800 4261 5828
rect 3844 5788 3850 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 5261 5831 5319 5837
rect 5261 5797 5273 5831
rect 5307 5828 5319 5831
rect 5442 5828 5448 5840
rect 5307 5800 5448 5828
rect 5307 5797 5319 5800
rect 5261 5791 5319 5797
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 5902 5788 5908 5840
rect 5960 5828 5966 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 5960 5800 6101 5828
rect 5960 5788 5966 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 6181 5831 6239 5837
rect 6181 5797 6193 5831
rect 6227 5828 6239 5831
rect 6270 5828 6276 5840
rect 6227 5800 6276 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 6730 5788 6736 5840
rect 6788 5837 6794 5840
rect 6788 5831 6852 5837
rect 6788 5797 6806 5831
rect 6840 5797 6852 5831
rect 6788 5791 6852 5797
rect 6788 5788 6794 5791
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7834 5828 7840 5840
rect 6972 5800 7840 5828
rect 6972 5788 6978 5800
rect 7834 5788 7840 5800
rect 7892 5788 7898 5840
rect 4709 5763 4767 5769
rect 3620 5732 4568 5760
rect 3513 5723 3571 5729
rect 2639 5664 3188 5692
rect 3237 5695 3295 5701
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 4154 5692 4160 5704
rect 3283 5664 4160 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4540 5701 4568 5732
rect 4709 5729 4721 5763
rect 4755 5760 4767 5763
rect 4890 5760 4896 5772
rect 4755 5732 4896 5760
rect 4755 5729 4767 5732
rect 4709 5723 4767 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5074 5760 5080 5772
rect 5035 5732 5080 5760
rect 5074 5720 5080 5732
rect 5132 5720 5138 5772
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7282 5760 7288 5772
rect 6595 5732 7288 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7944 5760 7972 5856
rect 8588 5772 8616 5868
rect 8938 5828 8944 5840
rect 8899 5800 8944 5828
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7944 5732 8033 5760
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8294 5760 8300 5772
rect 8251 5732 8300 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5729 8447 5763
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8389 5723 8447 5729
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 4571 5664 6377 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 1394 5624 1400 5636
rect 1355 5596 1400 5624
rect 1394 5584 1400 5596
rect 1452 5584 1458 5636
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3421 5627 3479 5633
rect 3108 5596 3372 5624
rect 3108 5584 3114 5596
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3234 5556 3240 5568
rect 3191 5528 3240 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3344 5556 3372 5596
rect 3421 5593 3433 5627
rect 3467 5624 3479 5627
rect 6086 5624 6092 5636
rect 3467 5596 6092 5624
rect 3467 5593 3479 5596
rect 3421 5587 3479 5593
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 6380 5624 6408 5655
rect 6546 5624 6552 5636
rect 6380 5596 6552 5624
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 7650 5584 7656 5636
rect 7708 5624 7714 5636
rect 7834 5624 7840 5636
rect 7708 5596 7840 5624
rect 7708 5584 7714 5596
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 8404 5624 8432 5723
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 8711 5732 9076 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8527 5664 8953 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 9048 5692 9076 5732
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9180 5732 9225 5760
rect 9180 5720 9186 5732
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9585 5763 9643 5769
rect 9585 5760 9597 5763
rect 9548 5732 9597 5760
rect 9548 5720 9554 5732
rect 9585 5729 9597 5732
rect 9631 5729 9643 5763
rect 9692 5760 9720 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11238 5828 11244 5840
rect 11103 5800 11244 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9692 5732 9781 5760
rect 9585 5723 9643 5729
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 10413 5763 10471 5769
rect 9916 5732 9961 5760
rect 9916 5720 9922 5732
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10778 5760 10784 5772
rect 10459 5732 10784 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 10919 5732 11897 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 11885 5729 11897 5732
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9048 5664 9229 5692
rect 8941 5655 8999 5661
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9723 5664 10149 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10689 5695 10747 5701
rect 10284 5664 10640 5692
rect 10284 5652 10290 5664
rect 9582 5624 9588 5636
rect 8404 5596 9588 5624
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 10505 5627 10563 5633
rect 10505 5624 10517 5627
rect 9968 5596 10517 5624
rect 5442 5556 5448 5568
rect 3344 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 8294 5556 8300 5568
rect 5675 5528 8300 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 9674 5556 9680 5568
rect 8803 5528 9680 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 9674 5516 9680 5528
rect 9732 5556 9738 5568
rect 9968 5565 9996 5596
rect 10505 5593 10517 5596
rect 10551 5593 10563 5627
rect 10612 5624 10640 5664
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 11790 5692 11796 5704
rect 10735 5664 11796 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 10778 5624 10784 5636
rect 10612 5596 10784 5624
rect 10505 5587 10563 5593
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11333 5627 11391 5633
rect 11333 5624 11345 5627
rect 10928 5596 11345 5624
rect 10928 5584 10934 5596
rect 11333 5593 11345 5596
rect 11379 5593 11391 5627
rect 11333 5587 11391 5593
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 9732 5528 9965 5556
rect 9732 5516 9738 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 10686 5556 10692 5568
rect 10091 5528 10692 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 11020 5528 11621 5556
rect 11020 5516 11026 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 11609 5519 11667 5525
rect 1104 5466 12328 5488
rect 1104 5414 2852 5466
rect 2904 5414 2916 5466
rect 2968 5414 2980 5466
rect 3032 5414 3044 5466
rect 3096 5414 6594 5466
rect 6646 5414 6658 5466
rect 6710 5414 6722 5466
rect 6774 5414 6786 5466
rect 6838 5414 10335 5466
rect 10387 5414 10399 5466
rect 10451 5414 10463 5466
rect 10515 5414 10527 5466
rect 10579 5414 12328 5466
rect 1104 5392 12328 5414
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2777 5355 2835 5361
rect 2777 5352 2789 5355
rect 2556 5324 2789 5352
rect 2556 5312 2562 5324
rect 2777 5321 2789 5324
rect 2823 5321 2835 5355
rect 2777 5315 2835 5321
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4396 5324 4537 5352
rect 4396 5312 4402 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 4525 5315 4583 5321
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 8665 5355 8723 5361
rect 6319 5324 8616 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 2961 5287 3019 5293
rect 2961 5284 2973 5287
rect 2740 5256 2973 5284
rect 2740 5244 2746 5256
rect 2961 5253 2973 5256
rect 3007 5253 3019 5287
rect 2961 5247 3019 5253
rect 4614 5244 4620 5296
rect 4672 5284 4678 5296
rect 4890 5284 4896 5296
rect 4672 5256 4896 5284
rect 4672 5244 4678 5256
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 5350 5284 5356 5296
rect 5307 5256 5356 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 7469 5287 7527 5293
rect 7469 5284 7481 5287
rect 6788 5256 7481 5284
rect 6788 5244 6794 5256
rect 7469 5253 7481 5256
rect 7515 5253 7527 5287
rect 7469 5247 7527 5253
rect 7098 5216 7104 5228
rect 7059 5188 7104 5216
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7699 5188 8309 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 661 5151 719 5157
rect 661 5117 673 5151
rect 707 5148 719 5151
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 707 5120 1409 5148
rect 707 5117 719 5120
rect 661 5111 719 5117
rect 1397 5117 1409 5120
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 1412 5012 1440 5111
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2096 5120 2881 5148
rect 2096 5108 2102 5120
rect 2869 5117 2881 5120
rect 2915 5117 2927 5151
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2869 5111 2927 5117
rect 3068 5120 3157 5148
rect 1664 5083 1722 5089
rect 1664 5049 1676 5083
rect 1710 5080 1722 5083
rect 2406 5080 2412 5092
rect 1710 5052 2412 5080
rect 1710 5049 1722 5052
rect 1664 5043 1722 5049
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 3068 5012 3096 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3401 5151 3459 5157
rect 3401 5148 3413 5151
rect 3292 5120 3413 5148
rect 3292 5108 3298 5120
rect 3401 5117 3413 5120
rect 3447 5117 3459 5151
rect 3401 5111 3459 5117
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4706 5148 4712 5160
rect 4663 5120 4712 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4706 5108 4712 5120
rect 4764 5148 4770 5160
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 4764 5120 5641 5148
rect 4764 5108 4770 5120
rect 5629 5117 5641 5120
rect 5675 5148 5687 5151
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5675 5120 5825 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5813 5117 5825 5120
rect 5859 5148 5871 5151
rect 6822 5148 6828 5160
rect 5859 5120 6828 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 6880 5120 7144 5148
rect 6880 5108 6886 5120
rect 5074 5080 5080 5092
rect 5035 5052 5080 5080
rect 5074 5040 5080 5052
rect 5132 5080 5138 5092
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 5132 5052 5457 5080
rect 5132 5040 5138 5052
rect 5445 5049 5457 5052
rect 5491 5049 5503 5083
rect 5445 5043 5503 5049
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6328 5052 7021 5080
rect 6328 5040 6334 5052
rect 7009 5049 7021 5052
rect 7055 5049 7067 5083
rect 7116 5080 7144 5120
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 7929 5151 7987 5157
rect 7432 5120 7477 5148
rect 7432 5108 7438 5120
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 8202 5148 8208 5160
rect 8163 5120 8208 5148
rect 7929 5111 7987 5117
rect 7944 5080 7972 5111
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8386 5148 8392 5160
rect 8299 5120 8392 5148
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8404 5080 8432 5108
rect 7116 5052 7972 5080
rect 8128 5052 8432 5080
rect 8588 5080 8616 5324
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 9122 5352 9128 5364
rect 8711 5324 9128 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 9858 5352 9864 5364
rect 9631 5324 9864 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 9968 5324 11529 5352
rect 9490 5284 9496 5296
rect 9140 5256 9496 5284
rect 9140 5225 9168 5256
rect 9490 5244 9496 5256
rect 9548 5284 9554 5296
rect 9968 5284 9996 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 9548 5256 9996 5284
rect 9548 5244 9554 5256
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9306 5216 9312 5228
rect 9267 5188 9312 5216
rect 9125 5179 9183 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10042 5216 10048 5228
rect 9732 5188 10048 5216
rect 9732 5176 9738 5188
rect 10042 5176 10048 5188
rect 10100 5216 10106 5228
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 10100 5188 10149 5216
rect 10100 5176 10106 5188
rect 10137 5185 10149 5188
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8996 5120 9045 5148
rect 8996 5108 9002 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10226 5148 10232 5160
rect 9539 5120 10232 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10404 5151 10462 5157
rect 10404 5117 10416 5151
rect 10450 5148 10462 5151
rect 10686 5148 10692 5160
rect 10450 5120 10692 5148
rect 10450 5117 10462 5120
rect 10404 5111 10462 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11572 5120 11805 5148
rect 11572 5108 11578 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 9122 5080 9128 5092
rect 8588 5052 9128 5080
rect 7009 5043 7067 5049
rect 3602 5012 3608 5024
rect 1412 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4120 4984 4813 5012
rect 4120 4972 4126 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 5902 5012 5908 5024
rect 5863 4984 5908 5012
rect 4801 4975 4859 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6822 5012 6828 5024
rect 6595 4984 6828 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 7466 5012 7472 5024
rect 6963 4984 7472 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7650 5012 7656 5024
rect 7611 4984 7656 5012
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8128 5021 8156 5052
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 9858 5080 9864 5092
rect 9819 5052 9864 5080
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 10318 5080 10324 5092
rect 10244 5052 10324 5080
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7984 4984 8125 5012
rect 7984 4972 7990 4984
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10244 5012 10272 5052
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 11977 5083 12035 5089
rect 11977 5049 11989 5083
rect 12023 5080 12035 5083
rect 13262 5080 13268 5092
rect 12023 5052 13268 5080
rect 12023 5049 12035 5052
rect 11977 5043 12035 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 9999 4984 10272 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 1104 4922 12328 4944
rect 1104 4870 4723 4922
rect 4775 4870 4787 4922
rect 4839 4870 4851 4922
rect 4903 4870 4915 4922
rect 4967 4870 8464 4922
rect 8516 4870 8528 4922
rect 8580 4870 8592 4922
rect 8644 4870 8656 4922
rect 8708 4870 12328 4922
rect 1104 4848 12328 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 2556 4780 2820 4808
rect 2556 4768 2562 4780
rect 2593 4743 2651 4749
rect 2593 4740 2605 4743
rect 2148 4712 2605 4740
rect 198 4632 204 4684
rect 256 4672 262 4684
rect 2148 4681 2176 4712
rect 2593 4709 2605 4712
rect 2639 4709 2651 4743
rect 2593 4703 2651 4709
rect 1489 4675 1547 4681
rect 1489 4672 1501 4675
rect 256 4644 1501 4672
rect 256 4632 262 4644
rect 1489 4641 1501 4644
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4641 2191 4675
rect 2498 4672 2504 4684
rect 2459 4644 2504 4672
rect 2133 4635 2191 4641
rect 1872 4604 1900 4635
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 2792 4681 2820 4780
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 3970 4808 3976 4820
rect 3292 4780 3976 4808
rect 3292 4768 3298 4780
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4212 4780 4353 4808
rect 4212 4768 4218 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 5350 4808 5356 4820
rect 4341 4771 4399 4777
rect 4908 4780 5356 4808
rect 4080 4740 4108 4768
rect 4908 4749 4936 4780
rect 5350 4768 5356 4780
rect 5408 4808 5414 4820
rect 5408 4780 6684 4808
rect 5408 4768 5414 4780
rect 4893 4743 4951 4749
rect 3160 4712 4476 4740
rect 3160 4684 3188 4712
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4641 2835 4675
rect 2777 4635 2835 4641
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 3142 4672 3148 4684
rect 3007 4644 3148 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3418 4672 3424 4684
rect 3283 4644 3424 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3786 4672 3792 4684
rect 3559 4644 3792 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 3970 4672 3976 4684
rect 3931 4644 3976 4672
rect 3970 4632 3976 4644
rect 4028 4632 4034 4684
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 4120 4644 4169 4672
rect 4120 4632 4126 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4338 4672 4344 4684
rect 4295 4644 4344 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4448 4681 4476 4712
rect 4893 4709 4905 4743
rect 4939 4709 4951 4743
rect 4893 4703 4951 4709
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 6546 4740 6552 4752
rect 5684 4712 6552 4740
rect 5684 4700 5690 4712
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 6656 4740 6684 4780
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7466 4808 7472 4820
rect 7340 4780 7472 4808
rect 7340 4768 7346 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8260 4780 8677 4808
rect 8260 4768 8266 4780
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 6716 4743 6774 4749
rect 6716 4740 6728 4743
rect 6656 4712 6728 4740
rect 6716 4709 6728 4712
rect 6762 4709 6774 4743
rect 6716 4703 6774 4709
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 7552 4743 7610 4749
rect 6972 4712 7512 4740
rect 6972 4700 6978 4712
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5425 4675 5483 4681
rect 5425 4672 5437 4675
rect 5040 4644 5437 4672
rect 5040 4632 5046 4644
rect 5425 4641 5437 4644
rect 5471 4641 5483 4675
rect 5425 4635 5483 4641
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6880 4644 7021 4672
rect 6880 4632 6886 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 7009 4635 7067 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7484 4672 7512 4712
rect 7552 4709 7564 4743
rect 7598 4740 7610 4743
rect 7650 4740 7656 4752
rect 7598 4712 7656 4740
rect 7598 4709 7610 4712
rect 7552 4703 7610 4709
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 8757 4675 8815 4681
rect 7484 4644 8340 4672
rect 2314 4604 2320 4616
rect 1872 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2455 4576 2881 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 3752 4576 5181 4604
rect 3752 4564 3758 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 6748 4576 7236 4604
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 6748 4536 6776 4576
rect 6914 4536 6920 4548
rect 4755 4508 5212 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2225 4471 2283 4477
rect 2225 4437 2237 4471
rect 2271 4468 2283 4471
rect 3418 4468 3424 4480
rect 2271 4440 3424 4468
rect 2271 4437 2283 4440
rect 2225 4431 2283 4437
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 3602 4428 3608 4480
rect 3660 4468 3666 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 3660 4440 4077 4468
rect 3660 4428 3666 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 4065 4431 4123 4437
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4948 4440 4997 4468
rect 4948 4428 4954 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 5184 4468 5212 4508
rect 6104 4508 6776 4536
rect 6875 4508 6920 4536
rect 6104 4480 6132 4508
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 5442 4468 5448 4480
rect 5184 4440 5448 4468
rect 4985 4431 5043 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 6086 4428 6092 4480
rect 6144 4428 6150 4480
rect 6362 4428 6368 4480
rect 6420 4468 6426 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6420 4440 6561 4468
rect 6420 4428 6426 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 7098 4468 7104 4480
rect 7059 4440 7104 4468
rect 6549 4431 6607 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7208 4468 7236 4576
rect 8312 4536 8340 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9140 4672 9168 4771
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 10284 4780 10425 4808
rect 10284 4768 10290 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10413 4771 10471 4777
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 10652 4780 10793 4808
rect 10652 4768 10658 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 10781 4771 10839 4777
rect 9582 4740 9588 4752
rect 9543 4712 9588 4740
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 10045 4743 10103 4749
rect 10045 4709 10057 4743
rect 10091 4740 10103 4743
rect 10870 4740 10876 4752
rect 10091 4712 10876 4740
rect 10091 4709 10103 4712
rect 10045 4703 10103 4709
rect 10870 4700 10876 4712
rect 10928 4700 10934 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11388 4712 11437 4740
rect 11388 4700 11394 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 9490 4672 9496 4684
rect 8803 4644 9168 4672
rect 9451 4644 9496 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 11793 4675 11851 4681
rect 9692 4644 11008 4672
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9692 4613 9720 4644
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9364 4576 9689 4604
rect 9364 4564 9370 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 9677 4567 9735 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 10980 4613 11008 4644
rect 11793 4641 11805 4675
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11808 4536 11836 4635
rect 8312 4508 11836 4536
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12526 4536 12532 4548
rect 12023 4508 12532 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 8570 4468 8576 4480
rect 7208 4440 8576 4468
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8849 4471 8907 4477
rect 8849 4437 8861 4471
rect 8895 4468 8907 4471
rect 8938 4468 8944 4480
rect 8895 4440 8944 4468
rect 8895 4437 8907 4440
rect 8849 4431 8907 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9490 4428 9496 4480
rect 9548 4468 9554 4480
rect 9674 4468 9680 4480
rect 9548 4440 9680 4468
rect 9548 4428 9554 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 10008 4440 10149 4468
rect 10008 4428 10014 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 12894 4468 12900 4480
rect 11563 4440 12900 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 1104 4378 12328 4400
rect 1104 4326 2852 4378
rect 2904 4326 2916 4378
rect 2968 4326 2980 4378
rect 3032 4326 3044 4378
rect 3096 4326 6594 4378
rect 6646 4326 6658 4378
rect 6710 4326 6722 4378
rect 6774 4326 6786 4378
rect 6838 4326 10335 4378
rect 10387 4326 10399 4378
rect 10451 4326 10463 4378
rect 10515 4326 10527 4378
rect 10579 4326 12328 4378
rect 1104 4304 12328 4326
rect 474 4264 480 4276
rect 435 4236 480 4264
rect 474 4224 480 4236
rect 532 4224 538 4276
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2498 4264 2504 4276
rect 2271 4236 2504 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 3418 4264 3424 4276
rect 3331 4236 3424 4264
rect 3418 4224 3424 4236
rect 3476 4264 3482 4276
rect 4890 4264 4896 4276
rect 3476 4236 4896 4264
rect 3476 4224 3482 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5626 4264 5632 4276
rect 5491 4236 5632 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 5810 4264 5816 4276
rect 5767 4236 5816 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 6641 4267 6699 4273
rect 6641 4264 6653 4267
rect 5920 4236 6653 4264
rect 2130 4156 2136 4208
rect 2188 4196 2194 4208
rect 2188 4168 2820 4196
rect 2188 4156 2194 4168
rect 106 4088 112 4140
rect 164 4088 170 4140
rect 474 4088 480 4140
rect 532 4128 538 4140
rect 934 4128 940 4140
rect 532 4100 940 4128
rect 532 4088 538 4100
rect 934 4088 940 4100
rect 992 4088 998 4140
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2498 4128 2504 4140
rect 2004 4100 2504 4128
rect 2004 4088 2010 4100
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2792 4137 2820 4168
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3436 4196 3464 4224
rect 3016 4168 3464 4196
rect 3016 4156 3022 4168
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 3660 4100 3705 4128
rect 3660 4088 3666 4100
rect 124 4060 152 4088
rect 1118 4060 1124 4072
rect 124 4032 1124 4060
rect 1118 4020 1124 4032
rect 1176 4020 1182 4072
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 2130 4060 2136 4072
rect 1719 4032 2136 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3050 4060 3056 4072
rect 2731 4032 3056 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3200 4032 3249 4060
rect 3200 4020 3206 4032
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3694 4060 3700 4072
rect 3384 4032 3429 4060
rect 3655 4032 3700 4060
rect 3384 4020 3390 4032
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 5920 4060 5948 4236
rect 6641 4233 6653 4236
rect 6687 4233 6699 4267
rect 6641 4227 6699 4233
rect 6748 4236 7052 4264
rect 5997 4199 6055 4205
rect 5997 4165 6009 4199
rect 6043 4196 6055 4199
rect 6086 4196 6092 4208
rect 6043 4168 6092 4196
rect 6043 4165 6055 4168
rect 5997 4159 6055 4165
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 6362 4156 6368 4208
rect 6420 4196 6426 4208
rect 6748 4196 6776 4236
rect 6420 4168 6776 4196
rect 6420 4156 6426 4168
rect 6546 4128 6552 4140
rect 3844 4032 5396 4060
rect 3844 4020 3850 4032
rect 106 3952 112 4004
rect 164 3992 170 4004
rect 1489 3995 1547 4001
rect 1489 3992 1501 3995
rect 164 3964 1501 3992
rect 164 3952 170 3964
rect 1489 3961 1501 3964
rect 1535 3961 1547 3995
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 1489 3955 1547 3961
rect 1596 3964 1869 3992
rect 14 3884 20 3936
rect 72 3924 78 3936
rect 1596 3924 1624 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 1857 3955 1915 3961
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 3942 3995 4000 4001
rect 3942 3992 3954 3995
rect 3651 3964 3954 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 3942 3961 3954 3964
rect 3988 3961 4000 3995
rect 3942 3955 4000 3961
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5368 3992 5396 4032
rect 5736 4032 5948 4060
rect 6012 4100 6552 4128
rect 5534 3992 5540 4004
rect 5040 3964 5304 3992
rect 5368 3964 5540 3992
rect 5040 3952 5046 3964
rect 1946 3924 1952 3936
rect 72 3896 1624 3924
rect 1907 3896 1952 3924
rect 72 3884 78 3896
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4120 3896 5089 3924
rect 4120 3884 4126 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5276 3924 5304 3964
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 5736 3924 5764 4032
rect 5276 3896 5764 3924
rect 6012 3924 6040 4100
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6736 4131 6794 4137
rect 6736 4097 6748 4131
rect 6782 4097 6794 4131
rect 7024 4128 7052 4236
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7432 4236 7573 4264
rect 7432 4224 7438 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 9490 4264 9496 4276
rect 7561 4227 7619 4233
rect 9148 4236 9496 4264
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 9033 4199 9091 4205
rect 9033 4196 9045 4199
rect 7340 4168 9045 4196
rect 7340 4156 7346 4168
rect 9033 4165 9045 4168
rect 9079 4165 9091 4199
rect 9033 4159 9091 4165
rect 6736 4091 6794 4097
rect 6932 4100 7052 4128
rect 7377 4131 7435 4137
rect 6086 4020 6092 4072
rect 6144 4060 6150 4072
rect 6273 4063 6331 4069
rect 6273 4060 6285 4063
rect 6144 4032 6285 4060
rect 6144 4020 6150 4032
rect 6273 4029 6285 4032
rect 6319 4029 6331 4063
rect 6273 4023 6331 4029
rect 6457 4063 6515 4069
rect 6457 4029 6469 4063
rect 6503 4060 6515 4063
rect 6503 4032 6684 4060
rect 6503 4029 6515 4032
rect 6457 4023 6515 4029
rect 6086 3924 6092 3936
rect 6012 3896 6092 3924
rect 5077 3887 5135 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6656 3924 6684 4032
rect 6748 3992 6776 4091
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 6932 4060 6960 4100
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 8294 4128 8300 4140
rect 7423 4100 8300 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8846 4128 8852 4140
rect 8527 4100 8852 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 6871 4032 6960 4060
rect 7009 4063 7067 4069
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7055 4032 7420 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7392 4004 7420 4032
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 7524 4032 7569 4060
rect 7524 4020 7530 4032
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 8110 4060 8116 4072
rect 8071 4032 8116 4060
rect 7929 4023 7987 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8386 4060 8392 4072
rect 8312 4032 8392 4060
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 6748 3964 6929 3992
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 7374 3952 7380 4004
rect 7432 3952 7438 4004
rect 8312 4001 8340 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8662 4060 8668 4072
rect 8623 4032 8668 4060
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 8938 4060 8944 4072
rect 8899 4032 8944 4060
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9148 4060 9176 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 12158 4264 12164 4276
rect 9640 4236 12164 4264
rect 9640 4224 9646 4236
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 9306 4196 9312 4208
rect 9232 4168 9312 4196
rect 9232 4137 9260 4168
rect 9306 4156 9312 4168
rect 9364 4156 9370 4208
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 11974 4196 11980 4208
rect 10744 4168 11980 4196
rect 10744 4156 10750 4168
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 12618 4128 12624 4140
rect 11195 4100 12624 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 9148 4032 9321 4060
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10100 4032 10977 4060
rect 10100 4020 10106 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11698 4060 11704 4072
rect 11379 4032 11704 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 11882 4060 11888 4072
rect 11839 4032 11888 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 8297 3995 8355 4001
rect 8297 3961 8309 3995
rect 8343 3961 8355 3995
rect 8297 3955 8355 3961
rect 9217 3995 9275 4001
rect 9217 3961 9229 3995
rect 9263 3992 9275 3995
rect 9554 3995 9612 4001
rect 9554 3992 9566 3995
rect 9263 3964 9566 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 9554 3961 9566 3964
rect 9600 3961 9612 3995
rect 9554 3955 9612 3961
rect 10226 3952 10232 4004
rect 10284 3992 10290 4004
rect 11238 3992 11244 4004
rect 10284 3964 11244 3992
rect 10284 3952 10290 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 11517 3995 11575 4001
rect 11517 3961 11529 3995
rect 11563 3992 11575 3995
rect 12066 3992 12072 4004
rect 11563 3964 12072 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 7098 3924 7104 3936
rect 6656 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9674 3924 9680 3936
rect 8803 3896 9680 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10100 3896 10701 3924
rect 10100 3884 10106 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11756 3896 11897 3924
rect 11756 3884 11762 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 382 3816 388 3868
rect 440 3856 446 3868
rect 934 3856 940 3868
rect 440 3828 940 3856
rect 440 3816 446 3828
rect 934 3816 940 3828
rect 992 3816 998 3868
rect 1104 3834 12328 3856
rect 1104 3782 4723 3834
rect 4775 3782 4787 3834
rect 4839 3782 4851 3834
rect 4903 3782 4915 3834
rect 4967 3782 8464 3834
rect 8516 3782 8528 3834
rect 8580 3782 8592 3834
rect 8644 3782 8656 3834
rect 8708 3782 12328 3834
rect 1104 3760 12328 3782
rect 382 3680 388 3732
rect 440 3720 446 3732
rect 477 3723 535 3729
rect 477 3720 489 3723
rect 440 3692 489 3720
rect 440 3680 446 3692
rect 477 3689 489 3692
rect 523 3689 535 3723
rect 477 3683 535 3689
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3050 3720 3056 3732
rect 2823 3692 3056 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3384 3692 3985 3720
rect 3384 3680 3390 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 3973 3683 4031 3689
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 7282 3720 7288 3732
rect 4212 3692 4384 3720
rect 4212 3680 4218 3692
rect 1664 3655 1722 3661
rect 1664 3621 1676 3655
rect 1710 3652 1722 3655
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 1710 3624 3157 3652
rect 1710 3621 1722 3624
rect 1664 3615 1722 3621
rect 3145 3621 3157 3624
rect 3191 3621 3203 3655
rect 3252 3652 3280 3680
rect 3786 3652 3792 3664
rect 3252 3624 3792 3652
rect 3145 3615 3203 3621
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 661 3587 719 3593
rect 661 3553 673 3587
rect 707 3584 719 3587
rect 1397 3587 1455 3593
rect 1397 3584 1409 3587
rect 707 3556 1409 3584
rect 707 3553 719 3556
rect 661 3547 719 3553
rect 1397 3553 1409 3556
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 2884 3448 2912 3547
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 3016 3556 3061 3584
rect 3016 3544 3022 3556
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 3513 3587 3571 3593
rect 3292 3556 3337 3584
rect 3292 3544 3298 3556
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3602 3584 3608 3596
rect 3559 3556 3608 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 3878 3584 3884 3596
rect 3839 3556 3884 3584
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 4356 3593 4384 3692
rect 4724 3692 7288 3720
rect 4724 3593 4752 3692
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 7466 3720 7472 3732
rect 7423 3692 7472 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 7926 3720 7932 3732
rect 7791 3692 7932 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9398 3720 9404 3732
rect 9180 3692 9404 3720
rect 9180 3680 9186 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10781 3723 10839 3729
rect 9916 3692 10732 3720
rect 9916 3680 9922 3692
rect 5261 3655 5319 3661
rect 5261 3652 5273 3655
rect 4816 3624 5273 3652
rect 4816 3593 4844 3624
rect 5261 3621 5273 3624
rect 5307 3621 5319 3655
rect 6641 3655 6699 3661
rect 6641 3652 6653 3655
rect 5261 3615 5319 3621
rect 6196 3624 6653 3652
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4709 3587 4767 3593
rect 4387 3556 4660 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 4172 3516 4200 3547
rect 4430 3516 4436 3528
rect 4172 3488 4436 3516
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 3605 3451 3663 3457
rect 3605 3448 3617 3451
rect 2884 3420 3617 3448
rect 3605 3417 3617 3420
rect 3651 3417 3663 3451
rect 3605 3411 3663 3417
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4632 3448 4660 3556
rect 4709 3553 4721 3587
rect 4755 3553 4767 3587
rect 4709 3547 4767 3553
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 5166 3584 5172 3596
rect 4948 3556 4993 3584
rect 5127 3556 5172 3584
rect 4948 3544 4954 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5902 3584 5908 3596
rect 5675 3556 5908 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5123 3488 5549 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 5644 3448 5672 3547
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6086 3584 6092 3596
rect 6012 3556 6092 3584
rect 4212 3420 4384 3448
rect 4632 3420 5672 3448
rect 4212 3408 4218 3420
rect 845 3383 903 3389
rect 845 3349 857 3383
rect 891 3380 903 3383
rect 2682 3380 2688 3392
rect 891 3352 2688 3380
rect 891 3349 903 3352
rect 845 3343 903 3349
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 3510 3380 3516 3392
rect 3375 3352 3516 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 4028 3352 4261 3380
rect 4028 3340 4034 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 4356 3380 4384 3420
rect 4890 3380 4896 3392
rect 4356 3352 4896 3380
rect 4249 3343 4307 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5074 3380 5080 3392
rect 5031 3352 5080 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 6012 3380 6040 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6196 3593 6224 3624
rect 6641 3621 6653 3624
rect 6687 3621 6699 3655
rect 8757 3655 8815 3661
rect 8757 3652 8769 3655
rect 6641 3615 6699 3621
rect 8036 3624 8769 3652
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 7190 3584 7196 3596
rect 6595 3556 7196 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8036 3584 8064 3624
rect 8757 3621 8769 3624
rect 8803 3621 8815 3655
rect 8757 3615 8815 3621
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9217 3655 9275 3661
rect 9217 3652 9229 3655
rect 8996 3624 9229 3652
rect 8996 3612 9002 3624
rect 9217 3621 9229 3624
rect 9263 3621 9275 3655
rect 9217 3615 9275 3621
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 9548 3624 9597 3652
rect 9548 3612 9554 3624
rect 9585 3621 9597 3624
rect 9631 3621 9643 3655
rect 9585 3615 9643 3621
rect 9766 3612 9772 3664
rect 9824 3652 9830 3664
rect 9953 3655 10011 3661
rect 9953 3652 9965 3655
rect 9824 3624 9965 3652
rect 9824 3612 9830 3624
rect 9953 3621 9965 3624
rect 9999 3621 10011 3655
rect 10318 3652 10324 3664
rect 10279 3624 10324 3652
rect 9953 3615 10011 3621
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10704 3661 10732 3692
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 12250 3720 12256 3732
rect 10827 3692 12256 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 10689 3655 10747 3661
rect 10689 3621 10701 3655
rect 10735 3621 10747 3655
rect 11422 3652 11428 3664
rect 11383 3624 11428 3652
rect 10689 3615 10747 3621
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 11606 3652 11612 3664
rect 11567 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 12710 3652 12716 3664
rect 11716 3624 12716 3652
rect 7392 3556 8064 3584
rect 8205 3587 8263 3593
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6328 3488 6469 3516
rect 6328 3476 6334 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 7392 3516 7420 3556
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8251 3556 8708 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8680 3528 8708 3556
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10836 3556 11069 3584
rect 10836 3544 10842 3556
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11716 3584 11744 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 11057 3547 11115 3553
rect 11164 3556 11744 3584
rect 7834 3516 7840 3528
rect 6457 3479 6515 3485
rect 6932 3488 7420 3516
rect 7795 3488 7840 3516
rect 6089 3451 6147 3457
rect 6089 3417 6101 3451
rect 6135 3448 6147 3451
rect 6932 3448 6960 3488
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 7984 3488 8029 3516
rect 7984 3476 7990 3488
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8168 3488 8493 3516
rect 8168 3476 8174 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9401 3519 9459 3525
rect 8987 3488 9352 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 6135 3420 6960 3448
rect 7009 3451 7067 3457
rect 6135 3417 6147 3420
rect 6089 3411 6147 3417
rect 7009 3417 7021 3451
rect 7055 3448 7067 3451
rect 9122 3448 9128 3460
rect 7055 3420 9128 3448
rect 7055 3417 7067 3420
rect 7009 3411 7067 3417
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 9324 3448 9352 3488
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9674 3516 9680 3528
rect 9447 3488 9680 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11164 3516 11192 3556
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 11848 3556 11893 3584
rect 11848 3544 11854 3556
rect 10551 3488 11192 3516
rect 11241 3519 11299 3525
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11882 3516 11888 3528
rect 11287 3488 11888 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 9766 3448 9772 3460
rect 9324 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 10137 3451 10195 3457
rect 10137 3417 10149 3451
rect 10183 3448 10195 3451
rect 11054 3448 11060 3460
rect 10183 3420 11060 3448
rect 10183 3417 10195 3420
rect 10137 3411 10195 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 11480 3420 11989 3448
rect 11480 3408 11486 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 11977 3411 12035 3417
rect 6273 3383 6331 3389
rect 6273 3380 6285 3383
rect 6012 3352 6285 3380
rect 6273 3349 6285 3352
rect 6319 3349 6331 3383
rect 6273 3343 6331 3349
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6454 3380 6460 3392
rect 6411 3352 6460 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 7282 3380 7288 3392
rect 7243 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 7432 3352 8309 3380
rect 7432 3340 7438 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 9677 3383 9735 3389
rect 8444 3352 8489 3380
rect 8444 3340 8450 3352
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 13170 3380 13176 3392
rect 9723 3352 13176 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 1104 3290 12328 3312
rect 1104 3238 2852 3290
rect 2904 3238 2916 3290
rect 2968 3238 2980 3290
rect 3032 3238 3044 3290
rect 3096 3238 6594 3290
rect 6646 3238 6658 3290
rect 6710 3238 6722 3290
rect 6774 3238 6786 3290
rect 6838 3238 10335 3290
rect 10387 3238 10399 3290
rect 10451 3238 10463 3290
rect 10515 3238 10527 3290
rect 10579 3238 12328 3290
rect 1104 3216 12328 3238
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 3234 3176 3240 3188
rect 2731 3148 3240 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3878 3176 3884 3188
rect 3839 3148 3884 3176
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4154 3176 4160 3188
rect 3988 3148 4160 3176
rect 753 3111 811 3117
rect 753 3077 765 3111
rect 799 3108 811 3111
rect 1854 3108 1860 3120
rect 799 3080 1860 3108
rect 799 3077 811 3080
rect 753 3071 811 3077
rect 1854 3068 1860 3080
rect 1912 3068 1918 3120
rect 2038 3068 2044 3120
rect 2096 3108 2102 3120
rect 2774 3108 2780 3120
rect 2096 3080 2780 3108
rect 2096 3068 2102 3080
rect 2774 3068 2780 3080
rect 2832 3108 2838 3120
rect 3605 3111 3663 3117
rect 2832 3080 3280 3108
rect 2832 3068 2838 3080
rect 661 3043 719 3049
rect 661 3009 673 3043
rect 707 3040 719 3043
rect 1486 3040 1492 3052
rect 707 3012 1492 3040
rect 707 3009 719 3012
rect 661 3003 719 3009
rect 1486 3000 1492 3012
rect 1544 3000 1550 3052
rect 3050 3040 3056 3052
rect 2746 3012 3056 3040
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2130 2972 2136 2984
rect 2091 2944 2136 2972
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 2746 2972 2774 3012
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3252 3049 3280 3080
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 3988 3108 4016 3148
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 7374 3176 7380 3188
rect 6144 3148 7380 3176
rect 6144 3136 6150 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7558 3136 7564 3188
rect 7616 3136 7622 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 7892 3148 8953 3176
rect 7892 3136 7898 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 8941 3139 8999 3145
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 9456 3148 9781 3176
rect 9456 3136 9462 3148
rect 9769 3145 9781 3148
rect 9815 3145 9827 3179
rect 9769 3139 9827 3145
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 12342 3176 12348 3188
rect 10183 3148 12348 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 3651 3080 4016 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 6457 3111 6515 3117
rect 4120 3080 4476 3108
rect 4120 3068 4126 3080
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4154 3040 4160 3052
rect 3835 3012 4160 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4448 3049 4476 3080
rect 6457 3077 6469 3111
rect 6503 3108 6515 3111
rect 7190 3108 7196 3120
rect 6503 3080 7196 3108
rect 6503 3077 6515 3080
rect 6457 3071 6515 3077
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4433 3003 4491 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6420 3012 6929 3040
rect 6420 3000 6426 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 7282 3040 7288 3052
rect 7147 3012 7288 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 3142 2972 3148 2984
rect 2639 2944 2774 2972
rect 3103 2944 3148 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3568 2944 3613 2972
rect 3568 2932 3574 2944
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 1486 2904 1492 2916
rect 624 2876 1492 2904
rect 624 2864 630 2876
rect 1486 2864 1492 2876
rect 1544 2864 1550 2916
rect 3053 2907 3111 2913
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 3418 2904 3424 2916
rect 3099 2876 3424 2904
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 3418 2864 3424 2876
rect 3476 2864 3482 2916
rect 290 2796 296 2848
rect 348 2836 354 2848
rect 1854 2836 1860 2848
rect 348 2808 1860 2836
rect 348 2796 354 2808
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3712 2836 3740 3000
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 4816 2972 4844 3000
rect 5074 2981 5080 2984
rect 5068 2972 5080 2981
rect 3936 2944 4844 2972
rect 5035 2944 5080 2972
rect 3936 2932 3942 2944
rect 5068 2935 5080 2944
rect 5074 2932 5080 2935
rect 5132 2932 5138 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 7190 2972 7196 2984
rect 6871 2944 7196 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7576 2981 7604 3136
rect 10597 3111 10655 3117
rect 10597 3077 10609 3111
rect 10643 3108 10655 3111
rect 11974 3108 11980 3120
rect 10643 3080 11980 3108
rect 10643 3077 10655 3080
rect 10597 3071 10655 3077
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9490 3040 9496 3052
rect 9355 3012 9496 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11606 3040 11612 3052
rect 11011 3012 11612 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 11848 3012 12020 3040
rect 11848 3000 11854 3012
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7650 2972 7656 2984
rect 7607 2944 7656 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 4246 2904 4252 2916
rect 4207 2876 4252 2904
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 4764 2876 7420 2904
rect 4764 2864 4770 2876
rect 7392 2848 7420 2876
rect 3568 2808 3740 2836
rect 3789 2839 3847 2845
rect 3568 2796 3574 2808
rect 3789 2805 3801 2839
rect 3835 2836 3847 2839
rect 4154 2836 4160 2848
rect 3835 2808 4160 2836
rect 3835 2805 3847 2808
rect 3789 2799 3847 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 5442 2836 5448 2848
rect 4387 2808 5448 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 5442 2796 5448 2808
rect 5500 2836 5506 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5500 2808 6193 2836
rect 5500 2796 5506 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6181 2799 6239 2805
rect 7374 2796 7380 2848
rect 7432 2796 7438 2848
rect 7484 2836 7512 2935
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7828 2975 7886 2981
rect 7828 2941 7840 2975
rect 7874 2972 7886 2975
rect 8386 2972 8392 2984
rect 7874 2944 8392 2972
rect 7874 2941 7886 2944
rect 7828 2935 7886 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9122 2972 9128 2984
rect 9083 2944 9128 2972
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9916 2944 10057 2972
rect 9916 2932 9922 2944
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10744 2944 10793 2972
rect 10744 2932 10750 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11992 2981 12020 3012
rect 11977 2975 12035 2981
rect 11112 2944 11284 2972
rect 11112 2932 11118 2944
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 9493 2907 9551 2913
rect 9493 2904 9505 2907
rect 8720 2876 9505 2904
rect 8720 2864 8726 2876
rect 9493 2873 9505 2876
rect 9539 2873 9551 2907
rect 10396 2907 10454 2913
rect 10396 2904 10408 2907
rect 9493 2867 9551 2873
rect 10336 2876 10408 2904
rect 8938 2836 8944 2848
rect 7484 2808 8944 2836
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 9456 2808 9597 2836
rect 9456 2796 9462 2808
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 10336 2836 10364 2876
rect 10396 2873 10408 2876
rect 10442 2873 10454 2907
rect 10396 2867 10454 2873
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11149 2907 11207 2913
rect 11149 2904 11161 2907
rect 11020 2876 11161 2904
rect 11020 2864 11026 2876
rect 11149 2873 11161 2876
rect 11195 2873 11207 2907
rect 11256 2904 11284 2944
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 11793 2907 11851 2913
rect 11256 2876 11744 2904
rect 11149 2867 11207 2873
rect 9815 2808 10364 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 11112 2808 11253 2836
rect 11112 2796 11118 2808
rect 11241 2805 11253 2808
rect 11287 2805 11299 2839
rect 11716 2836 11744 2876
rect 11793 2873 11805 2907
rect 11839 2904 11851 2907
rect 12158 2904 12164 2916
rect 11839 2876 12164 2904
rect 11839 2873 11851 2876
rect 11793 2867 11851 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12986 2836 12992 2848
rect 11716 2808 12992 2836
rect 11241 2799 11299 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 1104 2746 12328 2768
rect 1104 2694 4723 2746
rect 4775 2694 4787 2746
rect 4839 2694 4851 2746
rect 4903 2694 4915 2746
rect 4967 2694 8464 2746
rect 8516 2694 8528 2746
rect 8580 2694 8592 2746
rect 8644 2694 8656 2746
rect 8708 2694 12328 2746
rect 1104 2672 12328 2694
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4062 2632 4068 2644
rect 3988 2604 4068 2632
rect 3988 2564 4016 2604
rect 4062 2592 4068 2604
rect 4120 2632 4126 2644
rect 4120 2604 4476 2632
rect 4120 2592 4126 2604
rect 4154 2573 4160 2576
rect 4148 2564 4160 2573
rect 3344 2536 4016 2564
rect 4115 2536 4160 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2130 2496 2136 2508
rect 2091 2468 2136 2496
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 2774 2496 2780 2508
rect 2731 2468 2780 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 2792 2428 2820 2456
rect 3344 2428 3372 2536
rect 4148 2527 4160 2536
rect 4154 2524 4160 2527
rect 4212 2524 4218 2576
rect 4448 2564 4476 2604
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5224 2604 5365 2632
rect 5224 2592 5230 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 5353 2595 5411 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 6380 2604 7941 2632
rect 6380 2564 6408 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8812 2604 8953 2632
rect 8812 2592 8818 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9140 2604 9536 2632
rect 4448 2536 5396 2564
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3878 2496 3884 2508
rect 3467 2468 3740 2496
rect 3839 2468 3884 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2792 2400 3525 2428
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3712 2428 3740 2468
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4522 2496 4528 2508
rect 3988 2468 4528 2496
rect 3988 2428 4016 2468
rect 4522 2456 4528 2468
rect 4580 2496 4586 2508
rect 4580 2468 5304 2496
rect 4580 2456 4586 2468
rect 3712 2400 4016 2428
rect 3513 2391 3571 2397
rect 2777 2363 2835 2369
rect 2777 2329 2789 2363
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 3602 2360 3608 2372
rect 3007 2332 3608 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 2792 2292 2820 2323
rect 3602 2320 3608 2332
rect 3660 2320 3666 2372
rect 5276 2369 5304 2468
rect 5368 2428 5396 2536
rect 6196 2536 6408 2564
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 6196 2505 6224 2536
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 6794 2567 6852 2573
rect 6794 2564 6806 2567
rect 6512 2536 6806 2564
rect 6512 2524 6518 2536
rect 6794 2533 6806 2536
rect 6840 2533 6852 2567
rect 6794 2527 6852 2533
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 7834 2564 7840 2576
rect 6972 2536 7840 2564
rect 6972 2524 6978 2536
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8386 2564 8392 2576
rect 8347 2536 8392 2564
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 8481 2567 8539 2573
rect 8481 2533 8493 2567
rect 8527 2564 8539 2567
rect 9140 2564 9168 2604
rect 8527 2536 9168 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 9309 2567 9367 2573
rect 9309 2564 9321 2567
rect 9272 2536 9321 2564
rect 9272 2524 9278 2536
rect 9309 2533 9321 2536
rect 9355 2533 9367 2567
rect 9508 2564 9536 2604
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 9640 2604 10149 2632
rect 9640 2592 9646 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10689 2567 10747 2573
rect 9508 2536 9996 2564
rect 9309 2527 9367 2533
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5500 2468 5733 2496
rect 5500 2456 5506 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 5859 2468 6193 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 7650 2496 7656 2508
rect 6595 2468 7656 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5368 2400 6009 2428
rect 5261 2363 5319 2369
rect 5261 2329 5273 2363
rect 5307 2329 5319 2363
rect 5261 2323 5319 2329
rect 5074 2292 5080 2304
rect 2792 2264 5080 2292
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5828 2292 5856 2400
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 6380 2360 6408 2459
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 8849 2499 8907 2505
rect 8849 2496 8861 2499
rect 8036 2468 8861 2496
rect 8036 2369 8064 2468
rect 8849 2465 8861 2468
rect 8895 2465 8907 2499
rect 8849 2459 8907 2465
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 9968 2505 9996 2536
rect 10689 2533 10701 2567
rect 10735 2564 10747 2567
rect 10962 2564 10968 2576
rect 10735 2536 10968 2564
rect 10735 2533 10747 2536
rect 10689 2527 10747 2533
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 11057 2567 11115 2573
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 11146 2564 11152 2576
rect 11103 2536 11152 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11425 2567 11483 2573
rect 11425 2533 11437 2567
rect 11471 2564 11483 2567
rect 11514 2564 11520 2576
rect 11471 2536 11520 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 8996 2468 9689 2496
rect 8996 2456 9002 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10042 2496 10048 2508
rect 9999 2468 10048 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 5960 2332 6408 2360
rect 8021 2363 8079 2369
rect 5960 2320 5966 2332
rect 8021 2329 8033 2363
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 7282 2292 7288 2304
rect 5828 2264 7288 2292
rect 7282 2252 7288 2264
rect 7340 2292 7346 2304
rect 8588 2292 8616 2391
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 10152 2428 10180 2459
rect 10226 2456 10232 2508
rect 10284 2456 10290 2508
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 12434 2496 12440 2508
rect 10367 2468 12440 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 9364 2400 10180 2428
rect 9364 2388 9370 2400
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 10244 2360 10272 2456
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 10836 2400 11621 2428
rect 10836 2388 10842 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 10100 2332 10272 2360
rect 10505 2363 10563 2369
rect 10100 2320 10106 2332
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 10962 2360 10968 2372
rect 10551 2332 10968 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 7340 2264 8616 2292
rect 7340 2252 7346 2264
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9180 2264 9413 2292
rect 9180 2252 9186 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9640 2264 9781 2292
rect 9640 2252 9646 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10686 2252 10692 2304
rect 10744 2292 10750 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10744 2264 10793 2292
rect 10744 2252 10750 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 10928 2264 11161 2292
rect 10928 2252 10934 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 1104 2202 12328 2224
rect 1104 2150 2852 2202
rect 2904 2150 2916 2202
rect 2968 2150 2980 2202
rect 3032 2150 3044 2202
rect 3096 2150 6594 2202
rect 6646 2150 6658 2202
rect 6710 2150 6722 2202
rect 6774 2150 6786 2202
rect 6838 2150 10335 2202
rect 10387 2150 10399 2202
rect 10451 2150 10463 2202
rect 10515 2150 10527 2202
rect 10579 2150 12328 2202
rect 1104 2128 12328 2150
rect 845 2091 903 2097
rect 845 2057 857 2091
rect 891 2088 903 2091
rect 5442 2088 5448 2100
rect 891 2060 5448 2088
rect 891 2057 903 2060
rect 845 2051 903 2057
rect 5442 2048 5448 2060
rect 5500 2048 5506 2100
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 5718 2020 5724 2032
rect 4764 1992 5724 2020
rect 4764 1980 4770 1992
rect 5718 1980 5724 1992
rect 5776 1980 5782 2032
rect 937 1955 995 1961
rect 937 1921 949 1955
rect 983 1952 995 1955
rect 4154 1952 4160 1964
rect 983 1924 4160 1952
rect 983 1921 995 1924
rect 937 1915 995 1921
rect 4154 1912 4160 1924
rect 4212 1912 4218 1964
rect 753 1887 811 1893
rect 753 1853 765 1887
rect 799 1884 811 1887
rect 5902 1884 5908 1896
rect 799 1856 5908 1884
rect 799 1853 811 1856
rect 753 1847 811 1853
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 661 1819 719 1825
rect 661 1785 673 1819
rect 707 1816 719 1819
rect 6086 1816 6092 1828
rect 707 1788 6092 1816
rect 707 1785 719 1788
rect 661 1779 719 1785
rect 6086 1776 6092 1788
rect 6144 1776 6150 1828
rect 3878 1504 3884 1556
rect 3936 1544 3942 1556
rect 5166 1544 5172 1556
rect 3936 1516 5172 1544
rect 3936 1504 3942 1516
rect 5166 1504 5172 1516
rect 5224 1504 5230 1556
rect 3050 1436 3056 1488
rect 3108 1476 3114 1488
rect 3786 1476 3792 1488
rect 3108 1448 3792 1476
rect 3108 1436 3114 1448
rect 3786 1436 3792 1448
rect 3844 1436 3850 1488
rect 2498 1368 2504 1420
rect 2556 1408 2562 1420
rect 2682 1408 2688 1420
rect 2556 1380 2688 1408
rect 2556 1368 2562 1380
rect 2682 1368 2688 1380
rect 2740 1368 2746 1420
rect 5166 1368 5172 1420
rect 5224 1408 5230 1420
rect 5350 1408 5356 1420
rect 5224 1380 5356 1408
rect 5224 1368 5230 1380
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 6546 1408 6552 1420
rect 6052 1380 6552 1408
rect 6052 1368 6058 1380
rect 6546 1368 6552 1380
rect 6604 1368 6610 1420
rect 9306 1368 9312 1420
rect 9364 1408 9370 1420
rect 9582 1408 9588 1420
rect 9364 1380 9588 1408
rect 9364 1368 9370 1380
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
rect 5534 1300 5540 1352
rect 5592 1340 5598 1352
rect 6270 1340 6276 1352
rect 5592 1312 6276 1340
rect 5592 1300 5598 1312
rect 6270 1300 6276 1312
rect 6328 1300 6334 1352
rect 10042 1300 10048 1352
rect 10100 1340 10106 1352
rect 10318 1340 10324 1352
rect 10100 1312 10324 1340
rect 10100 1300 10106 1312
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
rect 8938 1164 8944 1216
rect 8996 1204 9002 1216
rect 10410 1204 10416 1216
rect 8996 1176 10416 1204
rect 8996 1164 9002 1176
rect 10410 1164 10416 1176
rect 10468 1164 10474 1216
rect 10686 1028 10692 1080
rect 10744 1068 10750 1080
rect 10870 1068 10876 1080
rect 10744 1040 10876 1068
rect 10744 1028 10750 1040
rect 10870 1028 10876 1040
rect 10928 1028 10934 1080
rect 4154 960 4160 1012
rect 4212 1000 4218 1012
rect 5350 1000 5356 1012
rect 4212 972 5356 1000
rect 4212 960 4218 972
rect 5350 960 5356 972
rect 5408 960 5414 1012
<< via1 >>
rect 572 13404 624 13456
rect 9036 13404 9088 13456
rect 664 13336 716 13388
rect 7288 13336 7340 13388
rect 1216 13268 1268 13320
rect 6276 13268 6328 13320
rect 1124 13200 1176 13252
rect 5540 13200 5592 13252
rect 2688 13132 2740 13184
rect 7932 13132 7984 13184
rect 2852 13030 2904 13082
rect 2916 13030 2968 13082
rect 2980 13030 3032 13082
rect 3044 13030 3096 13082
rect 6594 13030 6646 13082
rect 6658 13030 6710 13082
rect 6722 13030 6774 13082
rect 6786 13030 6838 13082
rect 10335 13030 10387 13082
rect 10399 13030 10451 13082
rect 10463 13030 10515 13082
rect 10527 13030 10579 13082
rect 940 12928 992 12980
rect 756 12860 808 12912
rect 1308 12792 1360 12844
rect 1584 12588 1636 12640
rect 5172 12928 5224 12980
rect 6920 12928 6972 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 8024 12928 8076 12980
rect 4528 12792 4580 12844
rect 5264 12792 5316 12844
rect 4620 12767 4672 12776
rect 1860 12656 1912 12708
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5080 12724 5132 12776
rect 5172 12724 5224 12776
rect 6644 12792 6696 12844
rect 8208 12860 8260 12912
rect 8300 12860 8352 12912
rect 9680 12928 9732 12980
rect 11152 12928 11204 12980
rect 7932 12792 7984 12844
rect 12624 12860 12676 12912
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 6276 12724 6328 12776
rect 7196 12767 7248 12776
rect 3424 12656 3476 12708
rect 2044 12588 2096 12640
rect 2596 12588 2648 12640
rect 3240 12588 3292 12640
rect 4252 12588 4304 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 6184 12656 6236 12708
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7288 12724 7340 12776
rect 8392 12724 8444 12776
rect 8760 12767 8812 12776
rect 8208 12656 8260 12708
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9128 12724 9180 12776
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10968 12724 11020 12776
rect 8944 12656 8996 12708
rect 6644 12588 6696 12640
rect 9312 12588 9364 12640
rect 11152 12656 11204 12708
rect 11612 12656 11664 12708
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 4723 12486 4775 12538
rect 4787 12486 4839 12538
rect 4851 12486 4903 12538
rect 4915 12486 4967 12538
rect 8464 12486 8516 12538
rect 8528 12486 8580 12538
rect 8592 12486 8644 12538
rect 8656 12486 8708 12538
rect 5080 12384 5132 12436
rect 5632 12384 5684 12436
rect 6368 12384 6420 12436
rect 8208 12427 8260 12436
rect 3700 12359 3752 12368
rect 3700 12325 3709 12359
rect 3709 12325 3743 12359
rect 3743 12325 3752 12359
rect 3700 12316 3752 12325
rect 4252 12316 4304 12368
rect 4712 12316 4764 12368
rect 5172 12316 5224 12368
rect 1676 12291 1728 12300
rect 1676 12257 1710 12291
rect 1710 12257 1728 12291
rect 1676 12248 1728 12257
rect 2412 12248 2464 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 4436 12248 4488 12300
rect 4988 12248 5040 12300
rect 3700 12180 3752 12232
rect 2136 12044 2188 12096
rect 3608 12044 3660 12096
rect 5908 12248 5960 12300
rect 7748 12316 7800 12368
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 8760 12384 8812 12436
rect 8944 12384 8996 12436
rect 9220 12384 9272 12436
rect 11612 12384 11664 12436
rect 9772 12316 9824 12368
rect 6920 12248 6972 12300
rect 8944 12248 8996 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 9404 12180 9456 12232
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 9956 12180 10008 12232
rect 6368 12112 6420 12164
rect 8116 12044 8168 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 10784 12044 10836 12096
rect 2852 11942 2904 11994
rect 2916 11942 2968 11994
rect 2980 11942 3032 11994
rect 3044 11942 3096 11994
rect 6594 11942 6646 11994
rect 6658 11942 6710 11994
rect 6722 11942 6774 11994
rect 6786 11942 6838 11994
rect 10335 11942 10387 11994
rect 10399 11942 10451 11994
rect 10463 11942 10515 11994
rect 10527 11942 10579 11994
rect 112 11840 164 11892
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2412 11772 2464 11824
rect 4620 11840 4672 11892
rect 5908 11840 5960 11892
rect 6920 11840 6972 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9496 11840 9548 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 11244 11883 11296 11892
rect 10232 11840 10284 11849
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 1400 11500 1452 11552
rect 2044 11500 2096 11552
rect 2780 11611 2832 11620
rect 2780 11577 2814 11611
rect 2814 11577 2832 11611
rect 2780 11568 2832 11577
rect 3608 11568 3660 11620
rect 5356 11772 5408 11824
rect 5448 11772 5500 11824
rect 8944 11772 8996 11824
rect 4528 11704 4580 11756
rect 5080 11704 5132 11756
rect 5540 11704 5592 11756
rect 5816 11704 5868 11756
rect 4436 11679 4488 11688
rect 4436 11645 4445 11679
rect 4445 11645 4479 11679
rect 4479 11645 4488 11679
rect 4436 11636 4488 11645
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6368 11704 6420 11756
rect 5632 11568 5684 11620
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 7196 11636 7248 11688
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 8300 11636 8352 11688
rect 9128 11636 9180 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 10508 11704 10560 11756
rect 10416 11679 10468 11688
rect 3332 11500 3384 11552
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 5908 11500 5960 11552
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 8208 11568 8260 11620
rect 9588 11568 9640 11620
rect 10416 11645 10425 11679
rect 10425 11645 10459 11679
rect 10459 11645 10468 11679
rect 10416 11636 10468 11645
rect 10784 11704 10836 11756
rect 11152 11679 11204 11688
rect 7288 11500 7340 11552
rect 7564 11500 7616 11552
rect 9956 11500 10008 11552
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 11520 11636 11572 11688
rect 10968 11543 11020 11552
rect 10968 11509 10977 11543
rect 10977 11509 11011 11543
rect 11011 11509 11020 11543
rect 10968 11500 11020 11509
rect 4723 11398 4775 11450
rect 4787 11398 4839 11450
rect 4851 11398 4903 11450
rect 4915 11398 4967 11450
rect 8464 11398 8516 11450
rect 8528 11398 8580 11450
rect 8592 11398 8644 11450
rect 8656 11398 8708 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2228 11296 2280 11348
rect 2044 11228 2096 11280
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 3056 11339 3108 11348
rect 2780 11296 2832 11305
rect 3056 11305 3065 11339
rect 3065 11305 3099 11339
rect 3099 11305 3108 11339
rect 3056 11296 3108 11305
rect 5632 11296 5684 11348
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 4252 11228 4304 11280
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 3884 11203 3936 11212
rect 572 11024 624 11076
rect 848 11024 900 11076
rect 2504 11024 2556 11076
rect 3884 11169 3893 11203
rect 3893 11169 3927 11203
rect 3927 11169 3936 11203
rect 3884 11160 3936 11169
rect 4528 11160 4580 11212
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4344 11092 4396 11144
rect 4804 11160 4856 11212
rect 5264 11160 5316 11212
rect 5448 11160 5500 11212
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6184 11296 6236 11348
rect 6276 11228 6328 11280
rect 6552 11296 6604 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 9680 11296 9732 11348
rect 10048 11296 10100 11348
rect 10324 11296 10376 11348
rect 8300 11228 8352 11280
rect 8484 11271 8536 11280
rect 8484 11237 8493 11271
rect 8493 11237 8527 11271
rect 8527 11237 8536 11271
rect 8484 11228 8536 11237
rect 8944 11228 8996 11280
rect 6920 11160 6972 11212
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 9036 11160 9088 11212
rect 10416 11228 10468 11280
rect 10508 11228 10560 11280
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10324 11160 10376 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 4436 11024 4488 11076
rect 4068 10956 4120 11008
rect 4804 10956 4856 11008
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 5172 10956 5224 11008
rect 6000 10956 6052 11008
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 9864 11024 9916 11076
rect 10048 11024 10100 11076
rect 10876 11160 10928 11212
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 10692 11024 10744 11076
rect 10784 10956 10836 11008
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 2852 10854 2904 10906
rect 2916 10854 2968 10906
rect 2980 10854 3032 10906
rect 3044 10854 3096 10906
rect 6594 10854 6646 10906
rect 6658 10854 6710 10906
rect 6722 10854 6774 10906
rect 6786 10854 6838 10906
rect 10335 10854 10387 10906
rect 10399 10854 10451 10906
rect 10463 10854 10515 10906
rect 10527 10854 10579 10906
rect 1768 10752 1820 10804
rect 3424 10752 3476 10804
rect 3516 10752 3568 10804
rect 5540 10795 5592 10804
rect 2780 10684 2832 10736
rect 3240 10684 3292 10736
rect 3792 10684 3844 10736
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 2228 10616 2280 10668
rect 2412 10616 2464 10668
rect 3332 10616 3384 10668
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 6000 10684 6052 10736
rect 6368 10752 6420 10804
rect 7012 10752 7064 10804
rect 2964 10480 3016 10532
rect 3332 10480 3384 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3240 10412 3292 10464
rect 3608 10480 3660 10532
rect 4243 10523 4295 10532
rect 4243 10489 4252 10523
rect 4252 10489 4286 10523
rect 4286 10489 4295 10523
rect 4243 10480 4295 10489
rect 5540 10548 5592 10600
rect 8208 10752 8260 10804
rect 8484 10752 8536 10804
rect 10876 10752 10928 10804
rect 11244 10752 11296 10804
rect 9680 10684 9732 10736
rect 9864 10684 9916 10736
rect 3976 10412 4028 10464
rect 4620 10412 4672 10464
rect 5540 10412 5592 10464
rect 6184 10548 6236 10600
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 6552 10480 6604 10532
rect 8852 10548 8904 10600
rect 6000 10412 6052 10464
rect 6184 10412 6236 10464
rect 6368 10412 6420 10464
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 8300 10480 8352 10532
rect 9588 10480 9640 10532
rect 9772 10480 9824 10532
rect 9036 10412 9088 10464
rect 9680 10412 9732 10464
rect 10232 10548 10284 10600
rect 10784 10480 10836 10532
rect 11152 10548 11204 10600
rect 11244 10480 11296 10532
rect 10508 10412 10560 10464
rect 4723 10310 4775 10362
rect 4787 10310 4839 10362
rect 4851 10310 4903 10362
rect 4915 10310 4967 10362
rect 8464 10310 8516 10362
rect 8528 10310 8580 10362
rect 8592 10310 8644 10362
rect 8656 10310 8708 10362
rect 2872 10208 2924 10260
rect 3148 10140 3200 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 2412 10072 2464 10124
rect 3424 10115 3476 10124
rect 3424 10081 3433 10115
rect 3433 10081 3467 10115
rect 3467 10081 3476 10115
rect 3424 10072 3476 10081
rect 4160 10208 4212 10260
rect 9772 10208 9824 10260
rect 4896 10140 4948 10192
rect 5816 10183 5868 10192
rect 5816 10149 5850 10183
rect 5850 10149 5868 10183
rect 5816 10140 5868 10149
rect 7840 10140 7892 10192
rect 3884 10072 3936 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 4160 10072 4212 10124
rect 4436 10072 4488 10124
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 4712 10072 4764 10124
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5540 10115 5592 10124
rect 1768 10004 1820 10013
rect 1492 9868 1544 9920
rect 4896 10004 4948 10056
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 2964 9936 3016 9988
rect 4252 9936 4304 9988
rect 3516 9868 3568 9920
rect 3976 9868 4028 9920
rect 4712 9868 4764 9920
rect 5080 9868 5132 9920
rect 5540 9868 5592 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 7380 9868 7432 9920
rect 8208 10072 8260 10124
rect 8944 10115 8996 10124
rect 8392 10004 8444 10056
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9404 10072 9456 10124
rect 8852 10004 8904 10056
rect 8668 9936 8720 9988
rect 9128 9868 9180 9920
rect 9864 10140 9916 10192
rect 10692 10208 10744 10260
rect 10048 10140 10100 10192
rect 10324 10140 10376 10192
rect 11336 10140 11388 10192
rect 10876 10115 10928 10124
rect 10876 10081 10910 10115
rect 10910 10081 10928 10115
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 9864 10004 9916 10056
rect 10876 10072 10928 10081
rect 10232 9936 10284 9988
rect 9956 9868 10008 9920
rect 2852 9766 2904 9818
rect 2916 9766 2968 9818
rect 2980 9766 3032 9818
rect 3044 9766 3096 9818
rect 6594 9766 6646 9818
rect 6658 9766 6710 9818
rect 6722 9766 6774 9818
rect 6786 9766 6838 9818
rect 10335 9766 10387 9818
rect 10399 9766 10451 9818
rect 10463 9766 10515 9818
rect 10527 9766 10579 9818
rect 1400 9664 1452 9716
rect 2780 9596 2832 9648
rect 3424 9639 3476 9648
rect 3424 9605 3433 9639
rect 3433 9605 3467 9639
rect 3467 9605 3476 9639
rect 3424 9596 3476 9605
rect 4068 9664 4120 9716
rect 4712 9664 4764 9716
rect 4988 9664 5040 9716
rect 1032 9528 1084 9580
rect 2228 9528 2280 9580
rect 2688 9460 2740 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 3424 9460 3476 9512
rect 5816 9664 5868 9716
rect 6460 9664 6512 9716
rect 7104 9664 7156 9716
rect 8944 9664 8996 9716
rect 10232 9664 10284 9716
rect 10876 9664 10928 9716
rect 6368 9596 6420 9648
rect 4620 9460 4672 9512
rect 2780 9324 2832 9376
rect 3976 9324 4028 9376
rect 4804 9392 4856 9444
rect 5080 9460 5132 9512
rect 5356 9460 5408 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 6920 9528 6972 9580
rect 8392 9596 8444 9648
rect 9220 9596 9272 9648
rect 5448 9460 5500 9469
rect 5540 9392 5592 9444
rect 6184 9503 6236 9512
rect 6184 9469 6201 9503
rect 6201 9469 6235 9503
rect 6235 9469 6236 9503
rect 6184 9460 6236 9469
rect 6368 9460 6420 9512
rect 6644 9460 6696 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7196 9392 7248 9444
rect 7380 9503 7432 9512
rect 7380 9469 7414 9503
rect 7414 9469 7432 9503
rect 9956 9528 10008 9580
rect 7380 9460 7432 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 10784 9460 10836 9512
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 12072 9460 12124 9512
rect 7656 9324 7708 9376
rect 9404 9324 9456 9376
rect 9680 9324 9732 9376
rect 9956 9435 10008 9444
rect 9956 9401 9965 9435
rect 9965 9401 9999 9435
rect 9999 9401 10008 9435
rect 10140 9435 10192 9444
rect 9956 9392 10008 9401
rect 10140 9401 10149 9435
rect 10149 9401 10183 9435
rect 10183 9401 10192 9435
rect 10140 9392 10192 9401
rect 10692 9392 10744 9444
rect 10876 9324 10928 9376
rect 4723 9222 4775 9274
rect 4787 9222 4839 9274
rect 4851 9222 4903 9274
rect 4915 9222 4967 9274
rect 8464 9222 8516 9274
rect 8528 9222 8580 9274
rect 8592 9222 8644 9274
rect 8656 9222 8708 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 4068 9120 4120 9172
rect 6092 9120 6144 9172
rect 6920 9120 6972 9172
rect 8300 9120 8352 9172
rect 1768 9052 1820 9104
rect 2504 9052 2556 9104
rect 3240 9052 3292 9104
rect 3976 9052 4028 9104
rect 4620 9052 4672 9104
rect 4804 9052 4856 9104
rect 6276 9052 6328 9104
rect 9404 9120 9456 9172
rect 1676 9027 1728 9036
rect 1676 8993 1710 9027
rect 1710 8993 1728 9027
rect 1676 8984 1728 8993
rect 2228 8984 2280 9036
rect 2412 8916 2464 8968
rect 4712 8984 4764 9036
rect 6920 8984 6972 9036
rect 7196 9027 7248 9036
rect 7196 8993 7230 9027
rect 7230 8993 7248 9027
rect 7196 8984 7248 8993
rect 3240 8916 3292 8968
rect 2504 8780 2556 8832
rect 3332 8780 3384 8832
rect 5080 8916 5132 8968
rect 6644 8848 6696 8900
rect 4068 8780 4120 8832
rect 4804 8780 4856 8832
rect 6276 8780 6328 8832
rect 6920 8848 6972 8900
rect 7196 8848 7248 8900
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 8944 8984 8996 9036
rect 10140 9027 10192 9036
rect 9220 8916 9272 8968
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 11152 8984 11204 9036
rect 9956 8848 10008 8900
rect 8668 8780 8720 8832
rect 9036 8780 9088 8832
rect 11244 8916 11296 8968
rect 10140 8848 10192 8900
rect 10232 8780 10284 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 11704 8780 11756 8832
rect 2852 8678 2904 8730
rect 2916 8678 2968 8730
rect 2980 8678 3032 8730
rect 3044 8678 3096 8730
rect 6594 8678 6646 8730
rect 6658 8678 6710 8730
rect 6722 8678 6774 8730
rect 6786 8678 6838 8730
rect 10335 8678 10387 8730
rect 10399 8678 10451 8730
rect 10463 8678 10515 8730
rect 10527 8678 10579 8730
rect 1400 8619 1452 8628
rect 1400 8585 1409 8619
rect 1409 8585 1443 8619
rect 1443 8585 1452 8619
rect 1400 8576 1452 8585
rect 1676 8576 1728 8628
rect 3240 8576 3292 8628
rect 7012 8576 7064 8628
rect 7196 8576 7248 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 9772 8576 9824 8628
rect 848 8372 900 8424
rect 1768 8372 1820 8424
rect 2044 8372 2096 8424
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2872 8508 2924 8560
rect 2136 8304 2188 8356
rect 2688 8304 2740 8356
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 2044 8236 2096 8245
rect 3424 8372 3476 8424
rect 5356 8508 5408 8560
rect 6184 8508 6236 8560
rect 11060 8576 11112 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 11152 8508 11204 8560
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 6460 8440 6512 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 10048 8440 10100 8492
rect 10784 8440 10836 8492
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 5540 8372 5592 8424
rect 6644 8415 6696 8424
rect 2964 8304 3016 8356
rect 3056 8304 3108 8356
rect 3976 8304 4028 8356
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7104 8372 7156 8424
rect 7748 8372 7800 8424
rect 9220 8415 9272 8424
rect 6828 8304 6880 8356
rect 8300 8304 8352 8356
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 10232 8372 10284 8424
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 3884 8236 3936 8288
rect 4436 8236 4488 8288
rect 5448 8236 5500 8288
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 4723 8134 4775 8186
rect 4787 8134 4839 8186
rect 4851 8134 4903 8186
rect 4915 8134 4967 8186
rect 8464 8134 8516 8186
rect 8528 8134 8580 8186
rect 8592 8134 8644 8186
rect 8656 8134 8708 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 2136 8032 2188 8084
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 5356 8032 5408 8084
rect 6644 8032 6696 8084
rect 7288 8032 7340 8084
rect 9956 8032 10008 8084
rect 3976 8007 4028 8016
rect 3976 7973 3985 8007
rect 3985 7973 4019 8007
rect 4019 7973 4028 8007
rect 3976 7964 4028 7973
rect 1768 7828 1820 7880
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 388 7760 440 7812
rect 1308 7760 1360 7812
rect 2688 7896 2740 7948
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 3240 7939 3292 7948
rect 2872 7896 2924 7905
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 3884 7896 3936 7948
rect 4436 7939 4488 7948
rect 3148 7760 3200 7812
rect 3240 7760 3292 7812
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 5632 7964 5684 8016
rect 6184 8007 6236 8016
rect 6184 7973 6193 8007
rect 6193 7973 6227 8007
rect 6227 7973 6236 8007
rect 6184 7964 6236 7973
rect 6000 7896 6052 7948
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6828 7964 6880 8016
rect 9404 7964 9456 8016
rect 4068 7828 4120 7880
rect 9128 7939 9180 7948
rect 6460 7828 6512 7880
rect 6276 7760 6328 7812
rect 6552 7760 6604 7812
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 10048 7964 10100 8016
rect 10692 7964 10744 8016
rect 11060 7896 11112 7948
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 8300 7828 8352 7880
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 9036 7828 9088 7880
rect 9956 7828 10008 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 8852 7760 8904 7812
rect 9680 7760 9732 7812
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 9036 7692 9088 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 10232 7692 10284 7744
rect 10968 7692 11020 7744
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 2852 7590 2904 7642
rect 2916 7590 2968 7642
rect 2980 7590 3032 7642
rect 3044 7590 3096 7642
rect 6594 7590 6646 7642
rect 6658 7590 6710 7642
rect 6722 7590 6774 7642
rect 6786 7590 6838 7642
rect 10335 7590 10387 7642
rect 10399 7590 10451 7642
rect 10463 7590 10515 7642
rect 10527 7590 10579 7642
rect 2320 7488 2372 7540
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 1492 7420 1544 7472
rect 1952 7420 2004 7472
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 1860 7284 1912 7336
rect 2412 7284 2464 7336
rect 2872 7284 2924 7336
rect 2780 7216 2832 7268
rect 3240 7488 3292 7540
rect 3424 7488 3476 7540
rect 3148 7420 3200 7472
rect 3056 7284 3108 7336
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3976 7352 4028 7404
rect 5080 7488 5132 7540
rect 5540 7488 5592 7540
rect 6460 7488 6512 7540
rect 7196 7488 7248 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 10692 7488 10744 7540
rect 4160 7284 4212 7336
rect 4712 7284 4764 7336
rect 6828 7420 6880 7472
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 9680 7420 9732 7472
rect 6000 7352 6052 7404
rect 6184 7352 6236 7404
rect 7196 7352 7248 7404
rect 9864 7352 9916 7404
rect 12440 7352 12492 7404
rect 5540 7284 5592 7336
rect 5632 7284 5684 7336
rect 8300 7327 8352 7336
rect 5264 7148 5316 7200
rect 5632 7148 5684 7200
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 9312 7284 9364 7336
rect 6000 7216 6052 7268
rect 6184 7216 6236 7268
rect 6920 7216 6972 7268
rect 7380 7216 7432 7268
rect 8668 7216 8720 7268
rect 9864 7216 9916 7268
rect 10324 7284 10376 7336
rect 10416 7284 10468 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 11244 7284 11296 7336
rect 11428 7284 11480 7336
rect 6276 7148 6328 7200
rect 6644 7148 6696 7200
rect 8116 7148 8168 7200
rect 4723 7046 4775 7098
rect 4787 7046 4839 7098
rect 4851 7046 4903 7098
rect 4915 7046 4967 7098
rect 8464 7046 8516 7098
rect 8528 7046 8580 7098
rect 8592 7046 8644 7098
rect 8656 7046 8708 7098
rect 2596 6944 2648 6996
rect 3884 6944 3936 6996
rect 1676 6851 1728 6860
rect 1676 6817 1710 6851
rect 1710 6817 1728 6851
rect 1676 6808 1728 6817
rect 2136 6808 2188 6860
rect 5540 6876 5592 6928
rect 6000 6876 6052 6928
rect 6644 6944 6696 6996
rect 8852 6987 8904 6996
rect 8852 6953 8861 6987
rect 8861 6953 8895 6987
rect 8895 6953 8904 6987
rect 8852 6944 8904 6953
rect 9128 6944 9180 6996
rect 9588 6944 9640 6996
rect 10048 6944 10100 6996
rect 10324 6944 10376 6996
rect 10876 6944 10928 6996
rect 6920 6876 6972 6928
rect 7104 6919 7156 6928
rect 7104 6885 7138 6919
rect 7138 6885 7156 6919
rect 7104 6876 7156 6885
rect 9680 6876 9732 6928
rect 2872 6715 2924 6724
rect 2872 6681 2881 6715
rect 2881 6681 2915 6715
rect 2915 6681 2924 6715
rect 2872 6672 2924 6681
rect 2596 6604 2648 6656
rect 4160 6851 4212 6860
rect 4160 6817 4194 6851
rect 4194 6817 4212 6851
rect 3608 6740 3660 6792
rect 4160 6808 4212 6817
rect 5264 6808 5316 6860
rect 5632 6851 5684 6860
rect 5632 6817 5666 6851
rect 5666 6817 5684 6851
rect 5632 6808 5684 6817
rect 6184 6808 6236 6860
rect 3884 6604 3936 6656
rect 7840 6740 7892 6792
rect 9036 6808 9088 6860
rect 9312 6740 9364 6792
rect 9864 6740 9916 6792
rect 8300 6672 8352 6724
rect 10416 6740 10468 6792
rect 11152 6740 11204 6792
rect 7196 6604 7248 6656
rect 10784 6604 10836 6656
rect 11612 6604 11664 6656
rect 2852 6502 2904 6554
rect 2916 6502 2968 6554
rect 2980 6502 3032 6554
rect 3044 6502 3096 6554
rect 6594 6502 6646 6554
rect 6658 6502 6710 6554
rect 6722 6502 6774 6554
rect 6786 6502 6838 6554
rect 10335 6502 10387 6554
rect 10399 6502 10451 6554
rect 10463 6502 10515 6554
rect 10527 6502 10579 6554
rect 1676 6400 1728 6452
rect 3424 6400 3476 6452
rect 3976 6443 4028 6452
rect 3976 6409 3985 6443
rect 3985 6409 4019 6443
rect 4019 6409 4028 6443
rect 3976 6400 4028 6409
rect 2136 6264 2188 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2412 6196 2464 6248
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 3148 6264 3200 6316
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 3240 6128 3292 6180
rect 3424 6196 3476 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 4436 6239 4488 6248
rect 3976 6128 4028 6180
rect 1676 6060 1728 6112
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 3884 6060 3936 6112
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 5540 6400 5592 6452
rect 5816 6400 5868 6452
rect 6460 6400 6512 6452
rect 7840 6400 7892 6452
rect 8116 6400 8168 6452
rect 8300 6400 8352 6452
rect 5172 6264 5224 6316
rect 6092 6332 6144 6384
rect 5264 6060 5316 6112
rect 6184 6196 6236 6248
rect 6552 6196 6604 6248
rect 6644 6196 6696 6248
rect 7196 6264 7248 6316
rect 7380 6264 7432 6316
rect 7288 6196 7340 6248
rect 7840 6196 7892 6248
rect 10048 6264 10100 6316
rect 11060 6400 11112 6452
rect 11244 6264 11296 6316
rect 8116 6128 8168 6180
rect 8944 6128 8996 6180
rect 10692 6128 10744 6180
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 7380 6060 7432 6112
rect 7932 6060 7984 6112
rect 9588 6060 9640 6112
rect 11060 6060 11112 6112
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 4723 5958 4775 6010
rect 4787 5958 4839 6010
rect 4851 5958 4903 6010
rect 4915 5958 4967 6010
rect 8464 5958 8516 6010
rect 8528 5958 8580 6010
rect 8592 5958 8644 6010
rect 8656 5958 8708 6010
rect 1400 5856 1452 5908
rect 2044 5856 2096 5908
rect 3424 5856 3476 5908
rect 6644 5856 6696 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 8116 5899 8168 5908
rect 8116 5865 8125 5899
rect 8125 5865 8159 5899
rect 8159 5865 8168 5899
rect 8116 5856 8168 5865
rect 10692 5899 10744 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 2136 5720 2188 5772
rect 2412 5720 2464 5772
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 2688 5720 2740 5772
rect 3240 5788 3292 5840
rect 3792 5788 3844 5840
rect 5448 5788 5500 5840
rect 5908 5788 5960 5840
rect 6276 5788 6328 5840
rect 6736 5788 6788 5840
rect 6920 5788 6972 5840
rect 7840 5788 7892 5840
rect 4160 5652 4212 5704
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 4896 5720 4948 5772
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 7288 5720 7340 5772
rect 8944 5831 8996 5840
rect 8944 5797 8953 5831
rect 8953 5797 8987 5831
rect 8987 5797 8996 5831
rect 8944 5788 8996 5797
rect 8300 5720 8352 5772
rect 8576 5763 8628 5772
rect 1400 5627 1452 5636
rect 1400 5593 1409 5627
rect 1409 5593 1443 5627
rect 1443 5593 1452 5627
rect 1400 5584 1452 5593
rect 3056 5584 3108 5636
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 3240 5516 3292 5568
rect 6092 5584 6144 5636
rect 6552 5584 6604 5636
rect 7656 5584 7708 5636
rect 7840 5584 7892 5636
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 9496 5720 9548 5772
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 11244 5788 11296 5840
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10784 5720 10836 5772
rect 10232 5652 10284 5704
rect 9588 5584 9640 5636
rect 5448 5516 5500 5568
rect 8300 5516 8352 5568
rect 9680 5516 9732 5568
rect 11796 5652 11848 5704
rect 10784 5584 10836 5636
rect 10876 5584 10928 5636
rect 10692 5516 10744 5568
rect 10968 5516 11020 5568
rect 2852 5414 2904 5466
rect 2916 5414 2968 5466
rect 2980 5414 3032 5466
rect 3044 5414 3096 5466
rect 6594 5414 6646 5466
rect 6658 5414 6710 5466
rect 6722 5414 6774 5466
rect 6786 5414 6838 5466
rect 10335 5414 10387 5466
rect 10399 5414 10451 5466
rect 10463 5414 10515 5466
rect 10527 5414 10579 5466
rect 2504 5312 2556 5364
rect 4344 5312 4396 5364
rect 2688 5244 2740 5296
rect 4620 5244 4672 5296
rect 4896 5244 4948 5296
rect 5356 5244 5408 5296
rect 6736 5244 6788 5296
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 2044 5108 2096 5160
rect 2412 5040 2464 5092
rect 3240 5108 3292 5160
rect 4712 5108 4764 5160
rect 6828 5108 6880 5160
rect 5080 5083 5132 5092
rect 5080 5049 5089 5083
rect 5089 5049 5123 5083
rect 5123 5049 5132 5083
rect 5080 5040 5132 5049
rect 6276 5040 6328 5092
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 9128 5312 9180 5364
rect 9864 5312 9916 5364
rect 9496 5244 9548 5296
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9680 5176 9732 5228
rect 10048 5176 10100 5228
rect 8944 5108 8996 5160
rect 10232 5108 10284 5160
rect 10692 5108 10744 5160
rect 11520 5108 11572 5160
rect 3608 4972 3660 5024
rect 4068 4972 4120 5024
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 6828 4972 6880 5024
rect 7472 4972 7524 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 7932 4972 7984 5024
rect 9128 5040 9180 5092
rect 9864 5083 9916 5092
rect 9864 5049 9873 5083
rect 9873 5049 9907 5083
rect 9907 5049 9916 5083
rect 9864 5040 9916 5049
rect 10324 5040 10376 5092
rect 13268 5040 13320 5092
rect 4723 4870 4775 4922
rect 4787 4870 4839 4922
rect 4851 4870 4903 4922
rect 4915 4870 4967 4922
rect 8464 4870 8516 4922
rect 8528 4870 8580 4922
rect 8592 4870 8644 4922
rect 8656 4870 8708 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 2504 4768 2556 4820
rect 204 4632 256 4684
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 3240 4768 3292 4820
rect 3976 4768 4028 4820
rect 4068 4768 4120 4820
rect 4160 4768 4212 4820
rect 5356 4768 5408 4820
rect 3148 4632 3200 4684
rect 3424 4632 3476 4684
rect 3792 4632 3844 4684
rect 3976 4675 4028 4684
rect 3976 4641 3985 4675
rect 3985 4641 4019 4675
rect 4019 4641 4028 4675
rect 3976 4632 4028 4641
rect 4068 4632 4120 4684
rect 4344 4632 4396 4684
rect 5632 4700 5684 4752
rect 6552 4700 6604 4752
rect 7288 4768 7340 4820
rect 7472 4768 7524 4820
rect 8208 4768 8260 4820
rect 6920 4700 6972 4752
rect 4988 4632 5040 4684
rect 6828 4632 6880 4684
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 7656 4700 7708 4752
rect 2320 4564 2372 4616
rect 3700 4564 3752 4616
rect 6920 4539 6972 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 3424 4428 3476 4480
rect 3608 4428 3660 4480
rect 4896 4428 4948 4480
rect 6920 4505 6929 4539
rect 6929 4505 6963 4539
rect 6963 4505 6972 4539
rect 6920 4496 6972 4505
rect 5448 4428 5500 4480
rect 6092 4428 6144 4480
rect 6368 4428 6420 4480
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 10232 4768 10284 4820
rect 10600 4768 10652 4820
rect 9588 4743 9640 4752
rect 9588 4709 9597 4743
rect 9597 4709 9631 4743
rect 9631 4709 9640 4743
rect 9588 4700 9640 4709
rect 10876 4700 10928 4752
rect 11336 4700 11388 4752
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 9312 4564 9364 4616
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12532 4496 12584 4548
rect 8576 4428 8628 4480
rect 8944 4428 8996 4480
rect 9496 4428 9548 4480
rect 9680 4428 9732 4480
rect 9956 4428 10008 4480
rect 12900 4428 12952 4480
rect 2852 4326 2904 4378
rect 2916 4326 2968 4378
rect 2980 4326 3032 4378
rect 3044 4326 3096 4378
rect 6594 4326 6646 4378
rect 6658 4326 6710 4378
rect 6722 4326 6774 4378
rect 6786 4326 6838 4378
rect 10335 4326 10387 4378
rect 10399 4326 10451 4378
rect 10463 4326 10515 4378
rect 10527 4326 10579 4378
rect 480 4267 532 4276
rect 480 4233 489 4267
rect 489 4233 523 4267
rect 523 4233 532 4267
rect 480 4224 532 4233
rect 2504 4224 2556 4276
rect 3424 4267 3476 4276
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 4896 4224 4948 4276
rect 5632 4224 5684 4276
rect 5816 4224 5868 4276
rect 2136 4156 2188 4208
rect 112 4088 164 4140
rect 480 4088 532 4140
rect 940 4088 992 4140
rect 1952 4088 2004 4140
rect 2504 4088 2556 4140
rect 2964 4156 3016 4208
rect 3608 4131 3660 4140
rect 3608 4097 3620 4131
rect 3620 4097 3654 4131
rect 3654 4097 3660 4131
rect 3608 4088 3660 4097
rect 1124 4020 1176 4072
rect 2136 4020 2188 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3148 4020 3200 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3700 4063 3752 4072
rect 3332 4020 3384 4029
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 3792 4020 3844 4072
rect 6092 4156 6144 4208
rect 6368 4156 6420 4208
rect 6552 4131 6604 4140
rect 112 3952 164 4004
rect 20 3884 72 3936
rect 4988 3952 5040 4004
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 4068 3884 4120 3936
rect 5540 3952 5592 4004
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7380 4224 7432 4276
rect 7288 4156 7340 4208
rect 6092 4020 6144 4072
rect 6092 3884 6144 3936
rect 8300 4088 8352 4140
rect 8852 4088 8904 4140
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7840 4020 7892 4072
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 7380 3952 7432 4004
rect 8392 4020 8444 4072
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9496 4224 9548 4276
rect 9588 4224 9640 4276
rect 12164 4224 12216 4276
rect 9312 4156 9364 4208
rect 10692 4156 10744 4208
rect 11980 4156 12032 4208
rect 12624 4088 12676 4140
rect 10048 4020 10100 4072
rect 11704 4020 11756 4072
rect 11888 4020 11940 4072
rect 10232 3952 10284 4004
rect 11244 3952 11296 4004
rect 12072 3952 12124 4004
rect 7104 3884 7156 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 9680 3884 9732 3936
rect 10048 3884 10100 3936
rect 11704 3884 11756 3936
rect 388 3816 440 3868
rect 940 3816 992 3868
rect 4723 3782 4775 3834
rect 4787 3782 4839 3834
rect 4851 3782 4903 3834
rect 4915 3782 4967 3834
rect 8464 3782 8516 3834
rect 8528 3782 8580 3834
rect 8592 3782 8644 3834
rect 8656 3782 8708 3834
rect 388 3680 440 3732
rect 3056 3680 3108 3732
rect 3240 3680 3292 3732
rect 3332 3680 3384 3732
rect 4160 3680 4212 3732
rect 3792 3612 3844 3664
rect 2964 3587 3016 3596
rect 2964 3553 2973 3587
rect 2973 3553 3007 3587
rect 3007 3553 3016 3587
rect 2964 3544 3016 3553
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 3608 3544 3660 3596
rect 3884 3587 3936 3596
rect 3884 3553 3893 3587
rect 3893 3553 3927 3587
rect 3927 3553 3936 3587
rect 3884 3544 3936 3553
rect 7288 3680 7340 3732
rect 7472 3680 7524 3732
rect 7932 3680 7984 3732
rect 9128 3680 9180 3732
rect 9404 3680 9456 3732
rect 9864 3680 9916 3732
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 4436 3476 4488 3528
rect 4160 3408 4212 3460
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 5172 3587 5224 3596
rect 4896 3544 4948 3553
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5908 3544 5960 3596
rect 2688 3340 2740 3392
rect 3516 3340 3568 3392
rect 3976 3340 4028 3392
rect 4896 3340 4948 3392
rect 5080 3340 5132 3392
rect 6092 3544 6144 3596
rect 7196 3544 7248 3596
rect 8944 3612 8996 3664
rect 9496 3612 9548 3664
rect 9772 3612 9824 3664
rect 10324 3655 10376 3664
rect 10324 3621 10333 3655
rect 10333 3621 10367 3655
rect 10367 3621 10376 3655
rect 10324 3612 10376 3621
rect 12256 3680 12308 3732
rect 11428 3655 11480 3664
rect 11428 3621 11437 3655
rect 11437 3621 11471 3655
rect 11471 3621 11480 3655
rect 11428 3612 11480 3621
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 6276 3476 6328 3528
rect 10784 3544 10836 3596
rect 12716 3612 12768 3664
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8116 3476 8168 3528
rect 8668 3476 8720 3528
rect 9128 3408 9180 3460
rect 9680 3476 9732 3528
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 11888 3476 11940 3528
rect 9772 3408 9824 3460
rect 11060 3408 11112 3460
rect 11428 3408 11480 3460
rect 6460 3340 6512 3392
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7380 3340 7432 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 13176 3340 13228 3392
rect 2852 3238 2904 3290
rect 2916 3238 2968 3290
rect 2980 3238 3032 3290
rect 3044 3238 3096 3290
rect 6594 3238 6646 3290
rect 6658 3238 6710 3290
rect 6722 3238 6774 3290
rect 6786 3238 6838 3290
rect 10335 3238 10387 3290
rect 10399 3238 10451 3290
rect 10463 3238 10515 3290
rect 10527 3238 10579 3290
rect 3240 3136 3292 3188
rect 3884 3179 3936 3188
rect 3884 3145 3893 3179
rect 3893 3145 3927 3179
rect 3927 3145 3936 3179
rect 3884 3136 3936 3145
rect 1860 3068 1912 3120
rect 2044 3068 2096 3120
rect 2780 3068 2832 3120
rect 1492 3000 1544 3052
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 3056 3000 3108 3052
rect 4160 3136 4212 3188
rect 6092 3136 6144 3188
rect 7380 3136 7432 3188
rect 7564 3136 7616 3188
rect 7840 3136 7892 3188
rect 9404 3136 9456 3188
rect 12348 3136 12400 3188
rect 4068 3068 4120 3120
rect 3700 3000 3752 3052
rect 4160 3000 4212 3052
rect 7196 3068 7248 3120
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 6368 3000 6420 3052
rect 7288 3000 7340 3052
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 572 2864 624 2916
rect 1492 2864 1544 2916
rect 3424 2864 3476 2916
rect 296 2796 348 2848
rect 1860 2796 1912 2848
rect 3516 2796 3568 2848
rect 3884 2932 3936 2984
rect 5080 2975 5132 2984
rect 5080 2941 5114 2975
rect 5114 2941 5132 2975
rect 5080 2932 5132 2941
rect 7196 2932 7248 2984
rect 11980 3068 12032 3120
rect 9496 3000 9548 3052
rect 11612 3000 11664 3052
rect 11796 3000 11848 3052
rect 4252 2907 4304 2916
rect 4252 2873 4261 2907
rect 4261 2873 4295 2907
rect 4295 2873 4304 2907
rect 4252 2864 4304 2873
rect 4712 2864 4764 2916
rect 4160 2796 4212 2848
rect 5448 2796 5500 2848
rect 7380 2796 7432 2848
rect 7656 2932 7708 2984
rect 8392 2932 8444 2984
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 9864 2932 9916 2984
rect 10692 2932 10744 2984
rect 11060 2932 11112 2984
rect 8668 2864 8720 2916
rect 8944 2796 8996 2848
rect 9404 2796 9456 2848
rect 10968 2864 11020 2916
rect 11060 2796 11112 2848
rect 12164 2864 12216 2916
rect 12992 2796 13044 2848
rect 4723 2694 4775 2746
rect 4787 2694 4839 2746
rect 4851 2694 4903 2746
rect 4915 2694 4967 2746
rect 8464 2694 8516 2746
rect 8528 2694 8580 2746
rect 8592 2694 8644 2746
rect 8656 2694 8708 2746
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4068 2592 4120 2644
rect 4160 2567 4212 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 2136 2499 2188 2508
rect 2136 2465 2145 2499
rect 2145 2465 2179 2499
rect 2179 2465 2188 2499
rect 2136 2456 2188 2465
rect 2780 2456 2832 2508
rect 4160 2533 4194 2567
rect 4194 2533 4212 2567
rect 4160 2524 4212 2533
rect 5172 2592 5224 2644
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 8760 2592 8812 2644
rect 3884 2499 3936 2508
rect 3884 2465 3893 2499
rect 3893 2465 3927 2499
rect 3927 2465 3936 2499
rect 3884 2456 3936 2465
rect 4528 2456 4580 2508
rect 3608 2320 3660 2372
rect 5448 2456 5500 2508
rect 6460 2524 6512 2576
rect 6920 2524 6972 2576
rect 7840 2524 7892 2576
rect 8392 2567 8444 2576
rect 8392 2533 8401 2567
rect 8401 2533 8435 2567
rect 8435 2533 8444 2567
rect 8392 2524 8444 2533
rect 9220 2524 9272 2576
rect 9588 2592 9640 2644
rect 5080 2252 5132 2304
rect 5908 2320 5960 2372
rect 7656 2456 7708 2508
rect 8944 2456 8996 2508
rect 10968 2524 11020 2576
rect 11152 2524 11204 2576
rect 11520 2524 11572 2576
rect 10048 2456 10100 2508
rect 7288 2252 7340 2304
rect 9312 2388 9364 2440
rect 10232 2456 10284 2508
rect 12440 2456 12492 2508
rect 10048 2320 10100 2372
rect 10784 2388 10836 2440
rect 10968 2320 11020 2372
rect 9128 2252 9180 2304
rect 9588 2252 9640 2304
rect 10692 2252 10744 2304
rect 10876 2252 10928 2304
rect 2852 2150 2904 2202
rect 2916 2150 2968 2202
rect 2980 2150 3032 2202
rect 3044 2150 3096 2202
rect 6594 2150 6646 2202
rect 6658 2150 6710 2202
rect 6722 2150 6774 2202
rect 6786 2150 6838 2202
rect 10335 2150 10387 2202
rect 10399 2150 10451 2202
rect 10463 2150 10515 2202
rect 10527 2150 10579 2202
rect 5448 2048 5500 2100
rect 4712 1980 4764 2032
rect 5724 1980 5776 2032
rect 4160 1912 4212 1964
rect 5908 1844 5960 1896
rect 6092 1776 6144 1828
rect 3884 1504 3936 1556
rect 5172 1504 5224 1556
rect 3056 1436 3108 1488
rect 3792 1436 3844 1488
rect 2504 1368 2556 1420
rect 2688 1368 2740 1420
rect 5172 1368 5224 1420
rect 5356 1368 5408 1420
rect 6000 1368 6052 1420
rect 6552 1368 6604 1420
rect 9312 1368 9364 1420
rect 9588 1368 9640 1420
rect 5540 1300 5592 1352
rect 6276 1300 6328 1352
rect 10048 1300 10100 1352
rect 10324 1300 10376 1352
rect 8944 1164 8996 1216
rect 10416 1164 10468 1216
rect 10692 1028 10744 1080
rect 10876 1028 10928 1080
rect 4160 960 4212 1012
rect 5356 960 5408 1012
<< metal2 >>
rect 754 14818 810 15618
rect 2226 14818 2282 15618
rect 3698 14818 3754 15618
rect 5170 14818 5226 15618
rect 6642 14818 6698 15618
rect 8206 14818 8262 15618
rect 9678 14818 9734 15618
rect 11150 14818 11206 15618
rect 12622 14818 12678 15618
rect 572 13456 624 13462
rect 572 13398 624 13404
rect 584 12434 612 13398
rect 664 13388 716 13394
rect 664 13330 716 13336
rect 308 12406 612 12434
rect 112 11892 164 11898
rect 112 11834 164 11840
rect 124 4146 152 11834
rect 204 4684 256 4690
rect 204 4626 256 4632
rect 112 4140 164 4146
rect 112 4082 164 4088
rect 112 4004 164 4010
rect 112 3946 164 3952
rect 20 3936 72 3942
rect 20 3878 72 3884
rect 32 800 60 3878
rect 124 800 152 3946
rect 216 800 244 4626
rect 308 2854 336 12406
rect 572 11076 624 11082
rect 572 11018 624 11024
rect 478 10160 534 10169
rect 478 10095 534 10104
rect 388 7812 440 7818
rect 388 7754 440 7760
rect 400 3874 428 7754
rect 492 4282 520 10095
rect 584 7857 612 11018
rect 570 7848 626 7857
rect 570 7783 626 7792
rect 676 7698 704 13330
rect 768 13002 796 14818
rect 1216 13320 1268 13326
rect 1216 13262 1268 13268
rect 1124 13252 1176 13258
rect 1124 13194 1176 13200
rect 768 12974 888 13002
rect 756 12912 808 12918
rect 756 12854 808 12860
rect 584 7670 704 7698
rect 480 4276 532 4282
rect 480 4218 532 4224
rect 480 4140 532 4146
rect 480 4082 532 4088
rect 388 3868 440 3874
rect 388 3810 440 3816
rect 388 3732 440 3738
rect 388 3674 440 3680
rect 296 2848 348 2854
rect 296 2790 348 2796
rect 400 800 428 3674
rect 492 800 520 4082
rect 584 2922 612 7670
rect 768 7562 796 12854
rect 860 11082 888 12974
rect 940 12980 992 12986
rect 940 12922 992 12928
rect 848 11076 900 11082
rect 848 11018 900 11024
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 676 7534 796 7562
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 676 800 704 7534
rect 754 4040 810 4049
rect 754 3975 810 3984
rect 768 800 796 3975
rect 860 800 888 8366
rect 952 4146 980 12922
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 940 3868 992 3874
rect 940 3810 992 3816
rect 952 2825 980 3810
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1044 800 1072 9522
rect 1136 7562 1164 13194
rect 1228 7698 1256 13262
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 7818 1348 12786
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11558 1440 12174
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10130 1532 10950
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1412 9722 1440 10066
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1398 8936 1454 8945
rect 1398 8871 1454 8880
rect 1412 8634 1440 8871
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1228 7670 1348 7698
rect 1136 7534 1256 7562
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 1136 800 1164 4014
rect 1228 2774 1256 7534
rect 1320 4842 1348 7670
rect 1504 7478 1532 9862
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5914 1440 6190
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1398 5672 1454 5681
rect 1398 5607 1400 5616
rect 1452 5607 1454 5616
rect 1400 5578 1452 5584
rect 1320 4814 1440 4842
rect 1228 2746 1348 2774
rect 1320 800 1348 2746
rect 1412 800 1440 4814
rect 1504 3058 1532 7278
rect 1596 5658 1624 12582
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11354 1716 12242
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10810 1808 11154
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1780 10062 1808 10231
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9110 1808 9998
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8634 1716 8978
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 7886 1808 8366
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1872 7562 1900 12650
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12434 2084 12582
rect 1964 12406 2084 12434
rect 1964 8090 1992 12406
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11762 2176 12038
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 11286 2084 11494
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2148 11218 2176 11698
rect 2240 11354 2268 14818
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11830 2452 12242
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2424 10674 2452 11766
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2240 9586 2268 10610
rect 2516 10606 2544 11018
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10130 2452 10406
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2318 9752 2374 9761
rect 2318 9687 2374 9696
rect 2228 9580 2280 9586
rect 2056 9540 2228 9568
rect 2056 8430 2084 9540
rect 2228 9522 2280 9528
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8537 2268 8978
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1780 7534 1900 7562
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6458 1716 6802
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5778 1716 6054
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1596 5630 1716 5658
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1596 2990 1624 4422
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1492 2916 1544 2922
rect 1492 2858 1544 2864
rect 1504 800 1532 2858
rect 1596 2514 1624 2926
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1688 800 1716 5630
rect 1780 800 1808 7534
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 3126 1900 7278
rect 1964 4146 1992 7414
rect 2056 5914 2084 8230
rect 2148 8090 2176 8298
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 6866 2176 7822
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2148 6322 2176 6802
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2136 6112 2188 6118
rect 2134 6080 2136 6089
rect 2188 6080 2190 6089
rect 2134 6015 2190 6024
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5166 2084 5510
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2148 4214 2176 5714
rect 2136 4208 2188 4214
rect 2056 4168 2136 4196
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1964 2990 1992 3878
rect 2056 3126 2084 4168
rect 2136 4150 2188 4156
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 2148 2990 2176 4014
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 1034 1900 2790
rect 1964 2514 1992 2926
rect 2042 2816 2098 2825
rect 2042 2751 2098 2760
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1872 1006 1992 1034
rect 1964 800 1992 1006
rect 2056 800 2084 2751
rect 2148 2514 2176 2926
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2240 1442 2268 8366
rect 2332 7546 2360 9687
rect 2516 9110 2544 10542
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 7426 2452 8910
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2332 7398 2452 7426
rect 2332 4706 2360 7398
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 6361 2452 7278
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5778 2452 6190
rect 2516 6066 2544 8774
rect 2608 7002 2636 12582
rect 2700 9518 2728 13126
rect 2826 13084 3122 13104
rect 2882 13082 2906 13084
rect 2962 13082 2986 13084
rect 3042 13082 3066 13084
rect 2904 13030 2906 13082
rect 2968 13030 2980 13082
rect 3042 13030 3044 13082
rect 2882 13028 2906 13030
rect 2962 13028 2986 13030
rect 3042 13028 3066 13030
rect 2826 13008 3122 13028
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2826 11996 3122 12016
rect 2882 11994 2906 11996
rect 2962 11994 2986 11996
rect 3042 11994 3066 11996
rect 2904 11942 2906 11994
rect 2968 11942 2980 11994
rect 3042 11942 3044 11994
rect 2882 11940 2906 11942
rect 2962 11940 2986 11942
rect 3042 11940 3066 11942
rect 2826 11920 3122 11940
rect 3054 11656 3110 11665
rect 2780 11620 2832 11626
rect 3054 11591 3110 11600
rect 2780 11562 2832 11568
rect 2792 11354 2820 11562
rect 3068 11354 3096 11591
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2826 10908 3122 10928
rect 2882 10906 2906 10908
rect 2962 10906 2986 10908
rect 3042 10906 3066 10908
rect 2904 10854 2906 10906
rect 2968 10854 2980 10906
rect 3042 10854 3044 10906
rect 2882 10852 2906 10854
rect 2962 10852 2986 10854
rect 3042 10852 3066 10854
rect 2826 10832 3122 10852
rect 3252 10742 3280 12582
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 11218 3372 11494
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 2780 10736 2832 10742
rect 2778 10704 2780 10713
rect 3240 10736 3292 10742
rect 2832 10704 2834 10713
rect 3240 10678 3292 10684
rect 3344 10674 3372 11154
rect 3436 10810 3464 12650
rect 3712 12374 3740 14818
rect 5184 12986 5212 14818
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12374 4292 12582
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11626 3648 12038
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 2778 10639 2834 10648
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10441 2820 10542
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 2872 10464 2924 10470
rect 2778 10432 2834 10441
rect 2872 10406 2924 10412
rect 2778 10367 2834 10376
rect 2884 10266 2912 10406
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2976 9994 3004 10474
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3160 10198 3188 10406
rect 3252 10305 3280 10406
rect 3238 10296 3294 10305
rect 3238 10231 3294 10240
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 3252 9874 3280 10231
rect 3344 9897 3372 10474
rect 3422 10160 3478 10169
rect 3422 10095 3424 10104
rect 3476 10095 3478 10104
rect 3424 10066 3476 10072
rect 3528 10010 3556 10746
rect 3620 10538 3648 11562
rect 3712 10674 3740 12174
rect 4448 11694 4476 12242
rect 4540 11762 4568 12786
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4632 11898 4660 12718
rect 4697 12540 4993 12560
rect 4753 12538 4777 12540
rect 4833 12538 4857 12540
rect 4913 12538 4937 12540
rect 4775 12486 4777 12538
rect 4839 12486 4851 12538
rect 4913 12486 4915 12538
rect 4753 12484 4777 12486
rect 4833 12484 4857 12486
rect 4913 12484 4937 12486
rect 4697 12464 4993 12484
rect 5092 12442 5120 12718
rect 5080 12436 5132 12442
rect 5000 12406 5080 12434
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11688 4488 11694
rect 4724 11642 4752 12310
rect 5000 12306 5028 12406
rect 5080 12378 5132 12384
rect 5184 12374 5212 12718
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5078 11792 5134 11801
rect 5078 11727 5080 11736
rect 5132 11727 5134 11736
rect 5080 11698 5132 11704
rect 4436 11630 4488 11636
rect 4632 11614 4752 11642
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3606 10160 3662 10169
rect 3606 10095 3662 10104
rect 3436 9982 3556 10010
rect 3160 9846 3280 9874
rect 3330 9888 3386 9897
rect 2826 9820 3122 9840
rect 2882 9818 2906 9820
rect 2962 9818 2986 9820
rect 3042 9818 3066 9820
rect 2904 9766 2906 9818
rect 2968 9766 2980 9818
rect 3042 9766 3044 9818
rect 2882 9764 2906 9766
rect 2962 9764 2986 9766
rect 3042 9764 3066 9766
rect 2826 9744 3122 9764
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 9518 2820 9590
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 9178 2820 9318
rect 2780 9172 2832 9178
rect 2700 9132 2780 9160
rect 2700 8362 2728 9132
rect 2780 9114 2832 9120
rect 3160 8956 3188 9846
rect 3330 9823 3386 9832
rect 3436 9738 3464 9982
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3252 9710 3464 9738
rect 3252 9217 3280 9710
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3436 9518 3464 9590
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3238 9208 3294 9217
rect 3238 9143 3294 9152
rect 3240 9104 3292 9110
rect 3292 9064 3464 9092
rect 3240 9046 3292 9052
rect 3240 8968 3292 8974
rect 3160 8928 3240 8956
rect 2826 8732 3122 8752
rect 2882 8730 2906 8732
rect 2962 8730 2986 8732
rect 3042 8730 3066 8732
rect 2904 8678 2906 8730
rect 2968 8678 2980 8730
rect 3042 8678 3044 8730
rect 2882 8676 2906 8678
rect 2962 8676 2986 8678
rect 3042 8676 3066 8678
rect 2826 8656 3122 8676
rect 2872 8560 2924 8566
rect 3160 8514 3188 8928
rect 3240 8910 3292 8916
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2872 8502 2924 8508
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2884 7954 2912 8502
rect 2976 8486 3188 8514
rect 2976 8362 3004 8486
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 8090 3096 8298
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3252 7954 3280 8570
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 2700 7546 2728 7890
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 2826 7644 3122 7664
rect 2882 7642 2906 7644
rect 2962 7642 2986 7644
rect 3042 7642 3066 7644
rect 2904 7590 2906 7642
rect 2968 7590 2980 7642
rect 3042 7590 3044 7642
rect 2882 7588 2906 7590
rect 2962 7588 2986 7590
rect 3042 7588 3066 7590
rect 2826 7568 3122 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 3160 7478 3188 7754
rect 3252 7546 3280 7754
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2792 6769 2820 7210
rect 2778 6760 2834 6769
rect 2884 6730 2912 7278
rect 3068 6769 3096 7278
rect 3054 6760 3110 6769
rect 2778 6695 2834 6704
rect 2872 6724 2924 6730
rect 3054 6695 3110 6704
rect 2872 6666 2924 6672
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6254 2636 6598
rect 2826 6556 3122 6576
rect 2882 6554 2906 6556
rect 2962 6554 2986 6556
rect 3042 6554 3066 6556
rect 2904 6502 2906 6554
rect 2968 6502 2980 6554
rect 3042 6502 3044 6554
rect 2882 6500 2906 6502
rect 2962 6500 2986 6502
rect 3042 6500 3066 6502
rect 2826 6480 3122 6500
rect 3160 6474 3188 7414
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3252 6633 3280 7278
rect 3238 6624 3294 6633
rect 3238 6559 3294 6568
rect 3160 6446 3280 6474
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2516 6038 2636 6066
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5370 2544 5646
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2424 4826 2452 5034
rect 2516 4826 2544 5306
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2332 4678 2452 4706
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 3641 2360 4558
rect 2318 3632 2374 3641
rect 2318 3567 2374 3576
rect 2318 3496 2374 3505
rect 2318 3431 2374 3440
rect 2148 1414 2268 1442
rect 2148 800 2176 1414
rect 2332 800 2360 3431
rect 2424 800 2452 4678
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2516 4282 2544 4626
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 1426 2544 4082
rect 2608 4078 2636 6038
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5302 2728 5714
rect 3068 5642 3096 6190
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2826 5468 3122 5488
rect 2882 5466 2906 5468
rect 2962 5466 2986 5468
rect 3042 5466 3066 5468
rect 2904 5414 2906 5466
rect 2968 5414 2980 5466
rect 3042 5414 3044 5466
rect 2882 5412 2906 5414
rect 2962 5412 2986 5414
rect 3042 5412 3066 5414
rect 2826 5392 3122 5412
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2686 4856 2742 4865
rect 2686 4791 2742 4800
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2700 3924 2728 4791
rect 3160 4690 3188 6258
rect 3252 6186 3280 6446
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3252 5846 3280 6122
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5166 3280 5510
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2826 4380 3122 4400
rect 2882 4378 2906 4380
rect 2962 4378 2986 4380
rect 3042 4378 3066 4380
rect 2904 4326 2906 4378
rect 2968 4326 2980 4378
rect 3042 4326 3044 4378
rect 2882 4324 2906 4326
rect 2962 4324 2986 4326
rect 3042 4324 3066 4326
rect 2826 4304 3122 4324
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2608 3896 2728 3924
rect 2504 1420 2556 1426
rect 2504 1362 2556 1368
rect 2608 800 2636 3896
rect 2976 3602 3004 4150
rect 3160 4078 3188 4626
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3068 3738 3096 4014
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3160 3534 3188 3878
rect 3252 3738 3280 4762
rect 3344 4162 3372 8774
rect 3436 8430 3464 9064
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3436 7954 3464 8366
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3436 7546 3464 7890
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 6458 3464 7278
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3436 5914 3464 6190
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3422 4856 3478 4865
rect 3422 4791 3478 4800
rect 3436 4690 3464 4791
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 4282 3464 4422
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3344 4134 3464 4162
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3344 3738 3372 4014
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3618 3464 4134
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3344 3590 3464 3618
rect 3148 3528 3200 3534
rect 3054 3496 3110 3505
rect 3148 3470 3200 3476
rect 3054 3431 3110 3440
rect 2688 3392 2740 3398
rect 3068 3380 3096 3431
rect 3068 3352 3188 3380
rect 2688 3334 2740 3340
rect 2700 2088 2728 3334
rect 2826 3292 3122 3312
rect 2882 3290 2906 3292
rect 2962 3290 2986 3292
rect 3042 3290 3066 3292
rect 2904 3238 2906 3290
rect 2968 3238 2980 3290
rect 3042 3238 3044 3290
rect 2882 3236 2906 3238
rect 2962 3236 2986 3238
rect 3042 3236 3066 3238
rect 2826 3216 3122 3236
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3054 3088 3110 3097
rect 2792 2514 2820 3062
rect 3160 3074 3188 3352
rect 3252 3194 3280 3538
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3160 3046 3280 3074
rect 3054 3023 3056 3032
rect 3108 3023 3110 3032
rect 3056 2994 3108 3000
rect 3148 2984 3200 2990
rect 3146 2952 3148 2961
rect 3200 2952 3202 2961
rect 3146 2887 3202 2896
rect 3054 2680 3110 2689
rect 3054 2615 3110 2624
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 3068 2394 3096 2615
rect 3068 2366 3188 2394
rect 2826 2204 3122 2224
rect 2882 2202 2906 2204
rect 2962 2202 2986 2204
rect 3042 2202 3066 2204
rect 2904 2150 2906 2202
rect 2968 2150 2980 2202
rect 3042 2150 3044 2202
rect 2882 2148 2906 2150
rect 2962 2148 2986 2150
rect 3042 2148 3066 2150
rect 2826 2128 3122 2148
rect 2700 2060 2820 2088
rect 2688 1420 2740 1426
rect 2688 1362 2740 1368
rect 2700 800 2728 1362
rect 2792 800 2820 2060
rect 3160 1578 3188 2366
rect 2976 1550 3188 1578
rect 2976 800 3004 1550
rect 3056 1488 3108 1494
rect 3056 1430 3108 1436
rect 3068 800 3096 1430
rect 3252 800 3280 3046
rect 3344 2650 3372 3590
rect 3528 3482 3556 9862
rect 3620 6905 3648 10095
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3620 5030 3648 6734
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4570 3648 4966
rect 3712 4808 3740 10367
rect 3804 5846 3832 10678
rect 3896 10282 3924 11154
rect 3988 10470 4016 11494
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3896 10254 4016 10282
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 8537 3924 10066
rect 3988 9926 4016 10254
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 4080 9722 4108 10950
rect 4172 10266 4200 11086
rect 4264 10538 4292 11222
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4243 10532 4295 10538
rect 4243 10474 4295 10480
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9217 4016 9318
rect 3974 9208 4030 9217
rect 4080 9178 4108 9658
rect 3974 9143 4030 9152
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3988 8362 4016 9046
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 8129 3924 8230
rect 3882 8120 3938 8129
rect 3882 8055 3938 8064
rect 3988 8022 4016 8298
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3896 7002 3924 7890
rect 4080 7886 4108 8774
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4172 7426 4200 10066
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4080 7398 4200 7426
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6254 3924 6598
rect 3988 6458 4016 7346
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 6118 3924 6190
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3988 5273 4016 6122
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 4080 5114 4108 7398
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4172 6866 4200 7278
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3988 5086 4108 5114
rect 3988 4826 4016 5086
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4172 4826 4200 5646
rect 3976 4820 4028 4826
rect 3712 4780 3924 4808
rect 3792 4684 3844 4690
rect 3712 4622 3740 4653
rect 3792 4626 3844 4632
rect 3700 4616 3752 4622
rect 3620 4564 3700 4570
rect 3620 4558 3752 4564
rect 3620 4542 3740 4558
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4146 3648 4422
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3712 4078 3740 4542
rect 3804 4078 3832 4626
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3712 3913 3740 4014
rect 3698 3904 3754 3913
rect 3698 3839 3754 3848
rect 3896 3754 3924 4780
rect 3976 4762 4028 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 4068 4684 4120 4690
rect 4120 4644 4200 4672
rect 4068 4626 4120 4632
rect 3988 4593 4016 4626
rect 3974 4584 4030 4593
rect 3974 4519 4030 4528
rect 3988 3924 4016 4519
rect 4068 3936 4120 3942
rect 3988 3896 4068 3924
rect 4068 3878 4120 3884
rect 3712 3726 3924 3754
rect 4066 3768 4122 3777
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3436 3454 3556 3482
rect 3436 2922 3464 3454
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2990 3556 3334
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3516 2848 3568 2854
rect 3436 2796 3516 2802
rect 3436 2790 3568 2796
rect 3436 2774 3556 2790
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3330 2544 3386 2553
rect 3330 2479 3386 2488
rect 3344 800 3372 2479
rect 3436 800 3464 2774
rect 3620 2378 3648 3538
rect 3712 3058 3740 3726
rect 4172 3738 4200 4644
rect 4066 3703 4122 3712
rect 4160 3732 4212 3738
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3698 2952 3754 2961
rect 3698 2887 3754 2896
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3712 1442 3740 2887
rect 3804 1494 3832 3606
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3896 3194 3924 3538
rect 3976 3392 4028 3398
rect 3974 3360 3976 3369
rect 4028 3360 4030 3369
rect 3974 3295 4030 3304
rect 4080 3210 4108 3703
rect 4160 3674 4212 3680
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3988 3182 4108 3210
rect 4172 3194 4200 3402
rect 4160 3188 4212 3194
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3896 2514 3924 2926
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 3620 1414 3740 1442
rect 3792 1488 3844 1494
rect 3792 1430 3844 1436
rect 3620 800 3648 1414
rect 3698 1320 3754 1329
rect 3698 1255 3754 1264
rect 3712 800 3740 1255
rect 3896 800 3924 1498
rect 3988 800 4016 3182
rect 4160 3130 4212 3136
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4158 3088 4214 3097
rect 4080 2650 4108 3062
rect 4158 3023 4160 3032
rect 4212 3023 4214 3032
rect 4160 2994 4212 3000
rect 4264 2922 4292 9930
rect 4356 5794 4384 11086
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 10305 4476 11018
rect 4434 10296 4490 10305
rect 4434 10231 4490 10240
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4448 8378 4476 10066
rect 4540 8514 4568 11154
rect 4632 10849 4660 11614
rect 4697 11452 4993 11472
rect 4753 11450 4777 11452
rect 4833 11450 4857 11452
rect 4913 11450 4937 11452
rect 4775 11398 4777 11450
rect 4839 11398 4851 11450
rect 4913 11398 4915 11450
rect 4753 11396 4777 11398
rect 4833 11396 4857 11398
rect 4913 11396 4937 11398
rect 4697 11376 4993 11396
rect 5276 11370 5304 12786
rect 5552 12782 5580 13194
rect 6288 12782 6316 13262
rect 6656 13172 6684 14818
rect 8220 13682 8248 14818
rect 8220 13654 8432 13682
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6656 13144 6960 13172
rect 6568 13084 6864 13104
rect 6624 13082 6648 13084
rect 6704 13082 6728 13084
rect 6784 13082 6808 13084
rect 6646 13030 6648 13082
rect 6710 13030 6722 13082
rect 6784 13030 6786 13082
rect 6624 13028 6648 13030
rect 6704 13028 6728 13030
rect 6784 13028 6808 13030
rect 6568 13008 6864 13028
rect 6932 12986 6960 13144
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 11830 5396 12582
rect 5644 12442 5672 12718
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5460 11370 5488 11766
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5184 11342 5304 11370
rect 5368 11342 5488 11370
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 11098 4844 11154
rect 4724 11070 4844 11098
rect 4618 10840 4674 10849
rect 4618 10775 4674 10784
rect 4724 10577 4752 11070
rect 5184 11014 5212 11342
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4816 10713 4844 10950
rect 4802 10704 4858 10713
rect 4802 10639 4858 10648
rect 4908 10577 4936 10950
rect 4710 10568 4766 10577
rect 4710 10503 4766 10512
rect 4894 10568 4950 10577
rect 4894 10503 4950 10512
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10130 4660 10406
rect 4697 10364 4993 10384
rect 4753 10362 4777 10364
rect 4833 10362 4857 10364
rect 4913 10362 4937 10364
rect 4775 10310 4777 10362
rect 4839 10310 4851 10362
rect 4913 10310 4915 10362
rect 4753 10308 4777 10310
rect 4833 10308 4857 10310
rect 4913 10308 4937 10310
rect 4697 10288 4993 10308
rect 5170 10296 5226 10305
rect 5170 10231 5226 10240
rect 4896 10192 4948 10198
rect 4948 10140 5120 10146
rect 4896 10134 5120 10140
rect 4908 10130 5120 10134
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4712 10124 4764 10130
rect 4908 10124 5132 10130
rect 4908 10118 5080 10124
rect 4764 10084 4844 10112
rect 4712 10066 4764 10072
rect 4632 9518 4660 10066
rect 4712 9920 4764 9926
rect 4710 9888 4712 9897
rect 4764 9888 4766 9897
rect 4710 9823 4766 9832
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4724 9364 4752 9658
rect 4816 9450 4844 10084
rect 5080 10066 5132 10072
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9489 4936 9998
rect 5080 9920 5132 9926
rect 4986 9888 5042 9897
rect 5080 9862 5132 9868
rect 4986 9823 5042 9832
rect 5000 9722 5028 9823
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 5092 9625 5120 9862
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 5080 9512 5132 9518
rect 4894 9480 4950 9489
rect 4804 9444 4856 9450
rect 5080 9454 5132 9460
rect 4894 9415 4950 9424
rect 4804 9386 4856 9392
rect 4632 9336 4752 9364
rect 4632 9110 4660 9336
rect 4697 9276 4993 9296
rect 4753 9274 4777 9276
rect 4833 9274 4857 9276
rect 4913 9274 4937 9276
rect 4775 9222 4777 9274
rect 4839 9222 4851 9274
rect 4913 9222 4915 9274
rect 4753 9220 4777 9222
rect 4833 9220 4857 9222
rect 4913 9220 4937 9222
rect 4697 9200 4993 9220
rect 5092 9217 5120 9454
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 4816 9110 4844 9141
rect 4620 9104 4672 9110
rect 4804 9104 4856 9110
rect 4620 9046 4672 9052
rect 4802 9072 4804 9081
rect 4856 9072 4858 9081
rect 4712 9036 4764 9042
rect 4802 9007 4858 9016
rect 4986 9072 5042 9081
rect 4986 9007 5042 9016
rect 4712 8978 4764 8984
rect 4724 8945 4752 8978
rect 4710 8936 4766 8945
rect 4710 8871 4766 8880
rect 4816 8838 4844 9007
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4540 8486 4660 8514
rect 5000 8498 5028 9007
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 8498 5120 8910
rect 4448 8350 4568 8378
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7954 4476 8230
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4448 5953 4476 6190
rect 4434 5944 4490 5953
rect 4434 5879 4490 5888
rect 4356 5766 4476 5794
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 5370 4384 5646
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4356 4690 4384 5306
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4342 4584 4398 4593
rect 4342 4519 4398 4528
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4172 2582 4200 2790
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4066 2272 4122 2281
rect 4066 2207 4122 2216
rect 4080 800 4108 2207
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4172 1018 4200 1906
rect 4250 1184 4306 1193
rect 4250 1119 4306 1128
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 4264 800 4292 1119
rect 4356 800 4384 4519
rect 4448 3777 4476 5766
rect 4434 3768 4490 3777
rect 4434 3703 4490 3712
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4448 2836 4476 3470
rect 4540 2961 4568 8350
rect 4632 7426 4660 8486
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4697 8188 4993 8208
rect 4753 8186 4777 8188
rect 4833 8186 4857 8188
rect 4913 8186 4937 8188
rect 4775 8134 4777 8186
rect 4839 8134 4851 8186
rect 4913 8134 4915 8186
rect 4753 8132 4777 8134
rect 4833 8132 4857 8134
rect 4913 8132 4937 8134
rect 4697 8112 4993 8132
rect 5078 7576 5134 7585
rect 5078 7511 5080 7520
rect 5132 7511 5134 7520
rect 5080 7482 5132 7488
rect 4632 7398 5120 7426
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 7188 4752 7278
rect 4632 7160 4752 7188
rect 4632 6984 4660 7160
rect 4697 7100 4993 7120
rect 4753 7098 4777 7100
rect 4833 7098 4857 7100
rect 4913 7098 4937 7100
rect 4775 7046 4777 7098
rect 4839 7046 4851 7098
rect 4913 7046 4915 7098
rect 4753 7044 4777 7046
rect 4833 7044 4857 7046
rect 4913 7044 4937 7046
rect 4697 7024 4993 7044
rect 4632 6956 4752 6984
rect 4618 6760 4674 6769
rect 4618 6695 4674 6704
rect 4632 5386 4660 6695
rect 4724 6225 4752 6956
rect 4710 6216 4766 6225
rect 4710 6151 4766 6160
rect 4697 6012 4993 6032
rect 4753 6010 4777 6012
rect 4833 6010 4857 6012
rect 4913 6010 4937 6012
rect 4775 5958 4777 6010
rect 4839 5958 4851 6010
rect 4913 5958 4915 6010
rect 4753 5956 4777 5958
rect 4833 5956 4857 5958
rect 4913 5956 4937 5958
rect 4697 5936 4993 5956
rect 5092 5930 5120 7398
rect 5184 6322 5212 10231
rect 5276 7206 5304 11154
rect 5368 9518 5396 11342
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10588 5488 11154
rect 5552 10810 5580 11698
rect 5644 11626 5672 12378
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5920 11898 5948 12242
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5630 11384 5686 11393
rect 5630 11319 5632 11328
rect 5684 11319 5686 11328
rect 5632 11290 5684 11296
rect 5630 11248 5686 11257
rect 5630 11183 5632 11192
rect 5684 11183 5686 11192
rect 5632 11154 5684 11160
rect 5736 11121 5764 11630
rect 5722 11112 5778 11121
rect 5722 11047 5778 11056
rect 5630 10976 5686 10985
rect 5630 10911 5686 10920
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10600 5592 10606
rect 5460 10560 5540 10588
rect 5460 10441 5488 10560
rect 5540 10542 5592 10548
rect 5540 10464 5592 10470
rect 5446 10432 5502 10441
rect 5540 10406 5592 10412
rect 5446 10367 5502 10376
rect 5460 9518 5488 10367
rect 5552 10130 5580 10406
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9625 5580 9862
rect 5538 9616 5594 9625
rect 5538 9551 5594 9560
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5354 9344 5410 9353
rect 5354 9279 5410 9288
rect 5368 8566 5396 9279
rect 5552 9217 5580 9386
rect 5538 9208 5594 9217
rect 5538 9143 5594 9152
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5540 8424 5592 8430
rect 5644 8401 5672 10911
rect 5828 10282 5856 11698
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5736 10254 5856 10282
rect 5540 8366 5592 8372
rect 5630 8392 5686 8401
rect 5368 8090 5396 8366
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5460 7528 5488 8230
rect 5552 7546 5580 8366
rect 5630 8327 5686 8336
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8022 5672 8230
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5368 7500 5488 7528
rect 5540 7540 5592 7546
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5262 6896 5318 6905
rect 5262 6831 5264 6840
rect 5316 6831 5318 6840
rect 5264 6802 5316 6808
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5092 5902 5212 5930
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 4632 5358 4752 5386
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4526 2952 4582 2961
rect 4526 2887 4582 2896
rect 4448 2808 4568 2836
rect 4434 2544 4490 2553
rect 4540 2514 4568 2808
rect 4434 2479 4490 2488
rect 4528 2508 4580 2514
rect 4448 1306 4476 2479
rect 4528 2450 4580 2456
rect 4632 2122 4660 5238
rect 4724 5166 4752 5358
rect 4908 5302 4936 5714
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 5092 5098 5120 5714
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 4697 4924 4993 4944
rect 4753 4922 4777 4924
rect 4833 4922 4857 4924
rect 4913 4922 4937 4924
rect 4775 4870 4777 4922
rect 4839 4870 4851 4922
rect 4913 4870 4915 4922
rect 4753 4868 4777 4870
rect 4833 4868 4857 4870
rect 4913 4868 4937 4870
rect 4697 4848 4993 4868
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4282 4936 4422
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4908 4049 4936 4218
rect 4894 4040 4950 4049
rect 5000 4010 5028 4626
rect 4894 3975 4950 3984
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4697 3836 4993 3856
rect 4753 3834 4777 3836
rect 4833 3834 4857 3836
rect 4913 3834 4937 3836
rect 4775 3782 4777 3834
rect 4839 3782 4851 3834
rect 4913 3782 4915 3834
rect 4753 3780 4777 3782
rect 4833 3780 4857 3782
rect 4913 3780 4937 3782
rect 4697 3760 4993 3780
rect 5092 3720 5120 5034
rect 5184 3754 5212 5902
rect 5276 3856 5304 6054
rect 5368 5302 5396 7500
rect 5736 7528 5764 10254
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5828 9722 5856 10134
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5540 7482 5592 7488
rect 5644 7500 5764 7528
rect 5644 7426 5672 7500
rect 5460 7398 5672 7426
rect 5460 6712 5488 7398
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5632 7336 5684 7342
rect 5684 7296 5856 7324
rect 5632 7278 5684 7284
rect 5552 6934 5580 7278
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5644 6866 5672 7142
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5460 6684 5764 6712
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5460 5846 5488 6559
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5368 4826 5396 5238
rect 5460 5001 5488 5510
rect 5446 4992 5502 5001
rect 5446 4927 5502 4936
rect 5446 4856 5502 4865
rect 5356 4820 5408 4826
rect 5446 4791 5502 4800
rect 5356 4762 5408 4768
rect 5460 4486 5488 4791
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5552 4128 5580 6394
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5644 4282 5672 4694
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5552 4100 5672 4128
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5276 3828 5396 3856
rect 5184 3726 5304 3754
rect 5000 3692 5120 3720
rect 4710 3632 4766 3641
rect 4710 3567 4766 3576
rect 4894 3632 4950 3641
rect 4894 3567 4896 3576
rect 4724 2922 4752 3567
rect 4948 3567 4950 3576
rect 4896 3538 4948 3544
rect 4908 3398 4936 3538
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4802 3088 4858 3097
rect 4802 3023 4804 3032
rect 4856 3023 4858 3032
rect 4804 2994 4856 3000
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 5000 2836 5028 3692
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 2990 5120 3334
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5000 2808 5120 2836
rect 4697 2748 4993 2768
rect 4753 2746 4777 2748
rect 4833 2746 4857 2748
rect 4913 2746 4937 2748
rect 4775 2694 4777 2746
rect 4839 2694 4851 2746
rect 4913 2694 4915 2746
rect 4753 2692 4777 2694
rect 4833 2692 4857 2694
rect 4913 2692 4937 2694
rect 4697 2672 4993 2692
rect 5092 2310 5120 2808
rect 5184 2650 5212 3538
rect 5276 3233 5304 3726
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 5262 2952 5318 2961
rect 5262 2887 5318 2896
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5170 2408 5226 2417
rect 5170 2343 5226 2352
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4632 2094 5028 2122
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4448 1278 4568 1306
rect 4540 800 4568 1278
rect 4618 1048 4674 1057
rect 4618 983 4674 992
rect 4632 800 4660 983
rect 4724 800 4752 1974
rect 4894 1728 4950 1737
rect 4894 1663 4950 1672
rect 4908 800 4936 1663
rect 5000 800 5028 2094
rect 5184 1562 5212 2343
rect 5172 1556 5224 1562
rect 5172 1498 5224 1504
rect 5172 1420 5224 1426
rect 5172 1362 5224 1368
rect 5184 800 5212 1362
rect 5276 800 5304 2887
rect 5368 1426 5396 3828
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 2854 5488 3538
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 2106 5488 2450
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 5446 1592 5502 1601
rect 5446 1527 5502 1536
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 5460 1170 5488 1527
rect 5552 1358 5580 3946
rect 5644 2961 5672 4100
rect 5630 2952 5686 2961
rect 5630 2887 5686 2896
rect 5630 2544 5686 2553
rect 5630 2479 5686 2488
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5460 1142 5580 1170
rect 5356 1012 5408 1018
rect 5356 954 5408 960
rect 5368 800 5396 954
rect 5552 800 5580 1142
rect 5644 800 5672 2479
rect 5736 2038 5764 6684
rect 5828 6458 5856 7296
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5814 6352 5870 6361
rect 5814 6287 5870 6296
rect 5828 4593 5856 6287
rect 5920 5846 5948 11494
rect 6012 11121 6040 11630
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5998 11112 6054 11121
rect 5998 11047 6054 11056
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6012 10742 6040 10950
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 7954 6040 10406
rect 6104 9178 6132 11494
rect 6196 11354 6224 12650
rect 6656 12646 6684 12786
rect 7300 12782 7328 13330
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12986 7972 13126
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6380 12170 6408 12378
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6568 11996 6864 12016
rect 6624 11994 6648 11996
rect 6704 11994 6728 11996
rect 6784 11994 6808 11996
rect 6646 11942 6648 11994
rect 6710 11942 6722 11994
rect 6784 11942 6786 11994
rect 6624 11940 6648 11942
rect 6704 11940 6728 11942
rect 6784 11940 6808 11942
rect 6568 11920 6864 11940
rect 6932 11898 6960 12242
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6550 11792 6606 11801
rect 6368 11756 6420 11762
rect 6550 11727 6606 11736
rect 6368 11698 6420 11704
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6182 11112 6238 11121
rect 6182 11047 6238 11056
rect 6196 10606 6224 11047
rect 6288 10690 6316 11222
rect 6380 10810 6408 11698
rect 6564 11694 6592 11727
rect 7208 11694 7236 12718
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11694 7788 12310
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 6458 11384 6514 11393
rect 6564 11354 6592 11630
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 6458 11319 6514 11328
rect 6552 11348 6604 11354
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6288 10662 6408 10690
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6380 10470 6408 10662
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6196 9761 6224 10406
rect 6274 10160 6330 10169
rect 6274 10095 6330 10104
rect 6182 9752 6238 9761
rect 6182 9687 6238 9696
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6196 8566 6224 9454
rect 6288 9110 6316 10095
rect 6472 9874 6500 11319
rect 6552 11290 6604 11296
rect 6564 11121 6592 11290
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6550 11112 6606 11121
rect 6932 11098 6960 11154
rect 6932 11070 7052 11098
rect 6550 11047 6606 11056
rect 6568 10908 6864 10928
rect 6624 10906 6648 10908
rect 6704 10906 6728 10908
rect 6784 10906 6808 10908
rect 6646 10854 6648 10906
rect 6710 10854 6722 10906
rect 6784 10854 6786 10906
rect 6624 10852 6648 10854
rect 6704 10852 6728 10854
rect 6784 10852 6808 10854
rect 6568 10832 6864 10852
rect 7024 10810 7052 11070
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6550 10704 6606 10713
rect 6550 10639 6606 10648
rect 6564 10538 6592 10639
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6656 10441 6684 10542
rect 6736 10464 6788 10470
rect 6642 10432 6698 10441
rect 6736 10406 6788 10412
rect 6642 10367 6698 10376
rect 6748 10305 6776 10406
rect 6734 10296 6790 10305
rect 6734 10231 6790 10240
rect 6932 10169 6960 10542
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6380 9846 6500 9874
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6380 9654 6408 9846
rect 6568 9820 6864 9840
rect 6624 9818 6648 9820
rect 6704 9818 6728 9820
rect 6784 9818 6808 9820
rect 6646 9766 6648 9818
rect 6710 9766 6722 9818
rect 6784 9766 6786 9818
rect 6624 9764 6648 9766
rect 6704 9764 6728 9766
rect 6784 9764 6808 9766
rect 6568 9744 6864 9764
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6196 8022 6224 8502
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6288 7954 6316 8774
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6012 7274 6040 7346
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5814 4584 5870 4593
rect 5814 4519 5870 4528
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5828 4282 5856 4383
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5920 4185 5948 4966
rect 5906 4176 5962 4185
rect 5906 4111 5962 4120
rect 5814 3632 5870 3641
rect 5920 3602 5948 4111
rect 5814 3567 5870 3576
rect 5908 3596 5960 3602
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 5828 800 5856 3567
rect 5908 3538 5960 3544
rect 5920 2378 5948 3538
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5920 1034 5948 1838
rect 6012 1426 6040 6870
rect 6104 6390 6132 7686
rect 6196 7410 6224 7686
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6288 7290 6316 7754
rect 6196 7274 6316 7290
rect 6184 7268 6316 7274
rect 6236 7262 6316 7268
rect 6184 7210 6236 7216
rect 6196 6866 6224 7210
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6633 6224 6802
rect 6182 6624 6238 6633
rect 6182 6559 6238 6568
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 4593 6132 5578
rect 6090 4584 6146 4593
rect 6090 4519 6146 4528
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4214 6132 4422
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 6092 4072 6144 4078
rect 6090 4040 6092 4049
rect 6144 4040 6146 4049
rect 6090 3975 6146 3984
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3602 6132 3878
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6104 3194 6132 3538
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 5920 1006 6040 1034
rect 5906 912 5962 921
rect 5906 847 5962 856
rect 5920 800 5948 847
rect 6012 800 6040 1006
rect 6104 898 6132 1770
rect 6196 1442 6224 6190
rect 6288 5846 6316 7142
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6274 5128 6330 5137
rect 6274 5063 6276 5072
rect 6328 5063 6330 5072
rect 6276 5034 6328 5040
rect 6380 4570 6408 9454
rect 6472 8945 6500 9658
rect 6932 9586 6960 9862
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6550 9208 6606 9217
rect 6550 9143 6606 9152
rect 6458 8936 6514 8945
rect 6458 8871 6514 8880
rect 6564 8820 6592 9143
rect 6656 8906 6684 9454
rect 6932 9178 6960 9522
rect 7024 9500 7052 10746
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9722 7144 10066
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7104 9512 7156 9518
rect 7024 9472 7104 9500
rect 7104 9454 7156 9460
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6918 9072 6974 9081
rect 6918 9007 6920 9016
rect 6972 9007 6974 9016
rect 6920 8978 6972 8984
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6472 8792 6592 8820
rect 6472 8616 6500 8792
rect 6568 8732 6864 8752
rect 6624 8730 6648 8732
rect 6704 8730 6728 8732
rect 6784 8730 6808 8732
rect 6646 8678 6648 8730
rect 6710 8678 6722 8730
rect 6784 8678 6786 8730
rect 6624 8676 6648 8678
rect 6704 8676 6728 8678
rect 6784 8676 6808 8678
rect 6568 8656 6864 8676
rect 6472 8588 6592 8616
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 7886 6500 8434
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6564 7818 6592 8588
rect 6932 8498 6960 8842
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 8090 6684 8366
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6840 8022 6868 8298
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6568 7644 6864 7664
rect 6624 7642 6648 7644
rect 6704 7642 6728 7644
rect 6784 7642 6808 7644
rect 6646 7590 6648 7642
rect 6710 7590 6722 7642
rect 6784 7590 6786 7642
rect 6624 7588 6648 7590
rect 6704 7588 6728 7590
rect 6784 7588 6808 7590
rect 6568 7568 6864 7588
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6472 6458 6500 7482
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 7002 6684 7142
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6840 6644 6868 7414
rect 6918 7304 6974 7313
rect 6918 7239 6920 7248
rect 6972 7239 6974 7248
rect 6920 7210 6972 7216
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6932 6769 6960 6870
rect 6918 6760 6974 6769
rect 6918 6695 6974 6704
rect 6840 6616 6960 6644
rect 6568 6556 6864 6576
rect 6624 6554 6648 6556
rect 6704 6554 6728 6556
rect 6784 6554 6808 6556
rect 6646 6502 6648 6554
rect 6710 6502 6722 6554
rect 6784 6502 6786 6554
rect 6624 6500 6648 6502
rect 6704 6500 6728 6502
rect 6784 6500 6808 6502
rect 6568 6480 6864 6500
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6932 6338 6960 6616
rect 6288 4542 6408 4570
rect 6472 6310 6960 6338
rect 6288 3641 6316 4542
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4214 6408 4422
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6274 3632 6330 3641
rect 6274 3567 6330 3576
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 2650 6316 3470
rect 6380 3058 6408 4150
rect 6472 3505 6500 6310
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6564 5642 6592 6190
rect 6656 5914 6684 6190
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6748 5846 6776 6054
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6568 5468 6864 5488
rect 6624 5466 6648 5468
rect 6704 5466 6728 5468
rect 6784 5466 6808 5468
rect 6646 5414 6648 5466
rect 6710 5414 6722 5466
rect 6784 5414 6786 5466
rect 6624 5412 6648 5414
rect 6704 5412 6728 5414
rect 6784 5412 6808 5414
rect 6568 5392 6864 5412
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6564 4593 6592 4694
rect 6550 4584 6606 4593
rect 6550 4519 6606 4528
rect 6748 4536 6776 5238
rect 6828 5160 6880 5166
rect 6932 5148 6960 5782
rect 6880 5120 6960 5148
rect 6828 5102 6880 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4690 6868 4966
rect 6918 4856 6974 4865
rect 6918 4791 6974 4800
rect 6932 4758 6960 4791
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6920 4548 6972 4554
rect 6748 4508 6920 4536
rect 6920 4490 6972 4496
rect 6568 4380 6864 4400
rect 6624 4378 6648 4380
rect 6704 4378 6728 4380
rect 6784 4378 6808 4380
rect 6646 4326 6648 4378
rect 6710 4326 6722 4378
rect 6784 4326 6786 4378
rect 6624 4324 6648 4326
rect 6704 4324 6728 4326
rect 6784 4324 6808 4326
rect 6568 4304 6864 4324
rect 6552 4140 6604 4146
rect 6932 4128 6960 4490
rect 6604 4100 6960 4128
rect 6552 4082 6604 4088
rect 7024 4060 7052 8570
rect 7116 8430 7144 9454
rect 7208 9450 7236 9862
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9042 7236 9386
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8634 7236 8842
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7194 8528 7250 8537
rect 7194 8463 7250 8472
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7208 7970 7236 8463
rect 7300 8090 7328 11494
rect 7392 11257 7420 11630
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7378 11248 7434 11257
rect 7378 11183 7434 11192
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9518 7420 9862
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7470 9480 7526 9489
rect 7470 9415 7526 9424
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7208 7942 7328 7970
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 6934 7144 7686
rect 7208 7546 7236 7822
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7208 6662 7236 7346
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6322 7236 6598
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 5234 7144 6054
rect 7208 5760 7236 6258
rect 7300 6254 7328 7942
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 6322 7420 7210
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7392 6118 7420 6258
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7288 5772 7340 5778
rect 7208 5732 7288 5760
rect 7288 5714 7340 5720
rect 7194 5400 7250 5409
rect 7194 5335 7250 5344
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6932 4032 7052 4060
rect 6826 3904 6882 3913
rect 6826 3839 6882 3848
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 6460 3392 6512 3398
rect 6840 3380 6868 3839
rect 6932 3448 6960 4032
rect 7116 3942 7144 4422
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7208 3754 7236 5335
rect 7300 4826 7328 5714
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7300 4690 7328 4762
rect 7288 4684 7340 4690
rect 7392 4672 7420 5102
rect 7484 5030 7512 9415
rect 7576 9353 7604 11494
rect 7668 11121 7696 11630
rect 7944 11354 7972 12786
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7654 11112 7710 11121
rect 7654 11047 7710 11056
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7656 9376 7708 9382
rect 7562 9344 7618 9353
rect 7656 9318 7708 9324
rect 7562 9279 7618 9288
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7576 5409 7604 8978
rect 7668 5642 7696 9318
rect 7852 9217 7880 10134
rect 8036 9874 8064 12922
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8220 12714 8248 12854
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8220 12442 8248 12650
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11665 8156 12038
rect 8312 11694 8340 12854
rect 8404 12782 8432 13654
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9048 12782 9076 13398
rect 9692 12986 9720 14818
rect 10309 13084 10605 13104
rect 10365 13082 10389 13084
rect 10445 13082 10469 13084
rect 10525 13082 10549 13084
rect 10387 13030 10389 13082
rect 10451 13030 10463 13082
rect 10525 13030 10527 13082
rect 10365 13028 10389 13030
rect 10445 13028 10469 13030
rect 10525 13028 10549 13030
rect 10309 13008 10605 13028
rect 11164 12986 11192 14818
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 12636 12918 12664 14818
rect 12624 12912 12676 12918
rect 10046 12880 10102 12889
rect 12624 12854 12676 12860
rect 10046 12815 10102 12824
rect 10060 12782 10088 12815
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 8438 12540 8734 12560
rect 8494 12538 8518 12540
rect 8574 12538 8598 12540
rect 8654 12538 8678 12540
rect 8516 12486 8518 12538
rect 8580 12486 8592 12538
rect 8654 12486 8656 12538
rect 8494 12484 8518 12486
rect 8574 12484 8598 12486
rect 8654 12484 8678 12486
rect 8438 12464 8734 12484
rect 8772 12442 8800 12718
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8956 12442 8984 12650
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 11830 8984 12242
rect 9140 11898 9168 12718
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8300 11688 8352 11694
rect 8114 11656 8170 11665
rect 8300 11630 8352 11636
rect 8114 11591 8170 11600
rect 8208 11620 8260 11626
rect 8128 11218 8156 11591
rect 8208 11562 8260 11568
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8220 10810 8248 11562
rect 8438 11452 8734 11472
rect 8494 11450 8518 11452
rect 8574 11450 8598 11452
rect 8654 11450 8678 11452
rect 8516 11398 8518 11450
rect 8580 11398 8592 11450
rect 8654 11398 8656 11450
rect 8494 11396 8518 11398
rect 8574 11396 8598 11398
rect 8654 11396 8678 11398
rect 8438 11376 8734 11396
rect 8956 11286 8984 11766
rect 9140 11694 9168 11834
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8312 10538 8340 11222
rect 8496 10810 8524 11222
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8864 10606 8892 10950
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7944 9846 8064 9874
rect 7838 9208 7894 9217
rect 7838 9143 7894 9152
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7562 5264 7618 5273
rect 7562 5199 7618 5208
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7288 4626 7340 4632
rect 7383 4644 7420 4672
rect 7383 4536 7411 4644
rect 7383 4508 7420 4536
rect 7392 4282 7420 4508
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7288 4208 7340 4214
rect 7484 4196 7512 4762
rect 7576 4264 7604 5199
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4758 7696 4966
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7576 4236 7696 4264
rect 7288 4150 7340 4156
rect 7378 4176 7434 4185
rect 7300 3890 7328 4150
rect 7484 4168 7604 4196
rect 7378 4111 7434 4120
rect 7392 4010 7420 4111
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7300 3862 7420 3890
rect 7116 3726 7236 3754
rect 7288 3732 7340 3738
rect 6932 3420 7052 3448
rect 6840 3352 6960 3380
rect 6460 3334 6512 3340
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6472 2582 6500 3334
rect 6568 3292 6864 3312
rect 6624 3290 6648 3292
rect 6704 3290 6728 3292
rect 6784 3290 6808 3292
rect 6646 3238 6648 3290
rect 6710 3238 6722 3290
rect 6784 3238 6786 3290
rect 6624 3236 6648 3238
rect 6704 3236 6728 3238
rect 6784 3236 6808 3238
rect 6568 3216 6864 3236
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6840 2394 6868 2887
rect 6932 2582 6960 3352
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 6840 2366 6960 2394
rect 6568 2204 6864 2224
rect 6624 2202 6648 2204
rect 6704 2202 6728 2204
rect 6784 2202 6808 2204
rect 6646 2150 6648 2202
rect 6710 2150 6722 2202
rect 6784 2150 6786 2202
rect 6624 2148 6648 2150
rect 6704 2148 6728 2150
rect 6784 2148 6808 2150
rect 6568 2128 6864 2148
rect 6932 2088 6960 2366
rect 6840 2060 6960 2088
rect 6196 1414 6500 1442
rect 6276 1352 6328 1358
rect 6276 1294 6328 1300
rect 6104 870 6224 898
rect 6196 800 6224 870
rect 6288 800 6316 1294
rect 6472 800 6500 1414
rect 6552 1420 6604 1426
rect 6552 1362 6604 1368
rect 6564 800 6592 1362
rect 6734 1320 6790 1329
rect 6734 1255 6790 1264
rect 6748 800 6776 1255
rect 6840 800 6868 2060
rect 7024 2020 7052 3420
rect 6932 1992 7052 2020
rect 6932 800 6960 1992
rect 7116 800 7144 3726
rect 7288 3674 7340 3680
rect 7300 3641 7328 3674
rect 7286 3632 7342 3641
rect 7196 3596 7248 3602
rect 7286 3567 7342 3576
rect 7196 3538 7248 3544
rect 7208 3126 7236 3538
rect 7392 3398 7420 3862
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7470 3496 7526 3505
rect 7470 3431 7526 3440
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7300 3233 7328 3334
rect 7286 3224 7342 3233
rect 7392 3194 7420 3334
rect 7286 3159 7342 3168
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2984 7248 2990
rect 7194 2952 7196 2961
rect 7248 2952 7250 2961
rect 7194 2887 7250 2896
rect 7300 2310 7328 2994
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7194 1864 7250 1873
rect 7194 1799 7250 1808
rect 7208 800 7236 1799
rect 7392 800 7420 2790
rect 7484 800 7512 3431
rect 7576 3194 7604 4168
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7668 3074 7696 4236
rect 7576 3046 7696 3074
rect 7576 800 7604 3046
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7668 2514 7696 2926
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7760 800 7788 8366
rect 7944 7478 7972 9846
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 6458 7880 6734
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5846 7880 6190
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5914 7972 6054
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 4162 7880 5578
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4593 7972 4966
rect 7930 4584 7986 4593
rect 7930 4519 7986 4528
rect 7852 4134 7972 4162
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3534 7880 4014
rect 7944 3738 7972 4134
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7852 3194 7880 3470
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 2825 7972 3470
rect 7930 2816 7986 2825
rect 7930 2751 7986 2760
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7852 800 7880 2518
rect 8036 800 8064 8978
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6458 8156 7142
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 5914 8156 6122
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8220 5250 8248 10066
rect 8312 9178 8340 10474
rect 8438 10364 8734 10384
rect 8494 10362 8518 10364
rect 8574 10362 8598 10364
rect 8654 10362 8678 10364
rect 8516 10310 8518 10362
rect 8580 10310 8592 10362
rect 8654 10310 8656 10362
rect 8494 10308 8518 10310
rect 8574 10308 8598 10310
rect 8654 10308 8678 10310
rect 8438 10288 8734 10308
rect 8956 10130 8984 11222
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9048 10470 9076 11154
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8404 9654 8432 9998
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8680 9674 8708 9930
rect 8392 9648 8444 9654
rect 8680 9646 8800 9674
rect 8392 9590 8444 9596
rect 8438 9276 8734 9296
rect 8494 9274 8518 9276
rect 8574 9274 8598 9276
rect 8654 9274 8678 9276
rect 8516 9222 8518 9274
rect 8580 9222 8592 9274
rect 8654 9222 8656 9274
rect 8494 9220 8518 9222
rect 8574 9220 8598 9222
rect 8654 9220 8678 9222
rect 8438 9200 8734 9220
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8390 9072 8446 9081
rect 8300 9036 8352 9042
rect 8390 9007 8446 9016
rect 8668 9036 8720 9042
rect 8300 8978 8352 8984
rect 8312 8362 8340 8978
rect 8404 8634 8432 9007
rect 8668 8978 8720 8984
rect 8680 8838 8708 8978
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 7993 8340 8298
rect 8438 8188 8734 8208
rect 8494 8186 8518 8188
rect 8574 8186 8598 8188
rect 8654 8186 8678 8188
rect 8516 8134 8518 8186
rect 8580 8134 8592 8186
rect 8654 8134 8656 8186
rect 8494 8132 8518 8134
rect 8574 8132 8598 8134
rect 8654 8132 8678 8134
rect 8438 8112 8734 8132
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8312 7342 8340 7822
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6730 8340 7278
rect 8680 7274 8708 7822
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8438 7100 8734 7120
rect 8494 7098 8518 7100
rect 8574 7098 8598 7100
rect 8654 7098 8678 7100
rect 8516 7046 8518 7098
rect 8580 7046 8592 7098
rect 8654 7046 8656 7098
rect 8494 7044 8518 7046
rect 8574 7044 8598 7046
rect 8654 7044 8678 7046
rect 8438 7024 8734 7044
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8312 5778 8340 6394
rect 8438 6012 8734 6032
rect 8494 6010 8518 6012
rect 8574 6010 8598 6012
rect 8654 6010 8678 6012
rect 8516 5958 8518 6010
rect 8580 5958 8592 6010
rect 8654 5958 8656 6010
rect 8494 5956 8518 5958
rect 8574 5956 8598 5958
rect 8654 5956 8678 5958
rect 8438 5936 8734 5956
rect 8300 5772 8352 5778
rect 8576 5772 8628 5778
rect 8300 5714 8352 5720
rect 8404 5732 8576 5760
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8128 5222 8248 5250
rect 8128 4706 8156 5222
rect 8208 5160 8260 5166
rect 8206 5128 8208 5137
rect 8260 5128 8262 5137
rect 8206 5063 8262 5072
rect 8220 4826 8248 5063
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8128 4678 8248 4706
rect 8114 4584 8170 4593
rect 8114 4519 8170 4528
rect 8128 4078 8156 4519
rect 8116 4072 8168 4078
rect 8114 4040 8116 4049
rect 8168 4040 8170 4049
rect 8114 3975 8170 3984
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3534 8156 3878
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8114 3360 8170 3369
rect 8114 3295 8170 3304
rect 8128 800 8156 3295
rect 8220 800 8248 4678
rect 8312 4264 8340 5510
rect 8404 5166 8432 5732
rect 8576 5714 8628 5720
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8438 4924 8734 4944
rect 8494 4922 8518 4924
rect 8574 4922 8598 4924
rect 8654 4922 8678 4924
rect 8516 4870 8518 4922
rect 8580 4870 8592 4922
rect 8654 4870 8656 4922
rect 8494 4868 8518 4870
rect 8574 4868 8598 4870
rect 8654 4868 8678 4870
rect 8438 4848 8734 4868
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4321 8616 4422
rect 8574 4312 8630 4321
rect 8312 4236 8432 4264
rect 8574 4247 8630 4256
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8312 3505 8340 4082
rect 8404 4078 8432 4236
rect 8666 4176 8722 4185
rect 8666 4111 8722 4120
rect 8680 4078 8708 4111
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8438 3836 8734 3856
rect 8494 3834 8518 3836
rect 8574 3834 8598 3836
rect 8654 3834 8678 3836
rect 8516 3782 8518 3834
rect 8580 3782 8592 3834
rect 8654 3782 8656 3834
rect 8494 3780 8518 3782
rect 8574 3780 8598 3782
rect 8654 3780 8678 3782
rect 8438 3760 8734 3780
rect 8772 3618 8800 9646
rect 8864 7936 8892 9998
rect 8956 9722 8984 10066
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9048 9518 9076 10406
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8956 8634 8984 8978
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8864 7908 8984 7936
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8864 7002 8892 7754
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8956 6474 8984 7908
rect 9048 7886 9076 8774
rect 9140 8106 9168 9862
rect 9232 9654 9260 12378
rect 9324 12306 9352 12582
rect 10980 12434 11008 12718
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 9876 12406 10180 12434
rect 10980 12406 11100 12434
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9588 12232 9640 12238
rect 9784 12209 9812 12310
rect 9876 12306 9904 12406
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9956 12232 10008 12238
rect 9588 12174 9640 12180
rect 9770 12200 9826 12209
rect 9416 11898 9444 12174
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11898 9536 12038
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9416 10130 9444 11834
rect 9600 11626 9628 12174
rect 9956 12174 10008 12180
rect 9770 12135 9826 12144
rect 9680 11688 9732 11694
rect 9968 11665 9996 12174
rect 9680 11630 9732 11636
rect 9954 11656 10010 11665
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9692 11354 9720 11630
rect 9954 11591 10010 11600
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 10736 9732 10742
rect 9678 10704 9680 10713
rect 9732 10704 9734 10713
rect 9678 10639 9734 10648
rect 9784 10538 9812 11086
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10742 9904 11018
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9494 10432 9550 10441
rect 9494 10367 9550 10376
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 9178 9444 9318
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 8430 9260 8910
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9140 8078 9260 8106
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 6866 9076 7686
rect 9140 7002 9168 7890
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8956 6446 9076 6474
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8956 5846 8984 6122
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8942 5264 8998 5273
rect 8942 5199 8998 5208
rect 8956 5166 8984 5199
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8588 3590 8800 3618
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8404 2990 8432 3334
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8588 2836 8616 3590
rect 8668 3528 8720 3534
rect 8720 3476 8800 3482
rect 8668 3470 8800 3476
rect 8680 3454 8800 3470
rect 8666 3224 8722 3233
rect 8666 3159 8722 3168
rect 8680 2922 8708 3159
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8312 2808 8616 2836
rect 8312 2428 8340 2808
rect 8438 2748 8734 2768
rect 8494 2746 8518 2748
rect 8574 2746 8598 2748
rect 8654 2746 8678 2748
rect 8516 2694 8518 2746
rect 8580 2694 8592 2746
rect 8654 2694 8656 2746
rect 8494 2692 8518 2694
rect 8574 2692 8598 2694
rect 8654 2692 8678 2694
rect 8438 2672 8734 2692
rect 8772 2650 8800 3454
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8392 2576 8444 2582
rect 8390 2544 8392 2553
rect 8444 2544 8446 2553
rect 8390 2479 8446 2488
rect 8312 2400 8432 2428
rect 8404 800 8432 2400
rect 8666 2408 8722 2417
rect 8666 2343 8722 2352
rect 8864 2360 8892 4082
rect 8956 4078 8984 4422
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8956 3505 8984 3606
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8956 2514 8984 2790
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8482 1592 8538 1601
rect 8482 1527 8538 1536
rect 8496 800 8524 1527
rect 8680 800 8708 2343
rect 8864 2332 8984 2360
rect 8850 2272 8906 2281
rect 8850 2207 8906 2216
rect 8758 2000 8814 2009
rect 8758 1935 8814 1944
rect 8772 800 8800 1935
rect 8864 800 8892 2207
rect 8956 1222 8984 2332
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 9048 800 9076 6446
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5370 9168 5714
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9140 3738 9168 5034
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9140 2990 9168 3402
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9232 2582 9260 8078
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7342 9352 7686
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 5234 9352 6734
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4622 9352 5170
rect 9312 4616 9364 4622
rect 9310 4584 9312 4593
rect 9364 4584 9366 4593
rect 9310 4519 9366 4528
rect 9312 4208 9364 4214
rect 9310 4176 9312 4185
rect 9364 4176 9366 4185
rect 9310 4111 9366 4120
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9324 2446 9352 3975
rect 9416 3856 9444 7958
rect 9508 6905 9536 10367
rect 9600 9058 9628 10474
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10146 9720 10406
rect 9784 10266 9812 10474
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9876 10198 9904 10678
rect 9864 10192 9916 10198
rect 9692 10118 9812 10146
rect 9864 10134 9916 10140
rect 9784 10044 9812 10118
rect 9864 10056 9916 10062
rect 9784 10016 9864 10044
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9382 9720 9862
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9600 9030 9720 9058
rect 9692 7936 9720 9030
rect 9784 8634 9812 10016
rect 9968 10033 9996 11494
rect 10060 11354 10088 12242
rect 10152 11914 10180 12406
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10309 11996 10605 12016
rect 10365 11994 10389 11996
rect 10445 11994 10469 11996
rect 10525 11994 10549 11996
rect 10387 11942 10389 11994
rect 10451 11942 10463 11994
rect 10525 11942 10527 11994
rect 10365 11940 10389 11942
rect 10445 11940 10469 11942
rect 10525 11940 10549 11942
rect 10309 11920 10605 11940
rect 10152 11898 10272 11914
rect 10152 11892 10284 11898
rect 10152 11886 10232 11892
rect 10232 11834 10284 11840
rect 10796 11762 10824 12038
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10416 11688 10468 11694
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 10414 11656 10416 11665
rect 10468 11656 10470 11665
rect 10414 11591 10470 11600
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 10282 10088 11018
rect 10152 10418 10180 11086
rect 10244 10713 10272 11591
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10336 11218 10364 11290
rect 10428 11286 10456 11591
rect 10520 11286 10548 11698
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10309 10908 10605 10928
rect 10365 10906 10389 10908
rect 10445 10906 10469 10908
rect 10525 10906 10549 10908
rect 10387 10854 10389 10906
rect 10451 10854 10463 10906
rect 10525 10854 10527 10906
rect 10365 10852 10389 10854
rect 10445 10852 10469 10854
rect 10525 10852 10549 10854
rect 10309 10832 10605 10852
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10244 10606 10272 10639
rect 10232 10600 10284 10606
rect 10284 10560 10364 10588
rect 10232 10542 10284 10548
rect 10152 10390 10272 10418
rect 10060 10254 10180 10282
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9864 9998 9916 10004
rect 9954 10024 10010 10033
rect 9954 9959 10010 9968
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9586 9996 9862
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9450 9996 9522
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9600 7908 9720 7936
rect 9600 7002 9628 7908
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7478 9720 7754
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9692 6934 9720 7414
rect 9680 6928 9732 6934
rect 9494 6896 9550 6905
rect 9680 6870 9732 6876
rect 9494 6831 9550 6840
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 5302 9536 5714
rect 9600 5642 9628 6054
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9600 4758 9628 5578
rect 9692 5574 9720 6870
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 4752 9640 4758
rect 9494 4720 9550 4729
rect 9588 4694 9640 4700
rect 9494 4655 9496 4664
rect 9548 4655 9550 4664
rect 9496 4626 9548 4632
rect 9692 4486 9720 5170
rect 9496 4480 9548 4486
rect 9680 4480 9732 4486
rect 9496 4422 9548 4428
rect 9586 4448 9642 4457
rect 9508 4282 9536 4422
rect 9680 4422 9732 4428
rect 9586 4383 9642 4392
rect 9600 4282 9628 4383
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9416 3828 9536 3856
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9416 3194 9444 3674
rect 9508 3670 9536 3828
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 800 9168 2246
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9324 800 9352 1362
rect 9416 800 9444 2790
rect 9508 800 9536 2994
rect 9600 2650 9628 4111
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3777 9720 3878
rect 9678 3768 9734 3777
rect 9678 3703 9734 3712
rect 9784 3670 9812 8366
rect 9968 8242 9996 8842
rect 10060 8498 10088 10134
rect 10152 9704 10180 10254
rect 10244 9994 10272 10390
rect 10336 10198 10364 10560
rect 10508 10464 10560 10470
rect 10506 10432 10508 10441
rect 10560 10432 10562 10441
rect 10506 10367 10562 10376
rect 10704 10266 10732 11018
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10538 10824 10950
rect 10888 10810 10916 11154
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10309 9820 10605 9840
rect 10365 9818 10389 9820
rect 10445 9818 10469 9820
rect 10525 9818 10549 9820
rect 10387 9766 10389 9818
rect 10451 9766 10463 9818
rect 10525 9766 10527 9818
rect 10365 9764 10389 9766
rect 10445 9764 10469 9766
rect 10525 9764 10549 9766
rect 10309 9744 10605 9764
rect 10232 9716 10284 9722
rect 10152 9676 10232 9704
rect 10232 9658 10284 9664
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10152 9042 10180 9386
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9876 8214 9996 8242
rect 9876 7410 9904 8214
rect 9954 8120 10010 8129
rect 9954 8055 9956 8064
rect 10008 8055 10010 8064
rect 9956 8026 10008 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6798 9904 7210
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9876 5370 9904 5714
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9862 5128 9918 5137
rect 9862 5063 9864 5072
rect 9916 5063 9918 5072
rect 9864 5034 9916 5040
rect 9968 4570 9996 7822
rect 10060 7546 10088 7958
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10060 7002 10088 7482
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5234 10088 6258
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10152 5114 10180 8842
rect 10244 8838 10272 9658
rect 10704 9450 10732 10202
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9722 10916 10066
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10796 8922 10824 9454
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10704 8894 10824 8922
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10309 8732 10605 8752
rect 10365 8730 10389 8732
rect 10445 8730 10469 8732
rect 10525 8730 10549 8732
rect 10387 8678 10389 8730
rect 10451 8678 10463 8730
rect 10525 8678 10527 8730
rect 10365 8676 10389 8678
rect 10445 8676 10469 8678
rect 10525 8676 10549 8678
rect 10309 8656 10605 8676
rect 10232 8424 10284 8430
rect 10284 8372 10364 8378
rect 10232 8366 10364 8372
rect 10244 8350 10364 8366
rect 10336 7886 10364 8350
rect 10704 8106 10732 8894
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8498 10824 8774
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10888 8378 10916 9318
rect 10796 8350 10916 8378
rect 10796 8129 10824 8350
rect 10980 8242 11008 11494
rect 11072 8634 11100 12406
rect 11164 11694 11192 12650
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11256 11898 11284 12135
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11532 11694 11560 12582
rect 11624 12442 11652 12650
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 12306 11652 12378
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11152 11688 11204 11694
rect 11520 11688 11572 11694
rect 11152 11630 11204 11636
rect 11242 11656 11298 11665
rect 11164 10606 11192 11630
rect 11520 11630 11572 11636
rect 11242 11591 11298 11600
rect 11256 11218 11284 11591
rect 11532 11218 11560 11630
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11256 10810 11284 11154
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11256 10538 11284 10746
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11348 10198 11376 10950
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8566 11192 8978
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8634 11284 8910
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10980 8214 11192 8242
rect 10612 8078 10732 8106
rect 10782 8120 10838 8129
rect 10612 7993 10640 8078
rect 10782 8055 10838 8064
rect 10692 8016 10744 8022
rect 10598 7984 10654 7993
rect 10692 7958 10744 7964
rect 10598 7919 10654 7928
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 5710 10272 7686
rect 10309 7644 10605 7664
rect 10365 7642 10389 7644
rect 10445 7642 10469 7644
rect 10525 7642 10549 7644
rect 10387 7590 10389 7642
rect 10451 7590 10463 7642
rect 10525 7590 10527 7642
rect 10365 7588 10389 7590
rect 10445 7588 10469 7590
rect 10525 7588 10549 7590
rect 10309 7568 10605 7588
rect 10704 7546 10732 7958
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10876 7336 10928 7342
rect 10980 7324 11008 7686
rect 11072 7342 11100 7890
rect 10928 7296 11008 7324
rect 11060 7336 11112 7342
rect 10876 7278 10928 7284
rect 11060 7278 11112 7284
rect 10336 7002 10364 7278
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10428 6798 10456 7278
rect 10888 7002 10916 7278
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11164 6882 11192 8214
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11072 6854 11192 6882
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10309 6556 10605 6576
rect 10365 6554 10389 6556
rect 10445 6554 10469 6556
rect 10525 6554 10549 6556
rect 10387 6502 10389 6554
rect 10451 6502 10463 6554
rect 10525 6502 10527 6554
rect 10365 6500 10389 6502
rect 10445 6500 10469 6502
rect 10525 6500 10549 6502
rect 10309 6480 10605 6500
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5914 10732 6122
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5778 10824 6598
rect 11072 6458 11100 6854
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10309 5468 10605 5488
rect 10365 5466 10389 5468
rect 10445 5466 10469 5468
rect 10525 5466 10549 5468
rect 10387 5414 10389 5466
rect 10451 5414 10463 5466
rect 10525 5414 10527 5466
rect 10365 5412 10389 5414
rect 10445 5412 10469 5414
rect 10525 5412 10549 5414
rect 10309 5392 10605 5412
rect 10704 5166 10732 5510
rect 9876 4542 9996 4570
rect 10060 5086 10180 5114
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 9876 3738 9904 4542
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9600 1426 9628 2246
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9692 800 9720 3470
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 800 9812 3402
rect 9864 2984 9916 2990
rect 9862 2952 9864 2961
rect 9916 2952 9918 2961
rect 9862 2887 9918 2896
rect 9968 800 9996 4422
rect 10060 4078 10088 5086
rect 10244 4826 10272 5102
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10336 4468 10364 5034
rect 10598 4992 10654 5001
rect 10598 4927 10654 4936
rect 10612 4826 10640 4927
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10152 4440 10364 4468
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 2514 10088 3878
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 10060 1358 10088 2314
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10046 1184 10102 1193
rect 10046 1119 10102 1128
rect 10060 800 10088 1119
rect 10152 800 10180 4440
rect 10309 4380 10605 4400
rect 10365 4378 10389 4380
rect 10445 4378 10469 4380
rect 10525 4378 10549 4380
rect 10387 4326 10389 4378
rect 10451 4326 10463 4378
rect 10525 4326 10527 4378
rect 10365 4324 10389 4326
rect 10445 4324 10469 4326
rect 10525 4324 10549 4326
rect 10309 4304 10605 4324
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10322 4040 10378 4049
rect 10232 4004 10284 4010
rect 10322 3975 10378 3984
rect 10232 3946 10284 3952
rect 10244 2514 10272 3946
rect 10336 3670 10364 3975
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10309 3292 10605 3312
rect 10365 3290 10389 3292
rect 10445 3290 10469 3292
rect 10525 3290 10549 3292
rect 10387 3238 10389 3290
rect 10451 3238 10463 3290
rect 10525 3238 10527 3290
rect 10365 3236 10389 3238
rect 10445 3236 10469 3238
rect 10525 3236 10549 3238
rect 10309 3216 10605 3236
rect 10704 2990 10732 4150
rect 10796 3602 10824 5578
rect 10888 4758 10916 5578
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10980 5137 11008 5510
rect 10966 5128 11022 5137
rect 10966 5063 11022 5072
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10876 4616 10928 4622
rect 11072 4604 11100 6054
rect 10928 4576 11100 4604
rect 10876 4558 10928 4564
rect 10874 4176 10930 4185
rect 10874 4111 10930 4120
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10888 3074 10916 4111
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10796 3046 10916 3074
rect 10966 3088 11022 3097
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10796 2774 10824 3046
rect 10966 3023 11022 3032
rect 10980 2922 11008 3023
rect 11072 2990 11100 3402
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10796 2746 11008 2774
rect 10980 2582 11008 2746
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10309 2204 10605 2224
rect 10365 2202 10389 2204
rect 10445 2202 10469 2204
rect 10525 2202 10549 2204
rect 10387 2150 10389 2202
rect 10451 2150 10463 2202
rect 10525 2150 10527 2202
rect 10365 2148 10389 2150
rect 10445 2148 10469 2150
rect 10525 2148 10549 2150
rect 10309 2128 10605 2148
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10336 800 10364 1294
rect 10416 1216 10468 1222
rect 10704 1170 10732 2246
rect 10416 1158 10468 1164
rect 10428 800 10456 1158
rect 10612 1142 10732 1170
rect 10612 800 10640 1142
rect 10692 1080 10744 1086
rect 10692 1022 10744 1028
rect 10704 800 10732 1022
rect 10796 800 10824 2382
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 1086 10916 2246
rect 10876 1080 10928 1086
rect 10876 1022 10928 1028
rect 10980 800 11008 2314
rect 11072 800 11100 2790
rect 11164 2582 11192 6734
rect 11256 6322 11284 7278
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11256 4010 11284 5782
rect 11348 4758 11376 8774
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11440 3670 11468 7278
rect 11532 5166 11560 9454
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11624 4706 11652 6598
rect 11532 4678 11652 4706
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11334 3224 11390 3233
rect 11334 3159 11390 3168
rect 11242 2816 11298 2825
rect 11242 2751 11298 2760
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11256 800 11284 2751
rect 11348 800 11376 3159
rect 11440 800 11468 3402
rect 11532 2582 11560 4678
rect 11716 4078 11744 8774
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5710 11836 6054
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11900 4078 11928 8366
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 4214 12020 7686
rect 11980 4208 12032 4214
rect 12084 4185 12112 9454
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11980 4150 12032 4156
rect 12070 4176 12126 4185
rect 12070 4111 12126 4120
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11624 3233 11652 3606
rect 11610 3224 11666 3233
rect 11610 3159 11666 3168
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11624 800 11652 2994
rect 11716 800 11744 3878
rect 11794 3632 11850 3641
rect 11794 3567 11796 3576
rect 11848 3567 11850 3576
rect 11796 3538 11848 3544
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11808 2825 11836 2994
rect 11794 2816 11850 2825
rect 11794 2751 11850 2760
rect 11900 800 11928 3470
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11992 800 12020 3062
rect 12084 800 12112 3946
rect 12176 2922 12204 4218
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12268 800 12296 3674
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12360 800 12388 3130
rect 12452 2514 12480 7346
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12544 800 12572 4490
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 800 12664 4082
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12728 800 12756 3606
rect 12912 800 12940 4422
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13004 800 13032 2790
rect 13188 800 13216 3334
rect 13280 800 13308 5034
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 386 0 442 800
rect 478 0 534 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
<< via2 >>
rect 478 10104 534 10160
rect 570 7792 626 7848
rect 754 3984 810 4040
rect 938 2760 994 2816
rect 1398 8880 1454 8936
rect 1398 5636 1454 5672
rect 1398 5616 1400 5636
rect 1400 5616 1452 5636
rect 1452 5616 1454 5636
rect 1766 10240 1822 10296
rect 2318 9696 2374 9752
rect 2226 8472 2282 8528
rect 2134 6060 2136 6080
rect 2136 6060 2188 6080
rect 2188 6060 2190 6080
rect 2134 6024 2190 6060
rect 2042 2760 2098 2816
rect 2410 6296 2466 6352
rect 2826 13082 2882 13084
rect 2906 13082 2962 13084
rect 2986 13082 3042 13084
rect 3066 13082 3122 13084
rect 2826 13030 2852 13082
rect 2852 13030 2882 13082
rect 2906 13030 2916 13082
rect 2916 13030 2962 13082
rect 2986 13030 3032 13082
rect 3032 13030 3042 13082
rect 3066 13030 3096 13082
rect 3096 13030 3122 13082
rect 2826 13028 2882 13030
rect 2906 13028 2962 13030
rect 2986 13028 3042 13030
rect 3066 13028 3122 13030
rect 2826 11994 2882 11996
rect 2906 11994 2962 11996
rect 2986 11994 3042 11996
rect 3066 11994 3122 11996
rect 2826 11942 2852 11994
rect 2852 11942 2882 11994
rect 2906 11942 2916 11994
rect 2916 11942 2962 11994
rect 2986 11942 3032 11994
rect 3032 11942 3042 11994
rect 3066 11942 3096 11994
rect 3096 11942 3122 11994
rect 2826 11940 2882 11942
rect 2906 11940 2962 11942
rect 2986 11940 3042 11942
rect 3066 11940 3122 11942
rect 3054 11600 3110 11656
rect 2826 10906 2882 10908
rect 2906 10906 2962 10908
rect 2986 10906 3042 10908
rect 3066 10906 3122 10908
rect 2826 10854 2852 10906
rect 2852 10854 2882 10906
rect 2906 10854 2916 10906
rect 2916 10854 2962 10906
rect 2986 10854 3032 10906
rect 3032 10854 3042 10906
rect 3066 10854 3096 10906
rect 3096 10854 3122 10906
rect 2826 10852 2882 10854
rect 2906 10852 2962 10854
rect 2986 10852 3042 10854
rect 3066 10852 3122 10854
rect 2778 10684 2780 10704
rect 2780 10684 2832 10704
rect 2832 10684 2834 10704
rect 2778 10648 2834 10684
rect 2778 10376 2834 10432
rect 3238 10240 3294 10296
rect 3422 10124 3478 10160
rect 3422 10104 3424 10124
rect 3424 10104 3476 10124
rect 3476 10104 3478 10124
rect 4697 12538 4753 12540
rect 4777 12538 4833 12540
rect 4857 12538 4913 12540
rect 4937 12538 4993 12540
rect 4697 12486 4723 12538
rect 4723 12486 4753 12538
rect 4777 12486 4787 12538
rect 4787 12486 4833 12538
rect 4857 12486 4903 12538
rect 4903 12486 4913 12538
rect 4937 12486 4967 12538
rect 4967 12486 4993 12538
rect 4697 12484 4753 12486
rect 4777 12484 4833 12486
rect 4857 12484 4913 12486
rect 4937 12484 4993 12486
rect 5078 11756 5134 11792
rect 5078 11736 5080 11756
rect 5080 11736 5132 11756
rect 5132 11736 5134 11756
rect 3698 10376 3754 10432
rect 3606 10104 3662 10160
rect 2826 9818 2882 9820
rect 2906 9818 2962 9820
rect 2986 9818 3042 9820
rect 3066 9818 3122 9820
rect 2826 9766 2852 9818
rect 2852 9766 2882 9818
rect 2906 9766 2916 9818
rect 2916 9766 2962 9818
rect 2986 9766 3032 9818
rect 3032 9766 3042 9818
rect 3066 9766 3096 9818
rect 3096 9766 3122 9818
rect 2826 9764 2882 9766
rect 2906 9764 2962 9766
rect 2986 9764 3042 9766
rect 3066 9764 3122 9766
rect 3330 9832 3386 9888
rect 3238 9152 3294 9208
rect 2826 8730 2882 8732
rect 2906 8730 2962 8732
rect 2986 8730 3042 8732
rect 3066 8730 3122 8732
rect 2826 8678 2852 8730
rect 2852 8678 2882 8730
rect 2906 8678 2916 8730
rect 2916 8678 2962 8730
rect 2986 8678 3032 8730
rect 3032 8678 3042 8730
rect 3066 8678 3096 8730
rect 3096 8678 3122 8730
rect 2826 8676 2882 8678
rect 2906 8676 2962 8678
rect 2986 8676 3042 8678
rect 3066 8676 3122 8678
rect 2826 7642 2882 7644
rect 2906 7642 2962 7644
rect 2986 7642 3042 7644
rect 3066 7642 3122 7644
rect 2826 7590 2852 7642
rect 2852 7590 2882 7642
rect 2906 7590 2916 7642
rect 2916 7590 2962 7642
rect 2986 7590 3032 7642
rect 3032 7590 3042 7642
rect 3066 7590 3096 7642
rect 3096 7590 3122 7642
rect 2826 7588 2882 7590
rect 2906 7588 2962 7590
rect 2986 7588 3042 7590
rect 3066 7588 3122 7590
rect 2778 6704 2834 6760
rect 3054 6704 3110 6760
rect 2826 6554 2882 6556
rect 2906 6554 2962 6556
rect 2986 6554 3042 6556
rect 3066 6554 3122 6556
rect 2826 6502 2852 6554
rect 2852 6502 2882 6554
rect 2906 6502 2916 6554
rect 2916 6502 2962 6554
rect 2986 6502 3032 6554
rect 3032 6502 3042 6554
rect 3066 6502 3096 6554
rect 3096 6502 3122 6554
rect 2826 6500 2882 6502
rect 2906 6500 2962 6502
rect 2986 6500 3042 6502
rect 3066 6500 3122 6502
rect 3238 6568 3294 6624
rect 2318 3576 2374 3632
rect 2318 3440 2374 3496
rect 2826 5466 2882 5468
rect 2906 5466 2962 5468
rect 2986 5466 3042 5468
rect 3066 5466 3122 5468
rect 2826 5414 2852 5466
rect 2852 5414 2882 5466
rect 2906 5414 2916 5466
rect 2916 5414 2962 5466
rect 2986 5414 3032 5466
rect 3032 5414 3042 5466
rect 3066 5414 3096 5466
rect 3096 5414 3122 5466
rect 2826 5412 2882 5414
rect 2906 5412 2962 5414
rect 2986 5412 3042 5414
rect 3066 5412 3122 5414
rect 2686 4800 2742 4856
rect 2826 4378 2882 4380
rect 2906 4378 2962 4380
rect 2986 4378 3042 4380
rect 3066 4378 3122 4380
rect 2826 4326 2852 4378
rect 2852 4326 2882 4378
rect 2906 4326 2916 4378
rect 2916 4326 2962 4378
rect 2986 4326 3032 4378
rect 3032 4326 3042 4378
rect 3066 4326 3096 4378
rect 3096 4326 3122 4378
rect 2826 4324 2882 4326
rect 2906 4324 2962 4326
rect 2986 4324 3042 4326
rect 3066 4324 3122 4326
rect 3422 4800 3478 4856
rect 3054 3440 3110 3496
rect 2826 3290 2882 3292
rect 2906 3290 2962 3292
rect 2986 3290 3042 3292
rect 3066 3290 3122 3292
rect 2826 3238 2852 3290
rect 2852 3238 2882 3290
rect 2906 3238 2916 3290
rect 2916 3238 2962 3290
rect 2986 3238 3032 3290
rect 3032 3238 3042 3290
rect 3066 3238 3096 3290
rect 3096 3238 3122 3290
rect 2826 3236 2882 3238
rect 2906 3236 2962 3238
rect 2986 3236 3042 3238
rect 3066 3236 3122 3238
rect 3054 3052 3110 3088
rect 3054 3032 3056 3052
rect 3056 3032 3108 3052
rect 3108 3032 3110 3052
rect 3146 2932 3148 2952
rect 3148 2932 3200 2952
rect 3200 2932 3202 2952
rect 3146 2896 3202 2932
rect 3054 2624 3110 2680
rect 2826 2202 2882 2204
rect 2906 2202 2962 2204
rect 2986 2202 3042 2204
rect 3066 2202 3122 2204
rect 2826 2150 2852 2202
rect 2852 2150 2882 2202
rect 2906 2150 2916 2202
rect 2916 2150 2962 2202
rect 2986 2150 3032 2202
rect 3032 2150 3042 2202
rect 3066 2150 3096 2202
rect 3096 2150 3122 2202
rect 2826 2148 2882 2150
rect 2906 2148 2962 2150
rect 2986 2148 3042 2150
rect 3066 2148 3122 2150
rect 3606 6840 3662 6896
rect 3974 9152 4030 9208
rect 3882 8472 3938 8528
rect 3882 8064 3938 8120
rect 3974 5208 4030 5264
rect 3698 3848 3754 3904
rect 3974 4528 4030 4584
rect 3330 2488 3386 2544
rect 4066 3712 4122 3768
rect 3698 2896 3754 2952
rect 3974 3340 3976 3360
rect 3976 3340 4028 3360
rect 4028 3340 4030 3360
rect 3974 3304 4030 3340
rect 3698 1264 3754 1320
rect 4158 3052 4214 3088
rect 4158 3032 4160 3052
rect 4160 3032 4212 3052
rect 4212 3032 4214 3052
rect 4434 10240 4490 10296
rect 4697 11450 4753 11452
rect 4777 11450 4833 11452
rect 4857 11450 4913 11452
rect 4937 11450 4993 11452
rect 4697 11398 4723 11450
rect 4723 11398 4753 11450
rect 4777 11398 4787 11450
rect 4787 11398 4833 11450
rect 4857 11398 4903 11450
rect 4903 11398 4913 11450
rect 4937 11398 4967 11450
rect 4967 11398 4993 11450
rect 4697 11396 4753 11398
rect 4777 11396 4833 11398
rect 4857 11396 4913 11398
rect 4937 11396 4993 11398
rect 6568 13082 6624 13084
rect 6648 13082 6704 13084
rect 6728 13082 6784 13084
rect 6808 13082 6864 13084
rect 6568 13030 6594 13082
rect 6594 13030 6624 13082
rect 6648 13030 6658 13082
rect 6658 13030 6704 13082
rect 6728 13030 6774 13082
rect 6774 13030 6784 13082
rect 6808 13030 6838 13082
rect 6838 13030 6864 13082
rect 6568 13028 6624 13030
rect 6648 13028 6704 13030
rect 6728 13028 6784 13030
rect 6808 13028 6864 13030
rect 4618 10784 4674 10840
rect 4802 10648 4858 10704
rect 4710 10512 4766 10568
rect 4894 10512 4950 10568
rect 4697 10362 4753 10364
rect 4777 10362 4833 10364
rect 4857 10362 4913 10364
rect 4937 10362 4993 10364
rect 4697 10310 4723 10362
rect 4723 10310 4753 10362
rect 4777 10310 4787 10362
rect 4787 10310 4833 10362
rect 4857 10310 4903 10362
rect 4903 10310 4913 10362
rect 4937 10310 4967 10362
rect 4967 10310 4993 10362
rect 4697 10308 4753 10310
rect 4777 10308 4833 10310
rect 4857 10308 4913 10310
rect 4937 10308 4993 10310
rect 5170 10240 5226 10296
rect 4710 9868 4712 9888
rect 4712 9868 4764 9888
rect 4764 9868 4766 9888
rect 4710 9832 4766 9868
rect 4986 9832 5042 9888
rect 5078 9560 5134 9616
rect 4894 9424 4950 9480
rect 4697 9274 4753 9276
rect 4777 9274 4833 9276
rect 4857 9274 4913 9276
rect 4937 9274 4993 9276
rect 4697 9222 4723 9274
rect 4723 9222 4753 9274
rect 4777 9222 4787 9274
rect 4787 9222 4833 9274
rect 4857 9222 4903 9274
rect 4903 9222 4913 9274
rect 4937 9222 4967 9274
rect 4967 9222 4993 9274
rect 4697 9220 4753 9222
rect 4777 9220 4833 9222
rect 4857 9220 4913 9222
rect 4937 9220 4993 9222
rect 5078 9152 5134 9208
rect 4802 9052 4804 9072
rect 4804 9052 4856 9072
rect 4856 9052 4858 9072
rect 4802 9016 4858 9052
rect 4986 9016 5042 9072
rect 4710 8880 4766 8936
rect 4434 5888 4490 5944
rect 4342 4528 4398 4584
rect 4066 2216 4122 2272
rect 4250 1128 4306 1184
rect 4434 3712 4490 3768
rect 4697 8186 4753 8188
rect 4777 8186 4833 8188
rect 4857 8186 4913 8188
rect 4937 8186 4993 8188
rect 4697 8134 4723 8186
rect 4723 8134 4753 8186
rect 4777 8134 4787 8186
rect 4787 8134 4833 8186
rect 4857 8134 4903 8186
rect 4903 8134 4913 8186
rect 4937 8134 4967 8186
rect 4967 8134 4993 8186
rect 4697 8132 4753 8134
rect 4777 8132 4833 8134
rect 4857 8132 4913 8134
rect 4937 8132 4993 8134
rect 5078 7540 5134 7576
rect 5078 7520 5080 7540
rect 5080 7520 5132 7540
rect 5132 7520 5134 7540
rect 4697 7098 4753 7100
rect 4777 7098 4833 7100
rect 4857 7098 4913 7100
rect 4937 7098 4993 7100
rect 4697 7046 4723 7098
rect 4723 7046 4753 7098
rect 4777 7046 4787 7098
rect 4787 7046 4833 7098
rect 4857 7046 4903 7098
rect 4903 7046 4913 7098
rect 4937 7046 4967 7098
rect 4967 7046 4993 7098
rect 4697 7044 4753 7046
rect 4777 7044 4833 7046
rect 4857 7044 4913 7046
rect 4937 7044 4993 7046
rect 4618 6704 4674 6760
rect 4710 6160 4766 6216
rect 4697 6010 4753 6012
rect 4777 6010 4833 6012
rect 4857 6010 4913 6012
rect 4937 6010 4993 6012
rect 4697 5958 4723 6010
rect 4723 5958 4753 6010
rect 4777 5958 4787 6010
rect 4787 5958 4833 6010
rect 4857 5958 4903 6010
rect 4903 5958 4913 6010
rect 4937 5958 4967 6010
rect 4967 5958 4993 6010
rect 4697 5956 4753 5958
rect 4777 5956 4833 5958
rect 4857 5956 4913 5958
rect 4937 5956 4993 5958
rect 5630 11348 5686 11384
rect 5630 11328 5632 11348
rect 5632 11328 5684 11348
rect 5684 11328 5686 11348
rect 5630 11212 5686 11248
rect 5630 11192 5632 11212
rect 5632 11192 5684 11212
rect 5684 11192 5686 11212
rect 5722 11056 5778 11112
rect 5630 10920 5686 10976
rect 5446 10376 5502 10432
rect 5538 9560 5594 9616
rect 5354 9288 5410 9344
rect 5538 9152 5594 9208
rect 5630 8336 5686 8392
rect 5262 6860 5318 6896
rect 5262 6840 5264 6860
rect 5264 6840 5316 6860
rect 5316 6840 5318 6860
rect 4526 2896 4582 2952
rect 4434 2488 4490 2544
rect 4697 4922 4753 4924
rect 4777 4922 4833 4924
rect 4857 4922 4913 4924
rect 4937 4922 4993 4924
rect 4697 4870 4723 4922
rect 4723 4870 4753 4922
rect 4777 4870 4787 4922
rect 4787 4870 4833 4922
rect 4857 4870 4903 4922
rect 4903 4870 4913 4922
rect 4937 4870 4967 4922
rect 4967 4870 4993 4922
rect 4697 4868 4753 4870
rect 4777 4868 4833 4870
rect 4857 4868 4913 4870
rect 4937 4868 4993 4870
rect 4894 3984 4950 4040
rect 4697 3834 4753 3836
rect 4777 3834 4833 3836
rect 4857 3834 4913 3836
rect 4937 3834 4993 3836
rect 4697 3782 4723 3834
rect 4723 3782 4753 3834
rect 4777 3782 4787 3834
rect 4787 3782 4833 3834
rect 4857 3782 4903 3834
rect 4903 3782 4913 3834
rect 4937 3782 4967 3834
rect 4967 3782 4993 3834
rect 4697 3780 4753 3782
rect 4777 3780 4833 3782
rect 4857 3780 4913 3782
rect 4937 3780 4993 3782
rect 5446 6568 5502 6624
rect 5446 4936 5502 4992
rect 5446 4800 5502 4856
rect 4710 3576 4766 3632
rect 4894 3596 4950 3632
rect 4894 3576 4896 3596
rect 4896 3576 4948 3596
rect 4948 3576 4950 3596
rect 4802 3052 4858 3088
rect 4802 3032 4804 3052
rect 4804 3032 4856 3052
rect 4856 3032 4858 3052
rect 4697 2746 4753 2748
rect 4777 2746 4833 2748
rect 4857 2746 4913 2748
rect 4937 2746 4993 2748
rect 4697 2694 4723 2746
rect 4723 2694 4753 2746
rect 4777 2694 4787 2746
rect 4787 2694 4833 2746
rect 4857 2694 4903 2746
rect 4903 2694 4913 2746
rect 4937 2694 4967 2746
rect 4967 2694 4993 2746
rect 4697 2692 4753 2694
rect 4777 2692 4833 2694
rect 4857 2692 4913 2694
rect 4937 2692 4993 2694
rect 5262 3168 5318 3224
rect 5262 2896 5318 2952
rect 5170 2352 5226 2408
rect 4618 992 4674 1048
rect 4894 1672 4950 1728
rect 5446 1536 5502 1592
rect 5630 2896 5686 2952
rect 5630 2488 5686 2544
rect 5814 6296 5870 6352
rect 5998 11056 6054 11112
rect 6568 11994 6624 11996
rect 6648 11994 6704 11996
rect 6728 11994 6784 11996
rect 6808 11994 6864 11996
rect 6568 11942 6594 11994
rect 6594 11942 6624 11994
rect 6648 11942 6658 11994
rect 6658 11942 6704 11994
rect 6728 11942 6774 11994
rect 6774 11942 6784 11994
rect 6808 11942 6838 11994
rect 6838 11942 6864 11994
rect 6568 11940 6624 11942
rect 6648 11940 6704 11942
rect 6728 11940 6784 11942
rect 6808 11940 6864 11942
rect 6550 11736 6606 11792
rect 6182 11056 6238 11112
rect 6458 11328 6514 11384
rect 6274 10104 6330 10160
rect 6182 9696 6238 9752
rect 6550 11056 6606 11112
rect 6568 10906 6624 10908
rect 6648 10906 6704 10908
rect 6728 10906 6784 10908
rect 6808 10906 6864 10908
rect 6568 10854 6594 10906
rect 6594 10854 6624 10906
rect 6648 10854 6658 10906
rect 6658 10854 6704 10906
rect 6728 10854 6774 10906
rect 6774 10854 6784 10906
rect 6808 10854 6838 10906
rect 6838 10854 6864 10906
rect 6568 10852 6624 10854
rect 6648 10852 6704 10854
rect 6728 10852 6784 10854
rect 6808 10852 6864 10854
rect 6550 10648 6606 10704
rect 6642 10376 6698 10432
rect 6734 10240 6790 10296
rect 6918 10104 6974 10160
rect 6568 9818 6624 9820
rect 6648 9818 6704 9820
rect 6728 9818 6784 9820
rect 6808 9818 6864 9820
rect 6568 9766 6594 9818
rect 6594 9766 6624 9818
rect 6648 9766 6658 9818
rect 6658 9766 6704 9818
rect 6728 9766 6774 9818
rect 6774 9766 6784 9818
rect 6808 9766 6838 9818
rect 6838 9766 6864 9818
rect 6568 9764 6624 9766
rect 6648 9764 6704 9766
rect 6728 9764 6784 9766
rect 6808 9764 6864 9766
rect 5814 4528 5870 4584
rect 5814 4392 5870 4448
rect 5906 4120 5962 4176
rect 5814 3576 5870 3632
rect 6182 6568 6238 6624
rect 6090 4528 6146 4584
rect 6090 4020 6092 4040
rect 6092 4020 6144 4040
rect 6144 4020 6146 4040
rect 6090 3984 6146 4020
rect 5906 856 5962 912
rect 6274 5092 6330 5128
rect 6274 5072 6276 5092
rect 6276 5072 6328 5092
rect 6328 5072 6330 5092
rect 6550 9152 6606 9208
rect 6458 8880 6514 8936
rect 6918 9036 6974 9072
rect 6918 9016 6920 9036
rect 6920 9016 6972 9036
rect 6972 9016 6974 9036
rect 6568 8730 6624 8732
rect 6648 8730 6704 8732
rect 6728 8730 6784 8732
rect 6808 8730 6864 8732
rect 6568 8678 6594 8730
rect 6594 8678 6624 8730
rect 6648 8678 6658 8730
rect 6658 8678 6704 8730
rect 6728 8678 6774 8730
rect 6774 8678 6784 8730
rect 6808 8678 6838 8730
rect 6838 8678 6864 8730
rect 6568 8676 6624 8678
rect 6648 8676 6704 8678
rect 6728 8676 6784 8678
rect 6808 8676 6864 8678
rect 6568 7642 6624 7644
rect 6648 7642 6704 7644
rect 6728 7642 6784 7644
rect 6808 7642 6864 7644
rect 6568 7590 6594 7642
rect 6594 7590 6624 7642
rect 6648 7590 6658 7642
rect 6658 7590 6704 7642
rect 6728 7590 6774 7642
rect 6774 7590 6784 7642
rect 6808 7590 6838 7642
rect 6838 7590 6864 7642
rect 6568 7588 6624 7590
rect 6648 7588 6704 7590
rect 6728 7588 6784 7590
rect 6808 7588 6864 7590
rect 6918 7268 6974 7304
rect 6918 7248 6920 7268
rect 6920 7248 6972 7268
rect 6972 7248 6974 7268
rect 6918 6704 6974 6760
rect 6568 6554 6624 6556
rect 6648 6554 6704 6556
rect 6728 6554 6784 6556
rect 6808 6554 6864 6556
rect 6568 6502 6594 6554
rect 6594 6502 6624 6554
rect 6648 6502 6658 6554
rect 6658 6502 6704 6554
rect 6728 6502 6774 6554
rect 6774 6502 6784 6554
rect 6808 6502 6838 6554
rect 6838 6502 6864 6554
rect 6568 6500 6624 6502
rect 6648 6500 6704 6502
rect 6728 6500 6784 6502
rect 6808 6500 6864 6502
rect 6274 3576 6330 3632
rect 6568 5466 6624 5468
rect 6648 5466 6704 5468
rect 6728 5466 6784 5468
rect 6808 5466 6864 5468
rect 6568 5414 6594 5466
rect 6594 5414 6624 5466
rect 6648 5414 6658 5466
rect 6658 5414 6704 5466
rect 6728 5414 6774 5466
rect 6774 5414 6784 5466
rect 6808 5414 6838 5466
rect 6838 5414 6864 5466
rect 6568 5412 6624 5414
rect 6648 5412 6704 5414
rect 6728 5412 6784 5414
rect 6808 5412 6864 5414
rect 6550 4528 6606 4584
rect 6918 4800 6974 4856
rect 6568 4378 6624 4380
rect 6648 4378 6704 4380
rect 6728 4378 6784 4380
rect 6808 4378 6864 4380
rect 6568 4326 6594 4378
rect 6594 4326 6624 4378
rect 6648 4326 6658 4378
rect 6658 4326 6704 4378
rect 6728 4326 6774 4378
rect 6774 4326 6784 4378
rect 6808 4326 6838 4378
rect 6838 4326 6864 4378
rect 6568 4324 6624 4326
rect 6648 4324 6704 4326
rect 6728 4324 6784 4326
rect 6808 4324 6864 4326
rect 7194 8472 7250 8528
rect 7378 11192 7434 11248
rect 7470 9424 7526 9480
rect 7194 5344 7250 5400
rect 6826 3848 6882 3904
rect 6458 3440 6514 3496
rect 7654 11056 7710 11112
rect 7562 9288 7618 9344
rect 10309 13082 10365 13084
rect 10389 13082 10445 13084
rect 10469 13082 10525 13084
rect 10549 13082 10605 13084
rect 10309 13030 10335 13082
rect 10335 13030 10365 13082
rect 10389 13030 10399 13082
rect 10399 13030 10445 13082
rect 10469 13030 10515 13082
rect 10515 13030 10525 13082
rect 10549 13030 10579 13082
rect 10579 13030 10605 13082
rect 10309 13028 10365 13030
rect 10389 13028 10445 13030
rect 10469 13028 10525 13030
rect 10549 13028 10605 13030
rect 10046 12824 10102 12880
rect 8438 12538 8494 12540
rect 8518 12538 8574 12540
rect 8598 12538 8654 12540
rect 8678 12538 8734 12540
rect 8438 12486 8464 12538
rect 8464 12486 8494 12538
rect 8518 12486 8528 12538
rect 8528 12486 8574 12538
rect 8598 12486 8644 12538
rect 8644 12486 8654 12538
rect 8678 12486 8708 12538
rect 8708 12486 8734 12538
rect 8438 12484 8494 12486
rect 8518 12484 8574 12486
rect 8598 12484 8654 12486
rect 8678 12484 8734 12486
rect 8114 11600 8170 11656
rect 8438 11450 8494 11452
rect 8518 11450 8574 11452
rect 8598 11450 8654 11452
rect 8678 11450 8734 11452
rect 8438 11398 8464 11450
rect 8464 11398 8494 11450
rect 8518 11398 8528 11450
rect 8528 11398 8574 11450
rect 8598 11398 8644 11450
rect 8644 11398 8654 11450
rect 8678 11398 8708 11450
rect 8708 11398 8734 11450
rect 8438 11396 8494 11398
rect 8518 11396 8574 11398
rect 8598 11396 8654 11398
rect 8678 11396 8734 11398
rect 7838 9152 7894 9208
rect 7562 5344 7618 5400
rect 7562 5208 7618 5264
rect 7378 4120 7434 4176
rect 6568 3290 6624 3292
rect 6648 3290 6704 3292
rect 6728 3290 6784 3292
rect 6808 3290 6864 3292
rect 6568 3238 6594 3290
rect 6594 3238 6624 3290
rect 6648 3238 6658 3290
rect 6658 3238 6704 3290
rect 6728 3238 6774 3290
rect 6774 3238 6784 3290
rect 6808 3238 6838 3290
rect 6838 3238 6864 3290
rect 6568 3236 6624 3238
rect 6648 3236 6704 3238
rect 6728 3236 6784 3238
rect 6808 3236 6864 3238
rect 6826 2896 6882 2952
rect 6568 2202 6624 2204
rect 6648 2202 6704 2204
rect 6728 2202 6784 2204
rect 6808 2202 6864 2204
rect 6568 2150 6594 2202
rect 6594 2150 6624 2202
rect 6648 2150 6658 2202
rect 6658 2150 6704 2202
rect 6728 2150 6774 2202
rect 6774 2150 6784 2202
rect 6808 2150 6838 2202
rect 6838 2150 6864 2202
rect 6568 2148 6624 2150
rect 6648 2148 6704 2150
rect 6728 2148 6784 2150
rect 6808 2148 6864 2150
rect 6734 1264 6790 1320
rect 7286 3576 7342 3632
rect 7470 3440 7526 3496
rect 7286 3168 7342 3224
rect 7194 2932 7196 2952
rect 7196 2932 7248 2952
rect 7248 2932 7250 2952
rect 7194 2896 7250 2932
rect 7194 1808 7250 1864
rect 7930 4528 7986 4584
rect 7930 2760 7986 2816
rect 8438 10362 8494 10364
rect 8518 10362 8574 10364
rect 8598 10362 8654 10364
rect 8678 10362 8734 10364
rect 8438 10310 8464 10362
rect 8464 10310 8494 10362
rect 8518 10310 8528 10362
rect 8528 10310 8574 10362
rect 8598 10310 8644 10362
rect 8644 10310 8654 10362
rect 8678 10310 8708 10362
rect 8708 10310 8734 10362
rect 8438 10308 8494 10310
rect 8518 10308 8574 10310
rect 8598 10308 8654 10310
rect 8678 10308 8734 10310
rect 8438 9274 8494 9276
rect 8518 9274 8574 9276
rect 8598 9274 8654 9276
rect 8678 9274 8734 9276
rect 8438 9222 8464 9274
rect 8464 9222 8494 9274
rect 8518 9222 8528 9274
rect 8528 9222 8574 9274
rect 8598 9222 8644 9274
rect 8644 9222 8654 9274
rect 8678 9222 8708 9274
rect 8708 9222 8734 9274
rect 8438 9220 8494 9222
rect 8518 9220 8574 9222
rect 8598 9220 8654 9222
rect 8678 9220 8734 9222
rect 8390 9016 8446 9072
rect 8438 8186 8494 8188
rect 8518 8186 8574 8188
rect 8598 8186 8654 8188
rect 8678 8186 8734 8188
rect 8438 8134 8464 8186
rect 8464 8134 8494 8186
rect 8518 8134 8528 8186
rect 8528 8134 8574 8186
rect 8598 8134 8644 8186
rect 8644 8134 8654 8186
rect 8678 8134 8708 8186
rect 8708 8134 8734 8186
rect 8438 8132 8494 8134
rect 8518 8132 8574 8134
rect 8598 8132 8654 8134
rect 8678 8132 8734 8134
rect 8298 7928 8354 7984
rect 8438 7098 8494 7100
rect 8518 7098 8574 7100
rect 8598 7098 8654 7100
rect 8678 7098 8734 7100
rect 8438 7046 8464 7098
rect 8464 7046 8494 7098
rect 8518 7046 8528 7098
rect 8528 7046 8574 7098
rect 8598 7046 8644 7098
rect 8644 7046 8654 7098
rect 8678 7046 8708 7098
rect 8708 7046 8734 7098
rect 8438 7044 8494 7046
rect 8518 7044 8574 7046
rect 8598 7044 8654 7046
rect 8678 7044 8734 7046
rect 8438 6010 8494 6012
rect 8518 6010 8574 6012
rect 8598 6010 8654 6012
rect 8678 6010 8734 6012
rect 8438 5958 8464 6010
rect 8464 5958 8494 6010
rect 8518 5958 8528 6010
rect 8528 5958 8574 6010
rect 8598 5958 8644 6010
rect 8644 5958 8654 6010
rect 8678 5958 8708 6010
rect 8708 5958 8734 6010
rect 8438 5956 8494 5958
rect 8518 5956 8574 5958
rect 8598 5956 8654 5958
rect 8678 5956 8734 5958
rect 8206 5108 8208 5128
rect 8208 5108 8260 5128
rect 8260 5108 8262 5128
rect 8206 5072 8262 5108
rect 8114 4528 8170 4584
rect 8114 4020 8116 4040
rect 8116 4020 8168 4040
rect 8168 4020 8170 4040
rect 8114 3984 8170 4020
rect 8114 3304 8170 3360
rect 8438 4922 8494 4924
rect 8518 4922 8574 4924
rect 8598 4922 8654 4924
rect 8678 4922 8734 4924
rect 8438 4870 8464 4922
rect 8464 4870 8494 4922
rect 8518 4870 8528 4922
rect 8528 4870 8574 4922
rect 8598 4870 8644 4922
rect 8644 4870 8654 4922
rect 8678 4870 8708 4922
rect 8708 4870 8734 4922
rect 8438 4868 8494 4870
rect 8518 4868 8574 4870
rect 8598 4868 8654 4870
rect 8678 4868 8734 4870
rect 8574 4256 8630 4312
rect 8666 4120 8722 4176
rect 8438 3834 8494 3836
rect 8518 3834 8574 3836
rect 8598 3834 8654 3836
rect 8678 3834 8734 3836
rect 8438 3782 8464 3834
rect 8464 3782 8494 3834
rect 8518 3782 8528 3834
rect 8528 3782 8574 3834
rect 8598 3782 8644 3834
rect 8644 3782 8654 3834
rect 8678 3782 8708 3834
rect 8708 3782 8734 3834
rect 8438 3780 8494 3782
rect 8518 3780 8574 3782
rect 8598 3780 8654 3782
rect 8678 3780 8734 3782
rect 9770 12144 9826 12200
rect 9954 11600 10010 11656
rect 9678 10684 9680 10704
rect 9680 10684 9732 10704
rect 9732 10684 9734 10704
rect 9678 10648 9734 10684
rect 9494 10376 9550 10432
rect 8942 5208 8998 5264
rect 8298 3440 8354 3496
rect 8666 3168 8722 3224
rect 8438 2746 8494 2748
rect 8518 2746 8574 2748
rect 8598 2746 8654 2748
rect 8678 2746 8734 2748
rect 8438 2694 8464 2746
rect 8464 2694 8494 2746
rect 8518 2694 8528 2746
rect 8528 2694 8574 2746
rect 8598 2694 8644 2746
rect 8644 2694 8654 2746
rect 8678 2694 8708 2746
rect 8708 2694 8734 2746
rect 8438 2692 8494 2694
rect 8518 2692 8574 2694
rect 8598 2692 8654 2694
rect 8678 2692 8734 2694
rect 8390 2524 8392 2544
rect 8392 2524 8444 2544
rect 8444 2524 8446 2544
rect 8390 2488 8446 2524
rect 8666 2352 8722 2408
rect 8942 3440 8998 3496
rect 8482 1536 8538 1592
rect 8850 2216 8906 2272
rect 8758 1944 8814 2000
rect 9310 4564 9312 4584
rect 9312 4564 9364 4584
rect 9364 4564 9366 4584
rect 9310 4528 9366 4564
rect 9310 4156 9312 4176
rect 9312 4156 9364 4176
rect 9364 4156 9366 4176
rect 9310 4120 9366 4156
rect 9310 3984 9366 4040
rect 10309 11994 10365 11996
rect 10389 11994 10445 11996
rect 10469 11994 10525 11996
rect 10549 11994 10605 11996
rect 10309 11942 10335 11994
rect 10335 11942 10365 11994
rect 10389 11942 10399 11994
rect 10399 11942 10445 11994
rect 10469 11942 10515 11994
rect 10515 11942 10525 11994
rect 10549 11942 10579 11994
rect 10579 11942 10605 11994
rect 10309 11940 10365 11942
rect 10389 11940 10445 11942
rect 10469 11940 10525 11942
rect 10549 11940 10605 11942
rect 10230 11600 10286 11656
rect 10414 11636 10416 11656
rect 10416 11636 10468 11656
rect 10468 11636 10470 11656
rect 10414 11600 10470 11636
rect 10309 10906 10365 10908
rect 10389 10906 10445 10908
rect 10469 10906 10525 10908
rect 10549 10906 10605 10908
rect 10309 10854 10335 10906
rect 10335 10854 10365 10906
rect 10389 10854 10399 10906
rect 10399 10854 10445 10906
rect 10469 10854 10515 10906
rect 10515 10854 10525 10906
rect 10549 10854 10579 10906
rect 10579 10854 10605 10906
rect 10309 10852 10365 10854
rect 10389 10852 10445 10854
rect 10469 10852 10525 10854
rect 10549 10852 10605 10854
rect 10230 10648 10286 10704
rect 9954 9968 10010 10024
rect 9494 6840 9550 6896
rect 9494 4684 9550 4720
rect 9494 4664 9496 4684
rect 9496 4664 9548 4684
rect 9548 4664 9550 4684
rect 9586 4392 9642 4448
rect 9586 4120 9642 4176
rect 9678 3712 9734 3768
rect 10506 10412 10508 10432
rect 10508 10412 10560 10432
rect 10560 10412 10562 10432
rect 10506 10376 10562 10412
rect 10309 9818 10365 9820
rect 10389 9818 10445 9820
rect 10469 9818 10525 9820
rect 10549 9818 10605 9820
rect 10309 9766 10335 9818
rect 10335 9766 10365 9818
rect 10389 9766 10399 9818
rect 10399 9766 10445 9818
rect 10469 9766 10515 9818
rect 10515 9766 10525 9818
rect 10549 9766 10579 9818
rect 10579 9766 10605 9818
rect 10309 9764 10365 9766
rect 10389 9764 10445 9766
rect 10469 9764 10525 9766
rect 10549 9764 10605 9766
rect 9954 8084 10010 8120
rect 9954 8064 9956 8084
rect 9956 8064 10008 8084
rect 10008 8064 10010 8084
rect 9862 5092 9918 5128
rect 9862 5072 9864 5092
rect 9864 5072 9916 5092
rect 9916 5072 9918 5092
rect 10309 8730 10365 8732
rect 10389 8730 10445 8732
rect 10469 8730 10525 8732
rect 10549 8730 10605 8732
rect 10309 8678 10335 8730
rect 10335 8678 10365 8730
rect 10389 8678 10399 8730
rect 10399 8678 10445 8730
rect 10469 8678 10515 8730
rect 10515 8678 10525 8730
rect 10549 8678 10579 8730
rect 10579 8678 10605 8730
rect 10309 8676 10365 8678
rect 10389 8676 10445 8678
rect 10469 8676 10525 8678
rect 10549 8676 10605 8678
rect 11242 12144 11298 12200
rect 11242 11600 11298 11656
rect 10782 8064 10838 8120
rect 10598 7928 10654 7984
rect 10309 7642 10365 7644
rect 10389 7642 10445 7644
rect 10469 7642 10525 7644
rect 10549 7642 10605 7644
rect 10309 7590 10335 7642
rect 10335 7590 10365 7642
rect 10389 7590 10399 7642
rect 10399 7590 10445 7642
rect 10469 7590 10515 7642
rect 10515 7590 10525 7642
rect 10549 7590 10579 7642
rect 10579 7590 10605 7642
rect 10309 7588 10365 7590
rect 10389 7588 10445 7590
rect 10469 7588 10525 7590
rect 10549 7588 10605 7590
rect 10309 6554 10365 6556
rect 10389 6554 10445 6556
rect 10469 6554 10525 6556
rect 10549 6554 10605 6556
rect 10309 6502 10335 6554
rect 10335 6502 10365 6554
rect 10389 6502 10399 6554
rect 10399 6502 10445 6554
rect 10469 6502 10515 6554
rect 10515 6502 10525 6554
rect 10549 6502 10579 6554
rect 10579 6502 10605 6554
rect 10309 6500 10365 6502
rect 10389 6500 10445 6502
rect 10469 6500 10525 6502
rect 10549 6500 10605 6502
rect 10309 5466 10365 5468
rect 10389 5466 10445 5468
rect 10469 5466 10525 5468
rect 10549 5466 10605 5468
rect 10309 5414 10335 5466
rect 10335 5414 10365 5466
rect 10389 5414 10399 5466
rect 10399 5414 10445 5466
rect 10469 5414 10515 5466
rect 10515 5414 10525 5466
rect 10549 5414 10579 5466
rect 10579 5414 10605 5466
rect 10309 5412 10365 5414
rect 10389 5412 10445 5414
rect 10469 5412 10525 5414
rect 10549 5412 10605 5414
rect 9862 2932 9864 2952
rect 9864 2932 9916 2952
rect 9916 2932 9918 2952
rect 9862 2896 9918 2932
rect 10598 4936 10654 4992
rect 10046 1128 10102 1184
rect 10309 4378 10365 4380
rect 10389 4378 10445 4380
rect 10469 4378 10525 4380
rect 10549 4378 10605 4380
rect 10309 4326 10335 4378
rect 10335 4326 10365 4378
rect 10389 4326 10399 4378
rect 10399 4326 10445 4378
rect 10469 4326 10515 4378
rect 10515 4326 10525 4378
rect 10549 4326 10579 4378
rect 10579 4326 10605 4378
rect 10309 4324 10365 4326
rect 10389 4324 10445 4326
rect 10469 4324 10525 4326
rect 10549 4324 10605 4326
rect 10322 3984 10378 4040
rect 10309 3290 10365 3292
rect 10389 3290 10445 3292
rect 10469 3290 10525 3292
rect 10549 3290 10605 3292
rect 10309 3238 10335 3290
rect 10335 3238 10365 3290
rect 10389 3238 10399 3290
rect 10399 3238 10445 3290
rect 10469 3238 10515 3290
rect 10515 3238 10525 3290
rect 10549 3238 10579 3290
rect 10579 3238 10605 3290
rect 10309 3236 10365 3238
rect 10389 3236 10445 3238
rect 10469 3236 10525 3238
rect 10549 3236 10605 3238
rect 10966 5072 11022 5128
rect 10874 4120 10930 4176
rect 10966 3032 11022 3088
rect 10309 2202 10365 2204
rect 10389 2202 10445 2204
rect 10469 2202 10525 2204
rect 10549 2202 10605 2204
rect 10309 2150 10335 2202
rect 10335 2150 10365 2202
rect 10389 2150 10399 2202
rect 10399 2150 10445 2202
rect 10469 2150 10515 2202
rect 10515 2150 10525 2202
rect 10549 2150 10579 2202
rect 10579 2150 10605 2202
rect 10309 2148 10365 2150
rect 10389 2148 10445 2150
rect 10469 2148 10525 2150
rect 10549 2148 10605 2150
rect 11334 3168 11390 3224
rect 11242 2760 11298 2816
rect 12070 4120 12126 4176
rect 11610 3168 11666 3224
rect 11794 3596 11850 3632
rect 11794 3576 11796 3596
rect 11796 3576 11848 3596
rect 11848 3576 11850 3596
rect 11794 2760 11850 2816
<< metal3 >>
rect 2814 13088 3134 13089
rect 2814 13024 2822 13088
rect 2886 13024 2902 13088
rect 2966 13024 2982 13088
rect 3046 13024 3062 13088
rect 3126 13024 3134 13088
rect 2814 13023 3134 13024
rect 6556 13088 6876 13089
rect 6556 13024 6564 13088
rect 6628 13024 6644 13088
rect 6708 13024 6724 13088
rect 6788 13024 6804 13088
rect 6868 13024 6876 13088
rect 6556 13023 6876 13024
rect 10297 13088 10617 13089
rect 10297 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10465 13088
rect 10529 13024 10545 13088
rect 10609 13024 10617 13088
rect 10297 13023 10617 13024
rect 1158 12820 1164 12884
rect 1228 12882 1234 12884
rect 10041 12882 10107 12885
rect 1228 12880 10107 12882
rect 1228 12824 10046 12880
rect 10102 12824 10107 12880
rect 1228 12822 10107 12824
rect 1228 12820 1234 12822
rect 10041 12819 10107 12822
rect 4685 12544 5005 12545
rect 4685 12480 4693 12544
rect 4757 12480 4773 12544
rect 4837 12480 4853 12544
rect 4917 12480 4933 12544
rect 4997 12480 5005 12544
rect 4685 12479 5005 12480
rect 8426 12544 8746 12545
rect 8426 12480 8434 12544
rect 8498 12480 8514 12544
rect 8578 12480 8594 12544
rect 8658 12480 8674 12544
rect 8738 12480 8746 12544
rect 8426 12479 8746 12480
rect 9765 12202 9831 12205
rect 11237 12202 11303 12205
rect 9765 12200 11303 12202
rect 9765 12144 9770 12200
rect 9826 12144 11242 12200
rect 11298 12144 11303 12200
rect 9765 12142 11303 12144
rect 9765 12139 9831 12142
rect 11237 12139 11303 12142
rect 2814 12000 3134 12001
rect 2814 11936 2822 12000
rect 2886 11936 2902 12000
rect 2966 11936 2982 12000
rect 3046 11936 3062 12000
rect 3126 11936 3134 12000
rect 2814 11935 3134 11936
rect 6556 12000 6876 12001
rect 6556 11936 6564 12000
rect 6628 11936 6644 12000
rect 6708 11936 6724 12000
rect 6788 11936 6804 12000
rect 6868 11936 6876 12000
rect 6556 11935 6876 11936
rect 10297 12000 10617 12001
rect 10297 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10545 12000
rect 10609 11936 10617 12000
rect 10297 11935 10617 11936
rect 5073 11794 5139 11797
rect 6545 11794 6611 11797
rect 5073 11792 6611 11794
rect 5073 11736 5078 11792
rect 5134 11736 6550 11792
rect 6606 11736 6611 11792
rect 5073 11734 6611 11736
rect 5073 11731 5139 11734
rect 6545 11731 6611 11734
rect 3049 11658 3115 11661
rect 8109 11658 8175 11661
rect 3049 11656 8175 11658
rect 3049 11600 3054 11656
rect 3110 11600 8114 11656
rect 8170 11600 8175 11656
rect 3049 11598 8175 11600
rect 3049 11595 3115 11598
rect 8109 11595 8175 11598
rect 9949 11658 10015 11661
rect 10225 11658 10291 11661
rect 9949 11656 10291 11658
rect 9949 11600 9954 11656
rect 10010 11600 10230 11656
rect 10286 11600 10291 11656
rect 9949 11598 10291 11600
rect 9949 11595 10015 11598
rect 10225 11595 10291 11598
rect 10409 11658 10475 11661
rect 11237 11658 11303 11661
rect 10409 11656 11303 11658
rect 10409 11600 10414 11656
rect 10470 11600 11242 11656
rect 11298 11600 11303 11656
rect 10409 11598 11303 11600
rect 10409 11595 10475 11598
rect 11237 11595 11303 11598
rect 4685 11456 5005 11457
rect 4685 11392 4693 11456
rect 4757 11392 4773 11456
rect 4837 11392 4853 11456
rect 4917 11392 4933 11456
rect 4997 11392 5005 11456
rect 4685 11391 5005 11392
rect 8426 11456 8746 11457
rect 8426 11392 8434 11456
rect 8498 11392 8514 11456
rect 8578 11392 8594 11456
rect 8658 11392 8674 11456
rect 8738 11392 8746 11456
rect 8426 11391 8746 11392
rect 5625 11386 5691 11389
rect 6453 11386 6519 11389
rect 5625 11384 6519 11386
rect 5625 11328 5630 11384
rect 5686 11328 6458 11384
rect 6514 11328 6519 11384
rect 5625 11326 6519 11328
rect 5625 11323 5691 11326
rect 6453 11323 6519 11326
rect 5625 11250 5691 11253
rect 7230 11250 7236 11252
rect 5625 11248 7236 11250
rect 5625 11192 5630 11248
rect 5686 11192 7236 11248
rect 5625 11190 7236 11192
rect 5625 11187 5691 11190
rect 7230 11188 7236 11190
rect 7300 11188 7306 11252
rect 7373 11250 7439 11253
rect 7598 11250 7604 11252
rect 7373 11248 7604 11250
rect 7373 11192 7378 11248
rect 7434 11192 7604 11248
rect 7373 11190 7604 11192
rect 7373 11187 7439 11190
rect 7598 11188 7604 11190
rect 7668 11188 7674 11252
rect 5717 11116 5783 11117
rect 5717 11112 5764 11116
rect 5828 11114 5834 11116
rect 5993 11114 6059 11117
rect 5717 11056 5722 11112
rect 5717 11052 5764 11056
rect 5828 11054 5874 11114
rect 5950 11112 6059 11114
rect 5950 11056 5998 11112
rect 6054 11056 6059 11112
rect 5828 11052 5834 11054
rect 5717 11051 5783 11052
rect 5950 11051 6059 11056
rect 6177 11114 6243 11117
rect 6545 11114 6611 11117
rect 6177 11112 6611 11114
rect 6177 11056 6182 11112
rect 6238 11056 6550 11112
rect 6606 11056 6611 11112
rect 6177 11054 6611 11056
rect 6177 11051 6243 11054
rect 6545 11051 6611 11054
rect 7649 11114 7715 11117
rect 7782 11114 7788 11116
rect 7649 11112 7788 11114
rect 7649 11056 7654 11112
rect 7710 11056 7788 11112
rect 7649 11054 7788 11056
rect 7649 11051 7715 11054
rect 7782 11052 7788 11054
rect 7852 11052 7858 11116
rect 5625 10978 5691 10981
rect 5950 10978 6010 11051
rect 5625 10976 6010 10978
rect 5625 10920 5630 10976
rect 5686 10920 6010 10976
rect 5625 10918 6010 10920
rect 5625 10915 5691 10918
rect 2814 10912 3134 10913
rect 2814 10848 2822 10912
rect 2886 10848 2902 10912
rect 2966 10848 2982 10912
rect 3046 10848 3062 10912
rect 3126 10848 3134 10912
rect 2814 10847 3134 10848
rect 6556 10912 6876 10913
rect 6556 10848 6564 10912
rect 6628 10848 6644 10912
rect 6708 10848 6724 10912
rect 6788 10848 6804 10912
rect 6868 10848 6876 10912
rect 6556 10847 6876 10848
rect 10297 10912 10617 10913
rect 10297 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10545 10912
rect 10609 10848 10617 10912
rect 10297 10847 10617 10848
rect 4102 10780 4108 10844
rect 4172 10842 4178 10844
rect 4613 10842 4679 10845
rect 4172 10840 4679 10842
rect 4172 10784 4618 10840
rect 4674 10784 4679 10840
rect 4172 10782 4679 10784
rect 4172 10780 4178 10782
rect 4613 10779 4679 10782
rect 2773 10706 2839 10709
rect 4470 10706 4476 10708
rect 2773 10704 4476 10706
rect 2773 10648 2778 10704
rect 2834 10648 4476 10704
rect 2773 10646 4476 10648
rect 2773 10643 2839 10646
rect 4470 10644 4476 10646
rect 4540 10644 4546 10708
rect 4797 10706 4863 10709
rect 6545 10706 6611 10709
rect 4797 10704 6611 10706
rect 4797 10648 4802 10704
rect 4858 10648 6550 10704
rect 6606 10648 6611 10704
rect 4797 10646 6611 10648
rect 4797 10643 4863 10646
rect 6545 10643 6611 10646
rect 9673 10706 9739 10709
rect 10225 10706 10291 10709
rect 9673 10704 10291 10706
rect 9673 10648 9678 10704
rect 9734 10648 10230 10704
rect 10286 10648 10291 10704
rect 9673 10646 10291 10648
rect 9673 10643 9739 10646
rect 10225 10643 10291 10646
rect 4286 10508 4292 10572
rect 4356 10570 4362 10572
rect 4705 10570 4771 10573
rect 4356 10568 4771 10570
rect 4356 10512 4710 10568
rect 4766 10512 4771 10568
rect 4356 10510 4771 10512
rect 4356 10508 4362 10510
rect 4705 10507 4771 10510
rect 4889 10570 4955 10573
rect 8150 10570 8156 10572
rect 4889 10568 8156 10570
rect 4889 10512 4894 10568
rect 4950 10512 8156 10568
rect 4889 10510 8156 10512
rect 4889 10507 4955 10510
rect 8150 10508 8156 10510
rect 8220 10508 8226 10572
rect 2773 10434 2839 10437
rect 3693 10434 3759 10437
rect 2773 10432 3759 10434
rect 2773 10376 2778 10432
rect 2834 10376 3698 10432
rect 3754 10376 3759 10432
rect 2773 10374 3759 10376
rect 2773 10371 2839 10374
rect 3693 10371 3759 10374
rect 5441 10434 5507 10437
rect 6637 10434 6703 10437
rect 5441 10432 6703 10434
rect 5441 10376 5446 10432
rect 5502 10376 6642 10432
rect 6698 10376 6703 10432
rect 5441 10374 6703 10376
rect 5441 10371 5507 10374
rect 6637 10371 6703 10374
rect 9489 10434 9555 10437
rect 10501 10434 10567 10437
rect 9489 10432 10567 10434
rect 9489 10376 9494 10432
rect 9550 10376 10506 10432
rect 10562 10376 10567 10432
rect 9489 10374 10567 10376
rect 9489 10371 9555 10374
rect 10501 10371 10567 10374
rect 4685 10368 5005 10369
rect 4685 10304 4693 10368
rect 4757 10304 4773 10368
rect 4837 10304 4853 10368
rect 4917 10304 4933 10368
rect 4997 10304 5005 10368
rect 4685 10303 5005 10304
rect 8426 10368 8746 10369
rect 8426 10304 8434 10368
rect 8498 10304 8514 10368
rect 8578 10304 8594 10368
rect 8658 10304 8674 10368
rect 8738 10304 8746 10368
rect 8426 10303 8746 10304
rect 1761 10298 1827 10301
rect 3233 10298 3299 10301
rect 1761 10296 3299 10298
rect 1761 10240 1766 10296
rect 1822 10240 3238 10296
rect 3294 10240 3299 10296
rect 1761 10238 3299 10240
rect 1761 10235 1827 10238
rect 3233 10235 3299 10238
rect 4429 10296 4495 10301
rect 4429 10240 4434 10296
rect 4490 10240 4495 10296
rect 4429 10235 4495 10240
rect 5165 10298 5231 10301
rect 6729 10298 6795 10301
rect 5165 10296 6795 10298
rect 5165 10240 5170 10296
rect 5226 10240 6734 10296
rect 6790 10240 6795 10296
rect 5165 10238 6795 10240
rect 5165 10235 5231 10238
rect 6729 10235 6795 10238
rect 473 10162 539 10165
rect 3417 10162 3483 10165
rect 3601 10162 3667 10165
rect 473 10160 2790 10162
rect 473 10104 478 10160
rect 534 10104 2790 10160
rect 473 10102 2790 10104
rect 473 10099 539 10102
rect 2730 10026 2790 10102
rect 3417 10160 3667 10162
rect 3417 10104 3422 10160
rect 3478 10104 3606 10160
rect 3662 10104 3667 10160
rect 3417 10102 3667 10104
rect 4432 10162 4492 10235
rect 6269 10162 6335 10165
rect 4432 10160 6335 10162
rect 4432 10104 6274 10160
rect 6330 10104 6335 10160
rect 4432 10102 6335 10104
rect 3417 10099 3483 10102
rect 3601 10099 3667 10102
rect 6269 10099 6335 10102
rect 6913 10162 6979 10165
rect 7046 10162 7052 10164
rect 6913 10160 7052 10162
rect 6913 10104 6918 10160
rect 6974 10104 7052 10160
rect 6913 10102 7052 10104
rect 6913 10099 6979 10102
rect 7046 10100 7052 10102
rect 7116 10100 7122 10164
rect 9949 10026 10015 10029
rect 2730 10024 10015 10026
rect 2730 9968 9954 10024
rect 10010 9968 10015 10024
rect 2730 9966 10015 9968
rect 9949 9963 10015 9966
rect 3325 9890 3391 9893
rect 3550 9890 3556 9892
rect 3325 9888 3556 9890
rect 3325 9832 3330 9888
rect 3386 9832 3556 9888
rect 3325 9830 3556 9832
rect 3325 9827 3391 9830
rect 3550 9828 3556 9830
rect 3620 9828 3626 9892
rect 4705 9890 4771 9893
rect 4981 9890 5047 9893
rect 4705 9888 5047 9890
rect 4705 9832 4710 9888
rect 4766 9832 4986 9888
rect 5042 9832 5047 9888
rect 4705 9830 5047 9832
rect 4705 9827 4771 9830
rect 4981 9827 5047 9830
rect 2814 9824 3134 9825
rect 2814 9760 2822 9824
rect 2886 9760 2902 9824
rect 2966 9760 2982 9824
rect 3046 9760 3062 9824
rect 3126 9760 3134 9824
rect 2814 9759 3134 9760
rect 6556 9824 6876 9825
rect 6556 9760 6564 9824
rect 6628 9760 6644 9824
rect 6708 9760 6724 9824
rect 6788 9760 6804 9824
rect 6868 9760 6876 9824
rect 6556 9759 6876 9760
rect 10297 9824 10617 9825
rect 10297 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10545 9824
rect 10609 9760 10617 9824
rect 10297 9759 10617 9760
rect 2313 9754 2379 9757
rect 6177 9754 6243 9757
rect 2313 9752 2698 9754
rect 2313 9696 2318 9752
rect 2374 9696 2698 9752
rect 2313 9694 2698 9696
rect 2313 9691 2379 9694
rect 2638 9690 2698 9694
rect 3328 9752 6243 9754
rect 3328 9696 6182 9752
rect 6238 9696 6243 9752
rect 3328 9694 6243 9696
rect 3328 9690 3388 9694
rect 6177 9691 6243 9694
rect 2638 9630 3388 9690
rect 5073 9616 5139 9621
rect 5073 9560 5078 9616
rect 5134 9560 5139 9616
rect 5073 9555 5139 9560
rect 5533 9618 5599 9621
rect 8886 9618 8892 9620
rect 5533 9616 8892 9618
rect 5533 9560 5538 9616
rect 5594 9560 8892 9616
rect 5533 9558 8892 9560
rect 5533 9555 5599 9558
rect 8886 9556 8892 9558
rect 8956 9556 8962 9620
rect 3366 9420 3372 9484
rect 3436 9482 3442 9484
rect 4889 9482 4955 9485
rect 3436 9480 4955 9482
rect 3436 9424 4894 9480
rect 4950 9424 4955 9480
rect 3436 9422 4955 9424
rect 5076 9482 5136 9555
rect 7465 9482 7531 9485
rect 5076 9480 7531 9482
rect 5076 9424 7470 9480
rect 7526 9424 7531 9480
rect 5076 9422 7531 9424
rect 3436 9420 3442 9422
rect 4889 9419 4955 9422
rect 7465 9419 7531 9422
rect 5349 9346 5415 9349
rect 7557 9346 7623 9349
rect 5349 9344 7623 9346
rect 5349 9288 5354 9344
rect 5410 9288 7562 9344
rect 7618 9288 7623 9344
rect 5349 9286 7623 9288
rect 5349 9283 5415 9286
rect 7557 9283 7623 9286
rect 4685 9280 5005 9281
rect 4685 9216 4693 9280
rect 4757 9216 4773 9280
rect 4837 9216 4853 9280
rect 4917 9216 4933 9280
rect 4997 9216 5005 9280
rect 4685 9215 5005 9216
rect 8426 9280 8746 9281
rect 8426 9216 8434 9280
rect 8498 9216 8514 9280
rect 8578 9216 8594 9280
rect 8658 9216 8674 9280
rect 8738 9216 8746 9280
rect 8426 9215 8746 9216
rect 1526 9148 1532 9212
rect 1596 9210 1602 9212
rect 3233 9210 3299 9213
rect 1596 9208 3299 9210
rect 1596 9152 3238 9208
rect 3294 9152 3299 9208
rect 1596 9150 3299 9152
rect 1596 9148 1602 9150
rect 3233 9147 3299 9150
rect 3969 9210 4035 9213
rect 5073 9210 5139 9213
rect 5390 9210 5396 9212
rect 3969 9208 4584 9210
rect 3969 9152 3974 9208
rect 4030 9152 4584 9208
rect 3969 9150 4584 9152
rect 3969 9147 4035 9150
rect 4524 9074 4584 9150
rect 5073 9208 5396 9210
rect 5073 9152 5078 9208
rect 5134 9152 5396 9208
rect 5073 9150 5396 9152
rect 5073 9147 5139 9150
rect 5390 9148 5396 9150
rect 5460 9148 5466 9212
rect 5533 9210 5599 9213
rect 6545 9210 6611 9213
rect 7833 9210 7899 9213
rect 5533 9208 7899 9210
rect 5533 9152 5538 9208
rect 5594 9152 6550 9208
rect 6606 9152 7838 9208
rect 7894 9152 7899 9208
rect 5533 9150 7899 9152
rect 5533 9147 5599 9150
rect 6545 9147 6611 9150
rect 7833 9147 7899 9150
rect 4797 9074 4863 9077
rect 4524 9072 4863 9074
rect 4524 9016 4802 9072
rect 4858 9016 4863 9072
rect 4524 9014 4863 9016
rect 4797 9011 4863 9014
rect 4981 9074 5047 9077
rect 6913 9074 6979 9077
rect 8385 9074 8451 9077
rect 4981 9072 8451 9074
rect 4981 9016 4986 9072
rect 5042 9016 6918 9072
rect 6974 9016 8390 9072
rect 8446 9016 8451 9072
rect 4981 9014 8451 9016
rect 4981 9011 5047 9014
rect 6913 9011 6979 9014
rect 8385 9011 8451 9014
rect 1393 8938 1459 8941
rect 4705 8938 4771 8941
rect 1393 8936 4771 8938
rect 1393 8880 1398 8936
rect 1454 8880 4710 8936
rect 4766 8880 4771 8936
rect 1393 8878 4771 8880
rect 1393 8875 1459 8878
rect 4705 8875 4771 8878
rect 6453 8938 6519 8941
rect 7966 8938 7972 8940
rect 6453 8936 7972 8938
rect 6453 8880 6458 8936
rect 6514 8880 7972 8936
rect 6453 8878 7972 8880
rect 6453 8875 6519 8878
rect 7966 8876 7972 8878
rect 8036 8876 8042 8940
rect 2814 8736 3134 8737
rect 2814 8672 2822 8736
rect 2886 8672 2902 8736
rect 2966 8672 2982 8736
rect 3046 8672 3062 8736
rect 3126 8672 3134 8736
rect 2814 8671 3134 8672
rect 6556 8736 6876 8737
rect 6556 8672 6564 8736
rect 6628 8672 6644 8736
rect 6708 8672 6724 8736
rect 6788 8672 6804 8736
rect 6868 8672 6876 8736
rect 6556 8671 6876 8672
rect 10297 8736 10617 8737
rect 10297 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10545 8736
rect 10609 8672 10617 8736
rect 10297 8671 10617 8672
rect 2221 8532 2287 8533
rect 2221 8528 2268 8532
rect 2332 8530 2338 8532
rect 3877 8530 3943 8533
rect 7189 8530 7255 8533
rect 2221 8472 2226 8528
rect 2221 8468 2268 8472
rect 2332 8470 2378 8530
rect 3877 8528 7255 8530
rect 3877 8472 3882 8528
rect 3938 8472 7194 8528
rect 7250 8472 7255 8528
rect 3877 8470 7255 8472
rect 2332 8468 2338 8470
rect 2221 8467 2287 8468
rect 3877 8467 3943 8470
rect 7189 8467 7255 8470
rect 5625 8396 5691 8397
rect 5574 8394 5580 8396
rect 5534 8334 5580 8394
rect 5644 8392 5691 8396
rect 5686 8336 5691 8392
rect 5574 8332 5580 8334
rect 5644 8332 5691 8336
rect 5625 8331 5691 8332
rect 4685 8192 5005 8193
rect 4685 8128 4693 8192
rect 4757 8128 4773 8192
rect 4837 8128 4853 8192
rect 4917 8128 4933 8192
rect 4997 8128 5005 8192
rect 4685 8127 5005 8128
rect 8426 8192 8746 8193
rect 8426 8128 8434 8192
rect 8498 8128 8514 8192
rect 8578 8128 8594 8192
rect 8658 8128 8674 8192
rect 8738 8128 8746 8192
rect 8426 8127 8746 8128
rect 3877 8124 3943 8125
rect 9949 8124 10015 8125
rect 10777 8124 10843 8125
rect 3877 8120 3924 8124
rect 3988 8122 3994 8124
rect 3877 8064 3882 8120
rect 3877 8060 3924 8064
rect 3988 8062 4034 8122
rect 9949 8120 9996 8124
rect 10060 8122 10066 8124
rect 10726 8122 10732 8124
rect 9949 8064 9954 8120
rect 3988 8060 3994 8062
rect 9949 8060 9996 8064
rect 10060 8062 10106 8122
rect 10686 8062 10732 8122
rect 10796 8120 10843 8124
rect 10838 8064 10843 8120
rect 10060 8060 10066 8062
rect 10726 8060 10732 8062
rect 10796 8060 10843 8064
rect 3877 8059 3943 8060
rect 9949 8059 10015 8060
rect 10777 8059 10843 8060
rect 3734 7924 3740 7988
rect 3804 7986 3810 7988
rect 8293 7986 8359 7989
rect 3804 7984 8359 7986
rect 3804 7928 8298 7984
rect 8354 7928 8359 7984
rect 3804 7926 8359 7928
rect 3804 7924 3810 7926
rect 8293 7923 8359 7926
rect 9622 7924 9628 7988
rect 9692 7986 9698 7988
rect 10593 7986 10659 7989
rect 9692 7984 10659 7986
rect 9692 7928 10598 7984
rect 10654 7928 10659 7984
rect 9692 7926 10659 7928
rect 9692 7924 9698 7926
rect 10593 7923 10659 7926
rect 565 7850 631 7853
rect 565 7848 4722 7850
rect 565 7792 570 7848
rect 626 7792 4722 7848
rect 565 7790 4722 7792
rect 565 7787 631 7790
rect 2814 7648 3134 7649
rect 2814 7584 2822 7648
rect 2886 7584 2902 7648
rect 2966 7584 2982 7648
rect 3046 7584 3062 7648
rect 3126 7584 3134 7648
rect 2814 7583 3134 7584
rect 4662 7306 4722 7790
rect 6556 7648 6876 7649
rect 6556 7584 6564 7648
rect 6628 7584 6644 7648
rect 6708 7584 6724 7648
rect 6788 7584 6804 7648
rect 6868 7584 6876 7648
rect 6556 7583 6876 7584
rect 10297 7648 10617 7649
rect 10297 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10465 7648
rect 10529 7584 10545 7648
rect 10609 7584 10617 7648
rect 10297 7583 10617 7584
rect 5073 7578 5139 7581
rect 5942 7578 5948 7580
rect 5073 7576 5948 7578
rect 5073 7520 5078 7576
rect 5134 7520 5948 7576
rect 5073 7518 5948 7520
rect 5073 7515 5139 7518
rect 5942 7516 5948 7518
rect 6012 7516 6018 7580
rect 6913 7306 6979 7309
rect 4662 7304 6979 7306
rect 4662 7248 6918 7304
rect 6974 7248 6979 7304
rect 4662 7246 6979 7248
rect 6913 7243 6979 7246
rect 4685 7104 5005 7105
rect 4685 7040 4693 7104
rect 4757 7040 4773 7104
rect 4837 7040 4853 7104
rect 4917 7040 4933 7104
rect 4997 7040 5005 7104
rect 4685 7039 5005 7040
rect 8426 7104 8746 7105
rect 8426 7040 8434 7104
rect 8498 7040 8514 7104
rect 8578 7040 8594 7104
rect 8658 7040 8674 7104
rect 8738 7040 8746 7104
rect 8426 7039 8746 7040
rect 2446 6836 2452 6900
rect 2516 6898 2522 6900
rect 3601 6898 3667 6901
rect 2516 6896 3667 6898
rect 2516 6840 3606 6896
rect 3662 6840 3667 6896
rect 2516 6838 3667 6840
rect 2516 6836 2522 6838
rect 3601 6835 3667 6838
rect 5257 6898 5323 6901
rect 9489 6898 9555 6901
rect 5257 6896 9555 6898
rect 5257 6840 5262 6896
rect 5318 6840 9494 6896
rect 9550 6840 9555 6896
rect 5257 6838 9555 6840
rect 5257 6835 5323 6838
rect 9489 6835 9555 6838
rect 2630 6700 2636 6764
rect 2700 6762 2706 6764
rect 2773 6762 2839 6765
rect 2700 6760 2839 6762
rect 2700 6704 2778 6760
rect 2834 6704 2839 6760
rect 2700 6702 2839 6704
rect 2700 6700 2706 6702
rect 2773 6699 2839 6702
rect 3049 6762 3115 6765
rect 4613 6762 4679 6765
rect 3049 6760 4679 6762
rect 3049 6704 3054 6760
rect 3110 6704 4618 6760
rect 4674 6704 4679 6760
rect 3049 6702 4679 6704
rect 3049 6699 3115 6702
rect 4613 6699 4679 6702
rect 6913 6762 6979 6765
rect 7414 6762 7420 6764
rect 6913 6760 7420 6762
rect 6913 6704 6918 6760
rect 6974 6704 7420 6760
rect 6913 6702 7420 6704
rect 6913 6699 6979 6702
rect 7414 6700 7420 6702
rect 7484 6700 7490 6764
rect 3233 6626 3299 6629
rect 5206 6626 5212 6628
rect 3233 6624 5212 6626
rect 3233 6568 3238 6624
rect 3294 6568 5212 6624
rect 3233 6566 5212 6568
rect 3233 6563 3299 6566
rect 5206 6564 5212 6566
rect 5276 6564 5282 6628
rect 5441 6626 5507 6629
rect 6177 6626 6243 6629
rect 5441 6624 6243 6626
rect 5441 6568 5446 6624
rect 5502 6568 6182 6624
rect 6238 6568 6243 6624
rect 5441 6566 6243 6568
rect 5441 6563 5507 6566
rect 6177 6563 6243 6566
rect 2814 6560 3134 6561
rect 2814 6496 2822 6560
rect 2886 6496 2902 6560
rect 2966 6496 2982 6560
rect 3046 6496 3062 6560
rect 3126 6496 3134 6560
rect 2814 6495 3134 6496
rect 6556 6560 6876 6561
rect 6556 6496 6564 6560
rect 6628 6496 6644 6560
rect 6708 6496 6724 6560
rect 6788 6496 6804 6560
rect 6868 6496 6876 6560
rect 6556 6495 6876 6496
rect 10297 6560 10617 6561
rect 10297 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10465 6560
rect 10529 6496 10545 6560
rect 10609 6496 10617 6560
rect 10297 6495 10617 6496
rect 5574 6428 5580 6492
rect 5644 6490 5650 6492
rect 5644 6430 5872 6490
rect 5644 6428 5650 6430
rect 5812 6357 5872 6430
rect 2405 6354 2471 6357
rect 5574 6354 5580 6356
rect 2405 6352 5580 6354
rect 2405 6296 2410 6352
rect 2466 6296 5580 6352
rect 2405 6294 5580 6296
rect 2405 6291 2471 6294
rect 5574 6292 5580 6294
rect 5644 6292 5650 6356
rect 5809 6352 5875 6357
rect 5809 6296 5814 6352
rect 5870 6296 5875 6352
rect 5809 6291 5875 6296
rect 4705 6218 4771 6221
rect 6310 6218 6316 6220
rect 4705 6216 6316 6218
rect 4705 6160 4710 6216
rect 4766 6160 6316 6216
rect 4705 6158 6316 6160
rect 4705 6155 4771 6158
rect 6310 6156 6316 6158
rect 6380 6156 6386 6220
rect 2129 6082 2195 6085
rect 4102 6082 4108 6084
rect 2129 6080 4108 6082
rect 2129 6024 2134 6080
rect 2190 6024 4108 6080
rect 2129 6022 4108 6024
rect 2129 6019 2195 6022
rect 4102 6020 4108 6022
rect 4172 6020 4178 6084
rect 4685 6016 5005 6017
rect 4685 5952 4693 6016
rect 4757 5952 4773 6016
rect 4837 5952 4853 6016
rect 4917 5952 4933 6016
rect 4997 5952 5005 6016
rect 4685 5951 5005 5952
rect 8426 6016 8746 6017
rect 8426 5952 8434 6016
rect 8498 5952 8514 6016
rect 8578 5952 8594 6016
rect 8658 5952 8674 6016
rect 8738 5952 8746 6016
rect 8426 5951 8746 5952
rect 4102 5884 4108 5948
rect 4172 5946 4178 5948
rect 4429 5946 4495 5949
rect 4172 5944 4495 5946
rect 4172 5888 4434 5944
rect 4490 5888 4495 5944
rect 4172 5886 4495 5888
rect 4172 5884 4178 5886
rect 4429 5883 4495 5886
rect 1393 5674 1459 5677
rect 1526 5674 1532 5676
rect 1393 5672 1532 5674
rect 1393 5616 1398 5672
rect 1454 5616 1532 5672
rect 1393 5614 1532 5616
rect 1393 5611 1459 5614
rect 1526 5612 1532 5614
rect 1596 5612 1602 5676
rect 2814 5472 3134 5473
rect 2814 5408 2822 5472
rect 2886 5408 2902 5472
rect 2966 5408 2982 5472
rect 3046 5408 3062 5472
rect 3126 5408 3134 5472
rect 2814 5407 3134 5408
rect 6556 5472 6876 5473
rect 6556 5408 6564 5472
rect 6628 5408 6644 5472
rect 6708 5408 6724 5472
rect 6788 5408 6804 5472
rect 6868 5408 6876 5472
rect 6556 5407 6876 5408
rect 10297 5472 10617 5473
rect 10297 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10545 5472
rect 10609 5408 10617 5472
rect 10297 5407 10617 5408
rect 7189 5402 7255 5405
rect 7557 5402 7623 5405
rect 7189 5400 7623 5402
rect 7189 5344 7194 5400
rect 7250 5344 7562 5400
rect 7618 5344 7623 5400
rect 7189 5342 7623 5344
rect 7189 5339 7255 5342
rect 7557 5339 7623 5342
rect 3969 5266 4035 5269
rect 7557 5266 7623 5269
rect 3969 5264 7623 5266
rect 3969 5208 3974 5264
rect 4030 5208 7562 5264
rect 7618 5208 7623 5264
rect 3969 5206 7623 5208
rect 3969 5203 4035 5206
rect 7557 5203 7623 5206
rect 8150 5204 8156 5268
rect 8220 5266 8226 5268
rect 8937 5266 9003 5269
rect 8220 5264 9003 5266
rect 8220 5208 8942 5264
rect 8998 5208 9003 5264
rect 8220 5206 9003 5208
rect 8220 5204 8226 5206
rect 8937 5203 9003 5206
rect 6126 5130 6132 5132
rect 4524 5070 6132 5130
rect 2446 4796 2452 4860
rect 2516 4858 2522 4860
rect 2681 4858 2747 4861
rect 2516 4856 2747 4858
rect 2516 4800 2686 4856
rect 2742 4800 2747 4856
rect 2516 4798 2747 4800
rect 2516 4796 2522 4798
rect 2681 4795 2747 4798
rect 3417 4858 3483 4861
rect 4524 4858 4584 5070
rect 6126 5068 6132 5070
rect 6196 5068 6202 5132
rect 6269 5130 6335 5133
rect 8201 5130 8267 5133
rect 6269 5128 8267 5130
rect 6269 5072 6274 5128
rect 6330 5072 8206 5128
rect 8262 5072 8267 5128
rect 6269 5070 8267 5072
rect 6269 5067 6335 5070
rect 8201 5067 8267 5070
rect 9857 5130 9923 5133
rect 10961 5130 11027 5133
rect 9857 5128 11027 5130
rect 9857 5072 9862 5128
rect 9918 5072 10966 5128
rect 11022 5072 11027 5128
rect 9857 5070 11027 5072
rect 9857 5067 9923 5070
rect 10961 5067 11027 5070
rect 5441 4994 5507 4997
rect 7966 4994 7972 4996
rect 5441 4992 7972 4994
rect 5441 4936 5446 4992
rect 5502 4936 7972 4992
rect 5441 4934 7972 4936
rect 5441 4931 5507 4934
rect 7966 4932 7972 4934
rect 8036 4932 8042 4996
rect 10593 4994 10659 4997
rect 10726 4994 10732 4996
rect 10593 4992 10732 4994
rect 10593 4936 10598 4992
rect 10654 4936 10732 4992
rect 10593 4934 10732 4936
rect 10593 4931 10659 4934
rect 10726 4932 10732 4934
rect 10796 4932 10802 4996
rect 4685 4928 5005 4929
rect 4685 4864 4693 4928
rect 4757 4864 4773 4928
rect 4837 4864 4853 4928
rect 4917 4864 4933 4928
rect 4997 4864 5005 4928
rect 4685 4863 5005 4864
rect 8426 4928 8746 4929
rect 8426 4864 8434 4928
rect 8498 4864 8514 4928
rect 8578 4864 8594 4928
rect 8658 4864 8674 4928
rect 8738 4864 8746 4928
rect 8426 4863 8746 4864
rect 3417 4856 4584 4858
rect 3417 4800 3422 4856
rect 3478 4800 4584 4856
rect 3417 4798 4584 4800
rect 5441 4858 5507 4861
rect 6913 4858 6979 4861
rect 5441 4856 6979 4858
rect 5441 4800 5446 4856
rect 5502 4800 6918 4856
rect 6974 4800 6979 4856
rect 5441 4798 6979 4800
rect 3417 4795 3483 4798
rect 5441 4795 5507 4798
rect 6913 4795 6979 4798
rect 4470 4660 4476 4724
rect 4540 4722 4546 4724
rect 9489 4722 9555 4725
rect 4540 4720 9555 4722
rect 4540 4664 9494 4720
rect 9550 4664 9555 4720
rect 4540 4662 9555 4664
rect 4540 4660 4546 4662
rect 9489 4659 9555 4662
rect 2446 4524 2452 4588
rect 2516 4586 2522 4588
rect 3969 4586 4035 4589
rect 2516 4584 4035 4586
rect 2516 4528 3974 4584
rect 4030 4528 4035 4584
rect 2516 4526 4035 4528
rect 2516 4524 2522 4526
rect 3969 4523 4035 4526
rect 4337 4586 4403 4589
rect 5809 4586 5875 4589
rect 4337 4584 5875 4586
rect 4337 4528 4342 4584
rect 4398 4528 5814 4584
rect 5870 4528 5875 4584
rect 4337 4526 5875 4528
rect 4337 4523 4403 4526
rect 5809 4523 5875 4526
rect 6085 4584 6151 4589
rect 6085 4528 6090 4584
rect 6146 4528 6151 4584
rect 6085 4523 6151 4528
rect 6545 4586 6611 4589
rect 7925 4586 7991 4589
rect 8109 4586 8175 4589
rect 6545 4584 7114 4586
rect 6545 4528 6550 4584
rect 6606 4528 7114 4584
rect 6545 4526 7114 4528
rect 6545 4523 6611 4526
rect 5809 4450 5875 4453
rect 5628 4448 5875 4450
rect 5628 4392 5814 4448
rect 5870 4392 5875 4448
rect 5628 4390 5875 4392
rect 2814 4384 3134 4385
rect 2814 4320 2822 4384
rect 2886 4320 2902 4384
rect 2966 4320 2982 4384
rect 3046 4320 3062 4384
rect 3126 4320 3134 4384
rect 2814 4319 3134 4320
rect 749 4042 815 4045
rect 1158 4042 1164 4044
rect 749 4040 1164 4042
rect 749 3984 754 4040
rect 810 3984 1164 4040
rect 749 3982 1164 3984
rect 749 3979 815 3982
rect 1158 3980 1164 3982
rect 1228 3980 1234 4044
rect 4889 4042 4955 4045
rect 4889 4040 5228 4042
rect 4889 3984 4894 4040
rect 4950 3984 5228 4040
rect 4889 3982 5228 3984
rect 4889 3979 4955 3982
rect 3693 3906 3759 3909
rect 4470 3906 4476 3908
rect 3693 3904 4476 3906
rect 3693 3848 3698 3904
rect 3754 3848 4476 3904
rect 3693 3846 4476 3848
rect 3693 3843 3759 3846
rect 4470 3844 4476 3846
rect 4540 3844 4546 3908
rect 4685 3840 5005 3841
rect 4685 3776 4693 3840
rect 4757 3776 4773 3840
rect 4837 3776 4853 3840
rect 4917 3776 4933 3840
rect 4997 3776 5005 3840
rect 4685 3775 5005 3776
rect 4061 3770 4127 3773
rect 4429 3770 4495 3773
rect 4061 3768 4495 3770
rect 4061 3712 4066 3768
rect 4122 3712 4434 3768
rect 4490 3712 4495 3768
rect 4061 3710 4495 3712
rect 4061 3707 4127 3710
rect 4429 3707 4495 3710
rect 2313 3634 2379 3637
rect 4705 3634 4771 3637
rect 2313 3632 4771 3634
rect 2313 3576 2318 3632
rect 2374 3576 4710 3632
rect 4766 3576 4771 3632
rect 2313 3574 4771 3576
rect 2313 3571 2379 3574
rect 4705 3571 4771 3574
rect 4889 3634 4955 3637
rect 5168 3634 5228 3982
rect 4889 3632 5228 3634
rect 4889 3576 4894 3632
rect 4950 3576 5228 3632
rect 4889 3574 5228 3576
rect 4889 3571 4955 3574
rect 2313 3500 2379 3501
rect 2262 3436 2268 3500
rect 2332 3498 2379 3500
rect 3049 3498 3115 3501
rect 5390 3498 5396 3500
rect 2332 3496 2424 3498
rect 2374 3440 2424 3496
rect 2332 3438 2424 3440
rect 3049 3496 5396 3498
rect 3049 3440 3054 3496
rect 3110 3440 5396 3496
rect 3049 3438 5396 3440
rect 2332 3436 2379 3438
rect 2313 3435 2379 3436
rect 3049 3435 3115 3438
rect 5390 3436 5396 3438
rect 5460 3436 5466 3500
rect 3969 3362 4035 3365
rect 3969 3360 4170 3362
rect 3969 3304 3974 3360
rect 4030 3304 4170 3360
rect 3969 3302 4170 3304
rect 3969 3299 4035 3302
rect 2814 3296 3134 3297
rect 2814 3232 2822 3296
rect 2886 3232 2902 3296
rect 2966 3232 2982 3296
rect 3046 3232 3062 3296
rect 3126 3232 3134 3296
rect 2814 3231 3134 3232
rect 4110 3093 4170 3302
rect 5257 3226 5323 3229
rect 5390 3226 5396 3228
rect 5257 3224 5396 3226
rect 5257 3168 5262 3224
rect 5318 3168 5396 3224
rect 5257 3166 5396 3168
rect 5257 3163 5323 3166
rect 5390 3164 5396 3166
rect 5460 3164 5466 3228
rect 3049 3090 3115 3093
rect 3734 3090 3740 3092
rect 3049 3088 3740 3090
rect 3049 3032 3054 3088
rect 3110 3032 3740 3088
rect 3049 3030 3740 3032
rect 3049 3027 3115 3030
rect 3734 3028 3740 3030
rect 3804 3028 3810 3092
rect 4110 3088 4219 3093
rect 4110 3032 4158 3088
rect 4214 3032 4219 3088
rect 4110 3030 4219 3032
rect 4153 3027 4219 3030
rect 4470 3028 4476 3092
rect 4540 3090 4546 3092
rect 4797 3090 4863 3093
rect 4540 3088 4863 3090
rect 4540 3032 4802 3088
rect 4858 3032 4863 3088
rect 4540 3030 4863 3032
rect 5628 3090 5688 4390
rect 5809 4387 5875 4390
rect 6088 4314 6148 4523
rect 7054 4450 7114 4526
rect 7925 4584 8175 4586
rect 7925 4528 7930 4584
rect 7986 4528 8114 4584
rect 8170 4528 8175 4584
rect 7925 4526 8175 4528
rect 7925 4523 7991 4526
rect 8109 4523 8175 4526
rect 9070 4524 9076 4588
rect 9140 4586 9146 4588
rect 9305 4586 9371 4589
rect 9140 4584 9371 4586
rect 9140 4528 9310 4584
rect 9366 4528 9371 4584
rect 9140 4526 9371 4528
rect 9140 4524 9146 4526
rect 9305 4523 9371 4526
rect 9581 4450 9647 4453
rect 7054 4448 9647 4450
rect 7054 4392 9586 4448
rect 9642 4392 9647 4448
rect 7054 4390 9647 4392
rect 9581 4387 9647 4390
rect 6556 4384 6876 4385
rect 6556 4320 6564 4384
rect 6628 4320 6644 4384
rect 6708 4320 6724 4384
rect 6788 4320 6804 4384
rect 6868 4320 6876 4384
rect 6556 4319 6876 4320
rect 10297 4384 10617 4385
rect 10297 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10545 4384
rect 10609 4320 10617 4384
rect 10297 4319 10617 4320
rect 5766 4254 6148 4314
rect 8569 4314 8635 4317
rect 8569 4312 9920 4314
rect 8569 4256 8574 4312
rect 8630 4256 9920 4312
rect 8569 4254 9920 4256
rect 5766 3906 5826 4254
rect 8569 4251 8635 4254
rect 5901 4178 5967 4181
rect 7373 4178 7439 4181
rect 8661 4178 8727 4181
rect 5901 4176 7439 4178
rect 5901 4120 5906 4176
rect 5962 4120 7378 4176
rect 7434 4120 7439 4176
rect 5901 4118 7439 4120
rect 5901 4115 5967 4118
rect 7373 4115 7439 4118
rect 7974 4176 8727 4178
rect 7974 4120 8666 4176
rect 8722 4120 8727 4176
rect 7974 4118 8727 4120
rect 6085 4042 6151 4045
rect 7974 4042 8034 4118
rect 8661 4115 8727 4118
rect 9305 4178 9371 4181
rect 9581 4178 9647 4181
rect 9305 4176 9647 4178
rect 9305 4120 9310 4176
rect 9366 4120 9586 4176
rect 9642 4120 9647 4176
rect 9305 4118 9647 4120
rect 9860 4178 9920 4254
rect 10869 4178 10935 4181
rect 12065 4178 12131 4181
rect 9860 4176 10935 4178
rect 9860 4120 10874 4176
rect 10930 4120 10935 4176
rect 9860 4118 10935 4120
rect 9305 4115 9371 4118
rect 9581 4115 9647 4118
rect 10869 4115 10935 4118
rect 11102 4176 12131 4178
rect 11102 4120 12070 4176
rect 12126 4120 12131 4176
rect 11102 4118 12131 4120
rect 6085 4040 8034 4042
rect 6085 3984 6090 4040
rect 6146 3984 8034 4040
rect 6085 3982 8034 3984
rect 8109 4042 8175 4045
rect 9305 4042 9371 4045
rect 8109 4040 9371 4042
rect 8109 3984 8114 4040
rect 8170 3984 9310 4040
rect 9366 3984 9371 4040
rect 8109 3982 9371 3984
rect 6085 3979 6151 3982
rect 8109 3979 8175 3982
rect 9305 3979 9371 3982
rect 10317 4042 10383 4045
rect 11102 4042 11162 4118
rect 12065 4115 12131 4118
rect 10317 4040 11162 4042
rect 10317 3984 10322 4040
rect 10378 3984 11162 4040
rect 10317 3982 11162 3984
rect 10317 3979 10383 3982
rect 6821 3906 6887 3909
rect 5766 3904 6887 3906
rect 5766 3848 6826 3904
rect 6882 3848 6887 3904
rect 5766 3846 6887 3848
rect 6821 3843 6887 3846
rect 8426 3840 8746 3841
rect 8426 3776 8434 3840
rect 8498 3776 8514 3840
rect 8578 3776 8594 3840
rect 8658 3776 8674 3840
rect 8738 3776 8746 3840
rect 8426 3775 8746 3776
rect 9673 3770 9739 3773
rect 9806 3770 9812 3772
rect 9673 3768 9812 3770
rect 9673 3712 9678 3768
rect 9734 3712 9812 3768
rect 9673 3710 9812 3712
rect 9673 3707 9739 3710
rect 9806 3708 9812 3710
rect 9876 3708 9882 3772
rect 5809 3634 5875 3637
rect 6269 3634 6335 3637
rect 5809 3632 6335 3634
rect 5809 3576 5814 3632
rect 5870 3576 6274 3632
rect 6330 3576 6335 3632
rect 5809 3574 6335 3576
rect 5809 3571 5875 3574
rect 6269 3571 6335 3574
rect 7281 3634 7347 3637
rect 11789 3634 11855 3637
rect 7281 3632 11855 3634
rect 7281 3576 7286 3632
rect 7342 3576 11794 3632
rect 11850 3576 11855 3632
rect 7281 3574 11855 3576
rect 7281 3571 7347 3574
rect 11789 3571 11855 3574
rect 6453 3498 6519 3501
rect 7465 3498 7531 3501
rect 6453 3496 7531 3498
rect 6453 3440 6458 3496
rect 6514 3440 7470 3496
rect 7526 3440 7531 3496
rect 6453 3438 7531 3440
rect 6453 3435 6519 3438
rect 7465 3435 7531 3438
rect 8293 3498 8359 3501
rect 8937 3498 9003 3501
rect 8293 3496 9003 3498
rect 8293 3440 8298 3496
rect 8354 3440 8942 3496
rect 8998 3440 9003 3496
rect 8293 3438 9003 3440
rect 8293 3435 8359 3438
rect 8937 3435 9003 3438
rect 8109 3362 8175 3365
rect 9622 3362 9628 3364
rect 8109 3360 9628 3362
rect 8109 3304 8114 3360
rect 8170 3304 9628 3360
rect 8109 3302 9628 3304
rect 8109 3299 8175 3302
rect 9622 3300 9628 3302
rect 9692 3300 9698 3364
rect 6556 3296 6876 3297
rect 6556 3232 6564 3296
rect 6628 3232 6644 3296
rect 6708 3232 6724 3296
rect 6788 3232 6804 3296
rect 6868 3232 6876 3296
rect 6556 3231 6876 3232
rect 10297 3296 10617 3297
rect 10297 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10545 3296
rect 10609 3232 10617 3296
rect 10297 3231 10617 3232
rect 7281 3226 7347 3229
rect 8661 3226 8727 3229
rect 7281 3224 8727 3226
rect 7281 3168 7286 3224
rect 7342 3168 8666 3224
rect 8722 3168 8727 3224
rect 7281 3166 8727 3168
rect 7281 3163 7347 3166
rect 8661 3163 8727 3166
rect 11329 3226 11395 3229
rect 11605 3226 11671 3229
rect 11329 3224 11671 3226
rect 11329 3168 11334 3224
rect 11390 3168 11610 3224
rect 11666 3168 11671 3224
rect 11329 3166 11671 3168
rect 11329 3163 11395 3166
rect 11605 3163 11671 3166
rect 10961 3090 11027 3093
rect 5628 3088 11027 3090
rect 5628 3032 10966 3088
rect 11022 3032 11027 3088
rect 5628 3030 11027 3032
rect 4540 3028 4546 3030
rect 4797 3027 4863 3030
rect 10961 3027 11027 3030
rect 2446 2892 2452 2956
rect 2516 2954 2522 2956
rect 3141 2954 3207 2957
rect 2516 2952 3207 2954
rect 2516 2896 3146 2952
rect 3202 2896 3207 2952
rect 2516 2894 3207 2896
rect 2516 2892 2522 2894
rect 3141 2891 3207 2894
rect 3693 2954 3759 2957
rect 4286 2954 4292 2956
rect 3693 2952 4292 2954
rect 3693 2896 3698 2952
rect 3754 2896 4292 2952
rect 3693 2894 4292 2896
rect 3693 2891 3759 2894
rect 4286 2892 4292 2894
rect 4356 2892 4362 2956
rect 4521 2954 4587 2957
rect 5257 2956 5323 2957
rect 4478 2952 4587 2954
rect 4478 2896 4526 2952
rect 4582 2896 4587 2952
rect 4478 2891 4587 2896
rect 5206 2892 5212 2956
rect 5276 2954 5323 2956
rect 5625 2954 5691 2957
rect 6821 2954 6887 2957
rect 5276 2952 5368 2954
rect 5318 2896 5368 2952
rect 5276 2894 5368 2896
rect 5625 2952 6887 2954
rect 5625 2896 5630 2952
rect 5686 2896 6826 2952
rect 6882 2896 6887 2952
rect 5625 2894 6887 2896
rect 5276 2892 5323 2894
rect 5257 2891 5323 2892
rect 5625 2891 5691 2894
rect 6821 2891 6887 2894
rect 7189 2954 7255 2957
rect 8150 2954 8156 2956
rect 7189 2952 8156 2954
rect 7189 2896 7194 2952
rect 7250 2896 8156 2952
rect 7189 2894 8156 2896
rect 7189 2891 7255 2894
rect 8150 2892 8156 2894
rect 8220 2892 8226 2956
rect 9070 2954 9076 2956
rect 8296 2894 9076 2954
rect 933 2818 999 2821
rect 2037 2818 2103 2821
rect 933 2816 2103 2818
rect 933 2760 938 2816
rect 994 2760 2042 2816
rect 2098 2760 2103 2816
rect 933 2758 2103 2760
rect 933 2755 999 2758
rect 2037 2755 2103 2758
rect 3049 2682 3115 2685
rect 4478 2682 4538 2891
rect 7046 2818 7052 2820
rect 5214 2758 7052 2818
rect 4685 2752 5005 2753
rect 4685 2688 4693 2752
rect 4757 2688 4773 2752
rect 4837 2688 4853 2752
rect 4917 2688 4933 2752
rect 4997 2688 5005 2752
rect 4685 2687 5005 2688
rect 3049 2680 4538 2682
rect 3049 2624 3054 2680
rect 3110 2624 4538 2680
rect 3049 2622 4538 2624
rect 3049 2619 3115 2622
rect 3325 2548 3391 2549
rect 3325 2546 3372 2548
rect 3280 2544 3372 2546
rect 3280 2488 3330 2544
rect 3280 2486 3372 2488
rect 3325 2484 3372 2486
rect 3436 2484 3442 2548
rect 4429 2546 4495 2549
rect 5214 2546 5274 2758
rect 7046 2756 7052 2758
rect 7116 2756 7122 2820
rect 7925 2818 7991 2821
rect 8296 2818 8356 2894
rect 9070 2892 9076 2894
rect 9140 2892 9146 2956
rect 9857 2954 9923 2957
rect 9990 2954 9996 2956
rect 9857 2952 9996 2954
rect 9857 2896 9862 2952
rect 9918 2896 9996 2952
rect 9857 2894 9996 2896
rect 9857 2891 9923 2894
rect 9990 2892 9996 2894
rect 10060 2892 10066 2956
rect 7925 2816 8356 2818
rect 7925 2760 7930 2816
rect 7986 2760 8356 2816
rect 7925 2758 8356 2760
rect 11237 2818 11303 2821
rect 11789 2818 11855 2821
rect 11237 2816 11855 2818
rect 11237 2760 11242 2816
rect 11298 2760 11794 2816
rect 11850 2760 11855 2816
rect 11237 2758 11855 2760
rect 7925 2755 7991 2758
rect 11237 2755 11303 2758
rect 11789 2755 11855 2758
rect 8426 2752 8746 2753
rect 8426 2688 8434 2752
rect 8498 2688 8514 2752
rect 8578 2688 8594 2752
rect 8658 2688 8674 2752
rect 8738 2688 8746 2752
rect 8426 2687 8746 2688
rect 5625 2548 5691 2549
rect 4429 2544 5274 2546
rect 4429 2488 4434 2544
rect 4490 2488 5274 2544
rect 4429 2486 5274 2488
rect 3325 2483 3391 2484
rect 4429 2483 4495 2486
rect 5574 2484 5580 2548
rect 5644 2546 5691 2548
rect 8385 2546 8451 2549
rect 8886 2546 8892 2548
rect 5644 2544 5736 2546
rect 5686 2488 5736 2544
rect 5644 2486 5736 2488
rect 8385 2544 8892 2546
rect 8385 2488 8390 2544
rect 8446 2488 8892 2544
rect 8385 2486 8892 2488
rect 5644 2484 5691 2486
rect 5625 2483 5691 2484
rect 8385 2483 8451 2486
rect 8886 2484 8892 2486
rect 8956 2484 8962 2548
rect 5165 2410 5231 2413
rect 5390 2410 5396 2412
rect 5165 2408 5396 2410
rect 5165 2352 5170 2408
rect 5226 2352 5396 2408
rect 5165 2350 5396 2352
rect 5165 2347 5231 2350
rect 5390 2348 5396 2350
rect 5460 2348 5466 2412
rect 7966 2348 7972 2412
rect 8036 2410 8042 2412
rect 8661 2410 8727 2413
rect 8036 2408 8727 2410
rect 8036 2352 8666 2408
rect 8722 2352 8727 2408
rect 8036 2350 8727 2352
rect 8036 2348 8042 2350
rect 8661 2347 8727 2350
rect 4061 2274 4127 2277
rect 5758 2274 5764 2276
rect 4061 2272 5764 2274
rect 4061 2216 4066 2272
rect 4122 2216 5764 2272
rect 4061 2214 5764 2216
rect 4061 2211 4127 2214
rect 5758 2212 5764 2214
rect 5828 2212 5834 2276
rect 7414 2212 7420 2276
rect 7484 2274 7490 2276
rect 8845 2274 8911 2277
rect 7484 2272 8911 2274
rect 7484 2216 8850 2272
rect 8906 2216 8911 2272
rect 7484 2214 8911 2216
rect 7484 2212 7490 2214
rect 8845 2211 8911 2214
rect 2814 2208 3134 2209
rect 2814 2144 2822 2208
rect 2886 2144 2902 2208
rect 2966 2144 2982 2208
rect 3046 2144 3062 2208
rect 3126 2144 3134 2208
rect 2814 2143 3134 2144
rect 6556 2208 6876 2209
rect 6556 2144 6564 2208
rect 6628 2144 6644 2208
rect 6708 2144 6724 2208
rect 6788 2144 6804 2208
rect 6868 2144 6876 2208
rect 6556 2143 6876 2144
rect 10297 2208 10617 2209
rect 10297 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10545 2208
rect 10609 2144 10617 2208
rect 10297 2143 10617 2144
rect 5942 1940 5948 2004
rect 6012 2002 6018 2004
rect 8753 2002 8819 2005
rect 6012 2000 8819 2002
rect 6012 1944 8758 2000
rect 8814 1944 8819 2000
rect 6012 1942 8819 1944
rect 6012 1940 6018 1942
rect 8753 1939 8819 1942
rect 4102 1804 4108 1868
rect 4172 1866 4178 1868
rect 7189 1866 7255 1869
rect 4172 1864 7255 1866
rect 4172 1808 7194 1864
rect 7250 1808 7255 1864
rect 4172 1806 7255 1808
rect 4172 1804 4178 1806
rect 7189 1803 7255 1806
rect 4889 1730 4955 1733
rect 7598 1730 7604 1732
rect 4889 1728 7604 1730
rect 4889 1672 4894 1728
rect 4950 1672 7604 1728
rect 4889 1670 7604 1672
rect 4889 1667 4955 1670
rect 7598 1668 7604 1670
rect 7668 1668 7674 1732
rect 2630 1532 2636 1596
rect 2700 1594 2706 1596
rect 5441 1594 5507 1597
rect 2700 1592 5507 1594
rect 2700 1536 5446 1592
rect 5502 1536 5507 1592
rect 2700 1534 5507 1536
rect 2700 1532 2706 1534
rect 5441 1531 5507 1534
rect 6310 1532 6316 1596
rect 6380 1594 6386 1596
rect 8477 1594 8543 1597
rect 6380 1592 8543 1594
rect 6380 1536 8482 1592
rect 8538 1536 8543 1592
rect 6380 1534 8543 1536
rect 6380 1532 6386 1534
rect 8477 1531 8543 1534
rect 7230 1458 7236 1460
rect 3696 1398 7236 1458
rect 3696 1325 3756 1398
rect 7230 1396 7236 1398
rect 7300 1396 7306 1460
rect 3693 1320 3759 1325
rect 3693 1264 3698 1320
rect 3754 1264 3759 1320
rect 3693 1259 3759 1264
rect 6126 1260 6132 1324
rect 6196 1322 6202 1324
rect 6729 1322 6795 1325
rect 6196 1320 6795 1322
rect 6196 1264 6734 1320
rect 6790 1264 6795 1320
rect 6196 1262 6795 1264
rect 6196 1260 6202 1262
rect 6729 1259 6795 1262
rect 3550 1124 3556 1188
rect 3620 1186 3626 1188
rect 4245 1186 4311 1189
rect 3620 1184 4311 1186
rect 3620 1128 4250 1184
rect 4306 1128 4311 1184
rect 3620 1126 4311 1128
rect 3620 1124 3626 1126
rect 4245 1123 4311 1126
rect 9806 1124 9812 1188
rect 9876 1186 9882 1188
rect 10041 1186 10107 1189
rect 9876 1184 10107 1186
rect 9876 1128 10046 1184
rect 10102 1128 10107 1184
rect 9876 1126 10107 1128
rect 9876 1124 9882 1126
rect 10041 1123 10107 1126
rect 4613 1050 4679 1053
rect 7782 1050 7788 1052
rect 4613 1048 7788 1050
rect 4613 992 4618 1048
rect 4674 992 7788 1048
rect 4613 990 7788 992
rect 4613 987 4679 990
rect 7782 988 7788 990
rect 7852 988 7858 1052
rect 3918 852 3924 916
rect 3988 914 3994 916
rect 5901 914 5967 917
rect 3988 912 5967 914
rect 3988 856 5906 912
rect 5962 856 5967 912
rect 3988 854 5967 856
rect 3988 852 3994 854
rect 5901 851 5967 854
<< via3 >>
rect 2822 13084 2886 13088
rect 2822 13028 2826 13084
rect 2826 13028 2882 13084
rect 2882 13028 2886 13084
rect 2822 13024 2886 13028
rect 2902 13084 2966 13088
rect 2902 13028 2906 13084
rect 2906 13028 2962 13084
rect 2962 13028 2966 13084
rect 2902 13024 2966 13028
rect 2982 13084 3046 13088
rect 2982 13028 2986 13084
rect 2986 13028 3042 13084
rect 3042 13028 3046 13084
rect 2982 13024 3046 13028
rect 3062 13084 3126 13088
rect 3062 13028 3066 13084
rect 3066 13028 3122 13084
rect 3122 13028 3126 13084
rect 3062 13024 3126 13028
rect 6564 13084 6628 13088
rect 6564 13028 6568 13084
rect 6568 13028 6624 13084
rect 6624 13028 6628 13084
rect 6564 13024 6628 13028
rect 6644 13084 6708 13088
rect 6644 13028 6648 13084
rect 6648 13028 6704 13084
rect 6704 13028 6708 13084
rect 6644 13024 6708 13028
rect 6724 13084 6788 13088
rect 6724 13028 6728 13084
rect 6728 13028 6784 13084
rect 6784 13028 6788 13084
rect 6724 13024 6788 13028
rect 6804 13084 6868 13088
rect 6804 13028 6808 13084
rect 6808 13028 6864 13084
rect 6864 13028 6868 13084
rect 6804 13024 6868 13028
rect 10305 13084 10369 13088
rect 10305 13028 10309 13084
rect 10309 13028 10365 13084
rect 10365 13028 10369 13084
rect 10305 13024 10369 13028
rect 10385 13084 10449 13088
rect 10385 13028 10389 13084
rect 10389 13028 10445 13084
rect 10445 13028 10449 13084
rect 10385 13024 10449 13028
rect 10465 13084 10529 13088
rect 10465 13028 10469 13084
rect 10469 13028 10525 13084
rect 10525 13028 10529 13084
rect 10465 13024 10529 13028
rect 10545 13084 10609 13088
rect 10545 13028 10549 13084
rect 10549 13028 10605 13084
rect 10605 13028 10609 13084
rect 10545 13024 10609 13028
rect 1164 12820 1228 12884
rect 4693 12540 4757 12544
rect 4693 12484 4697 12540
rect 4697 12484 4753 12540
rect 4753 12484 4757 12540
rect 4693 12480 4757 12484
rect 4773 12540 4837 12544
rect 4773 12484 4777 12540
rect 4777 12484 4833 12540
rect 4833 12484 4837 12540
rect 4773 12480 4837 12484
rect 4853 12540 4917 12544
rect 4853 12484 4857 12540
rect 4857 12484 4913 12540
rect 4913 12484 4917 12540
rect 4853 12480 4917 12484
rect 4933 12540 4997 12544
rect 4933 12484 4937 12540
rect 4937 12484 4993 12540
rect 4993 12484 4997 12540
rect 4933 12480 4997 12484
rect 8434 12540 8498 12544
rect 8434 12484 8438 12540
rect 8438 12484 8494 12540
rect 8494 12484 8498 12540
rect 8434 12480 8498 12484
rect 8514 12540 8578 12544
rect 8514 12484 8518 12540
rect 8518 12484 8574 12540
rect 8574 12484 8578 12540
rect 8514 12480 8578 12484
rect 8594 12540 8658 12544
rect 8594 12484 8598 12540
rect 8598 12484 8654 12540
rect 8654 12484 8658 12540
rect 8594 12480 8658 12484
rect 8674 12540 8738 12544
rect 8674 12484 8678 12540
rect 8678 12484 8734 12540
rect 8734 12484 8738 12540
rect 8674 12480 8738 12484
rect 2822 11996 2886 12000
rect 2822 11940 2826 11996
rect 2826 11940 2882 11996
rect 2882 11940 2886 11996
rect 2822 11936 2886 11940
rect 2902 11996 2966 12000
rect 2902 11940 2906 11996
rect 2906 11940 2962 11996
rect 2962 11940 2966 11996
rect 2902 11936 2966 11940
rect 2982 11996 3046 12000
rect 2982 11940 2986 11996
rect 2986 11940 3042 11996
rect 3042 11940 3046 11996
rect 2982 11936 3046 11940
rect 3062 11996 3126 12000
rect 3062 11940 3066 11996
rect 3066 11940 3122 11996
rect 3122 11940 3126 11996
rect 3062 11936 3126 11940
rect 6564 11996 6628 12000
rect 6564 11940 6568 11996
rect 6568 11940 6624 11996
rect 6624 11940 6628 11996
rect 6564 11936 6628 11940
rect 6644 11996 6708 12000
rect 6644 11940 6648 11996
rect 6648 11940 6704 11996
rect 6704 11940 6708 11996
rect 6644 11936 6708 11940
rect 6724 11996 6788 12000
rect 6724 11940 6728 11996
rect 6728 11940 6784 11996
rect 6784 11940 6788 11996
rect 6724 11936 6788 11940
rect 6804 11996 6868 12000
rect 6804 11940 6808 11996
rect 6808 11940 6864 11996
rect 6864 11940 6868 11996
rect 6804 11936 6868 11940
rect 10305 11996 10369 12000
rect 10305 11940 10309 11996
rect 10309 11940 10365 11996
rect 10365 11940 10369 11996
rect 10305 11936 10369 11940
rect 10385 11996 10449 12000
rect 10385 11940 10389 11996
rect 10389 11940 10445 11996
rect 10445 11940 10449 11996
rect 10385 11936 10449 11940
rect 10465 11996 10529 12000
rect 10465 11940 10469 11996
rect 10469 11940 10525 11996
rect 10525 11940 10529 11996
rect 10465 11936 10529 11940
rect 10545 11996 10609 12000
rect 10545 11940 10549 11996
rect 10549 11940 10605 11996
rect 10605 11940 10609 11996
rect 10545 11936 10609 11940
rect 4693 11452 4757 11456
rect 4693 11396 4697 11452
rect 4697 11396 4753 11452
rect 4753 11396 4757 11452
rect 4693 11392 4757 11396
rect 4773 11452 4837 11456
rect 4773 11396 4777 11452
rect 4777 11396 4833 11452
rect 4833 11396 4837 11452
rect 4773 11392 4837 11396
rect 4853 11452 4917 11456
rect 4853 11396 4857 11452
rect 4857 11396 4913 11452
rect 4913 11396 4917 11452
rect 4853 11392 4917 11396
rect 4933 11452 4997 11456
rect 4933 11396 4937 11452
rect 4937 11396 4993 11452
rect 4993 11396 4997 11452
rect 4933 11392 4997 11396
rect 8434 11452 8498 11456
rect 8434 11396 8438 11452
rect 8438 11396 8494 11452
rect 8494 11396 8498 11452
rect 8434 11392 8498 11396
rect 8514 11452 8578 11456
rect 8514 11396 8518 11452
rect 8518 11396 8574 11452
rect 8574 11396 8578 11452
rect 8514 11392 8578 11396
rect 8594 11452 8658 11456
rect 8594 11396 8598 11452
rect 8598 11396 8654 11452
rect 8654 11396 8658 11452
rect 8594 11392 8658 11396
rect 8674 11452 8738 11456
rect 8674 11396 8678 11452
rect 8678 11396 8734 11452
rect 8734 11396 8738 11452
rect 8674 11392 8738 11396
rect 7236 11188 7300 11252
rect 7604 11188 7668 11252
rect 5764 11112 5828 11116
rect 5764 11056 5778 11112
rect 5778 11056 5828 11112
rect 5764 11052 5828 11056
rect 7788 11052 7852 11116
rect 2822 10908 2886 10912
rect 2822 10852 2826 10908
rect 2826 10852 2882 10908
rect 2882 10852 2886 10908
rect 2822 10848 2886 10852
rect 2902 10908 2966 10912
rect 2902 10852 2906 10908
rect 2906 10852 2962 10908
rect 2962 10852 2966 10908
rect 2902 10848 2966 10852
rect 2982 10908 3046 10912
rect 2982 10852 2986 10908
rect 2986 10852 3042 10908
rect 3042 10852 3046 10908
rect 2982 10848 3046 10852
rect 3062 10908 3126 10912
rect 3062 10852 3066 10908
rect 3066 10852 3122 10908
rect 3122 10852 3126 10908
rect 3062 10848 3126 10852
rect 6564 10908 6628 10912
rect 6564 10852 6568 10908
rect 6568 10852 6624 10908
rect 6624 10852 6628 10908
rect 6564 10848 6628 10852
rect 6644 10908 6708 10912
rect 6644 10852 6648 10908
rect 6648 10852 6704 10908
rect 6704 10852 6708 10908
rect 6644 10848 6708 10852
rect 6724 10908 6788 10912
rect 6724 10852 6728 10908
rect 6728 10852 6784 10908
rect 6784 10852 6788 10908
rect 6724 10848 6788 10852
rect 6804 10908 6868 10912
rect 6804 10852 6808 10908
rect 6808 10852 6864 10908
rect 6864 10852 6868 10908
rect 6804 10848 6868 10852
rect 10305 10908 10369 10912
rect 10305 10852 10309 10908
rect 10309 10852 10365 10908
rect 10365 10852 10369 10908
rect 10305 10848 10369 10852
rect 10385 10908 10449 10912
rect 10385 10852 10389 10908
rect 10389 10852 10445 10908
rect 10445 10852 10449 10908
rect 10385 10848 10449 10852
rect 10465 10908 10529 10912
rect 10465 10852 10469 10908
rect 10469 10852 10525 10908
rect 10525 10852 10529 10908
rect 10465 10848 10529 10852
rect 10545 10908 10609 10912
rect 10545 10852 10549 10908
rect 10549 10852 10605 10908
rect 10605 10852 10609 10908
rect 10545 10848 10609 10852
rect 4108 10780 4172 10844
rect 4476 10644 4540 10708
rect 4292 10508 4356 10572
rect 8156 10508 8220 10572
rect 4693 10364 4757 10368
rect 4693 10308 4697 10364
rect 4697 10308 4753 10364
rect 4753 10308 4757 10364
rect 4693 10304 4757 10308
rect 4773 10364 4837 10368
rect 4773 10308 4777 10364
rect 4777 10308 4833 10364
rect 4833 10308 4837 10364
rect 4773 10304 4837 10308
rect 4853 10364 4917 10368
rect 4853 10308 4857 10364
rect 4857 10308 4913 10364
rect 4913 10308 4917 10364
rect 4853 10304 4917 10308
rect 4933 10364 4997 10368
rect 4933 10308 4937 10364
rect 4937 10308 4993 10364
rect 4993 10308 4997 10364
rect 4933 10304 4997 10308
rect 8434 10364 8498 10368
rect 8434 10308 8438 10364
rect 8438 10308 8494 10364
rect 8494 10308 8498 10364
rect 8434 10304 8498 10308
rect 8514 10364 8578 10368
rect 8514 10308 8518 10364
rect 8518 10308 8574 10364
rect 8574 10308 8578 10364
rect 8514 10304 8578 10308
rect 8594 10364 8658 10368
rect 8594 10308 8598 10364
rect 8598 10308 8654 10364
rect 8654 10308 8658 10364
rect 8594 10304 8658 10308
rect 8674 10364 8738 10368
rect 8674 10308 8678 10364
rect 8678 10308 8734 10364
rect 8734 10308 8738 10364
rect 8674 10304 8738 10308
rect 7052 10100 7116 10164
rect 3556 9828 3620 9892
rect 2822 9820 2886 9824
rect 2822 9764 2826 9820
rect 2826 9764 2882 9820
rect 2882 9764 2886 9820
rect 2822 9760 2886 9764
rect 2902 9820 2966 9824
rect 2902 9764 2906 9820
rect 2906 9764 2962 9820
rect 2962 9764 2966 9820
rect 2902 9760 2966 9764
rect 2982 9820 3046 9824
rect 2982 9764 2986 9820
rect 2986 9764 3042 9820
rect 3042 9764 3046 9820
rect 2982 9760 3046 9764
rect 3062 9820 3126 9824
rect 3062 9764 3066 9820
rect 3066 9764 3122 9820
rect 3122 9764 3126 9820
rect 3062 9760 3126 9764
rect 6564 9820 6628 9824
rect 6564 9764 6568 9820
rect 6568 9764 6624 9820
rect 6624 9764 6628 9820
rect 6564 9760 6628 9764
rect 6644 9820 6708 9824
rect 6644 9764 6648 9820
rect 6648 9764 6704 9820
rect 6704 9764 6708 9820
rect 6644 9760 6708 9764
rect 6724 9820 6788 9824
rect 6724 9764 6728 9820
rect 6728 9764 6784 9820
rect 6784 9764 6788 9820
rect 6724 9760 6788 9764
rect 6804 9820 6868 9824
rect 6804 9764 6808 9820
rect 6808 9764 6864 9820
rect 6864 9764 6868 9820
rect 6804 9760 6868 9764
rect 10305 9820 10369 9824
rect 10305 9764 10309 9820
rect 10309 9764 10365 9820
rect 10365 9764 10369 9820
rect 10305 9760 10369 9764
rect 10385 9820 10449 9824
rect 10385 9764 10389 9820
rect 10389 9764 10445 9820
rect 10445 9764 10449 9820
rect 10385 9760 10449 9764
rect 10465 9820 10529 9824
rect 10465 9764 10469 9820
rect 10469 9764 10525 9820
rect 10525 9764 10529 9820
rect 10465 9760 10529 9764
rect 10545 9820 10609 9824
rect 10545 9764 10549 9820
rect 10549 9764 10605 9820
rect 10605 9764 10609 9820
rect 10545 9760 10609 9764
rect 8892 9556 8956 9620
rect 3372 9420 3436 9484
rect 4693 9276 4757 9280
rect 4693 9220 4697 9276
rect 4697 9220 4753 9276
rect 4753 9220 4757 9276
rect 4693 9216 4757 9220
rect 4773 9276 4837 9280
rect 4773 9220 4777 9276
rect 4777 9220 4833 9276
rect 4833 9220 4837 9276
rect 4773 9216 4837 9220
rect 4853 9276 4917 9280
rect 4853 9220 4857 9276
rect 4857 9220 4913 9276
rect 4913 9220 4917 9276
rect 4853 9216 4917 9220
rect 4933 9276 4997 9280
rect 4933 9220 4937 9276
rect 4937 9220 4993 9276
rect 4993 9220 4997 9276
rect 4933 9216 4997 9220
rect 8434 9276 8498 9280
rect 8434 9220 8438 9276
rect 8438 9220 8494 9276
rect 8494 9220 8498 9276
rect 8434 9216 8498 9220
rect 8514 9276 8578 9280
rect 8514 9220 8518 9276
rect 8518 9220 8574 9276
rect 8574 9220 8578 9276
rect 8514 9216 8578 9220
rect 8594 9276 8658 9280
rect 8594 9220 8598 9276
rect 8598 9220 8654 9276
rect 8654 9220 8658 9276
rect 8594 9216 8658 9220
rect 8674 9276 8738 9280
rect 8674 9220 8678 9276
rect 8678 9220 8734 9276
rect 8734 9220 8738 9276
rect 8674 9216 8738 9220
rect 1532 9148 1596 9212
rect 5396 9148 5460 9212
rect 7972 8876 8036 8940
rect 2822 8732 2886 8736
rect 2822 8676 2826 8732
rect 2826 8676 2882 8732
rect 2882 8676 2886 8732
rect 2822 8672 2886 8676
rect 2902 8732 2966 8736
rect 2902 8676 2906 8732
rect 2906 8676 2962 8732
rect 2962 8676 2966 8732
rect 2902 8672 2966 8676
rect 2982 8732 3046 8736
rect 2982 8676 2986 8732
rect 2986 8676 3042 8732
rect 3042 8676 3046 8732
rect 2982 8672 3046 8676
rect 3062 8732 3126 8736
rect 3062 8676 3066 8732
rect 3066 8676 3122 8732
rect 3122 8676 3126 8732
rect 3062 8672 3126 8676
rect 6564 8732 6628 8736
rect 6564 8676 6568 8732
rect 6568 8676 6624 8732
rect 6624 8676 6628 8732
rect 6564 8672 6628 8676
rect 6644 8732 6708 8736
rect 6644 8676 6648 8732
rect 6648 8676 6704 8732
rect 6704 8676 6708 8732
rect 6644 8672 6708 8676
rect 6724 8732 6788 8736
rect 6724 8676 6728 8732
rect 6728 8676 6784 8732
rect 6784 8676 6788 8732
rect 6724 8672 6788 8676
rect 6804 8732 6868 8736
rect 6804 8676 6808 8732
rect 6808 8676 6864 8732
rect 6864 8676 6868 8732
rect 6804 8672 6868 8676
rect 10305 8732 10369 8736
rect 10305 8676 10309 8732
rect 10309 8676 10365 8732
rect 10365 8676 10369 8732
rect 10305 8672 10369 8676
rect 10385 8732 10449 8736
rect 10385 8676 10389 8732
rect 10389 8676 10445 8732
rect 10445 8676 10449 8732
rect 10385 8672 10449 8676
rect 10465 8732 10529 8736
rect 10465 8676 10469 8732
rect 10469 8676 10525 8732
rect 10525 8676 10529 8732
rect 10465 8672 10529 8676
rect 10545 8732 10609 8736
rect 10545 8676 10549 8732
rect 10549 8676 10605 8732
rect 10605 8676 10609 8732
rect 10545 8672 10609 8676
rect 2268 8528 2332 8532
rect 2268 8472 2282 8528
rect 2282 8472 2332 8528
rect 2268 8468 2332 8472
rect 5580 8392 5644 8396
rect 5580 8336 5630 8392
rect 5630 8336 5644 8392
rect 5580 8332 5644 8336
rect 4693 8188 4757 8192
rect 4693 8132 4697 8188
rect 4697 8132 4753 8188
rect 4753 8132 4757 8188
rect 4693 8128 4757 8132
rect 4773 8188 4837 8192
rect 4773 8132 4777 8188
rect 4777 8132 4833 8188
rect 4833 8132 4837 8188
rect 4773 8128 4837 8132
rect 4853 8188 4917 8192
rect 4853 8132 4857 8188
rect 4857 8132 4913 8188
rect 4913 8132 4917 8188
rect 4853 8128 4917 8132
rect 4933 8188 4997 8192
rect 4933 8132 4937 8188
rect 4937 8132 4993 8188
rect 4993 8132 4997 8188
rect 4933 8128 4997 8132
rect 8434 8188 8498 8192
rect 8434 8132 8438 8188
rect 8438 8132 8494 8188
rect 8494 8132 8498 8188
rect 8434 8128 8498 8132
rect 8514 8188 8578 8192
rect 8514 8132 8518 8188
rect 8518 8132 8574 8188
rect 8574 8132 8578 8188
rect 8514 8128 8578 8132
rect 8594 8188 8658 8192
rect 8594 8132 8598 8188
rect 8598 8132 8654 8188
rect 8654 8132 8658 8188
rect 8594 8128 8658 8132
rect 8674 8188 8738 8192
rect 8674 8132 8678 8188
rect 8678 8132 8734 8188
rect 8734 8132 8738 8188
rect 8674 8128 8738 8132
rect 3924 8120 3988 8124
rect 3924 8064 3938 8120
rect 3938 8064 3988 8120
rect 3924 8060 3988 8064
rect 9996 8120 10060 8124
rect 9996 8064 10010 8120
rect 10010 8064 10060 8120
rect 9996 8060 10060 8064
rect 10732 8120 10796 8124
rect 10732 8064 10782 8120
rect 10782 8064 10796 8120
rect 10732 8060 10796 8064
rect 3740 7924 3804 7988
rect 9628 7924 9692 7988
rect 2822 7644 2886 7648
rect 2822 7588 2826 7644
rect 2826 7588 2882 7644
rect 2882 7588 2886 7644
rect 2822 7584 2886 7588
rect 2902 7644 2966 7648
rect 2902 7588 2906 7644
rect 2906 7588 2962 7644
rect 2962 7588 2966 7644
rect 2902 7584 2966 7588
rect 2982 7644 3046 7648
rect 2982 7588 2986 7644
rect 2986 7588 3042 7644
rect 3042 7588 3046 7644
rect 2982 7584 3046 7588
rect 3062 7644 3126 7648
rect 3062 7588 3066 7644
rect 3066 7588 3122 7644
rect 3122 7588 3126 7644
rect 3062 7584 3126 7588
rect 6564 7644 6628 7648
rect 6564 7588 6568 7644
rect 6568 7588 6624 7644
rect 6624 7588 6628 7644
rect 6564 7584 6628 7588
rect 6644 7644 6708 7648
rect 6644 7588 6648 7644
rect 6648 7588 6704 7644
rect 6704 7588 6708 7644
rect 6644 7584 6708 7588
rect 6724 7644 6788 7648
rect 6724 7588 6728 7644
rect 6728 7588 6784 7644
rect 6784 7588 6788 7644
rect 6724 7584 6788 7588
rect 6804 7644 6868 7648
rect 6804 7588 6808 7644
rect 6808 7588 6864 7644
rect 6864 7588 6868 7644
rect 6804 7584 6868 7588
rect 10305 7644 10369 7648
rect 10305 7588 10309 7644
rect 10309 7588 10365 7644
rect 10365 7588 10369 7644
rect 10305 7584 10369 7588
rect 10385 7644 10449 7648
rect 10385 7588 10389 7644
rect 10389 7588 10445 7644
rect 10445 7588 10449 7644
rect 10385 7584 10449 7588
rect 10465 7644 10529 7648
rect 10465 7588 10469 7644
rect 10469 7588 10525 7644
rect 10525 7588 10529 7644
rect 10465 7584 10529 7588
rect 10545 7644 10609 7648
rect 10545 7588 10549 7644
rect 10549 7588 10605 7644
rect 10605 7588 10609 7644
rect 10545 7584 10609 7588
rect 5948 7516 6012 7580
rect 4693 7100 4757 7104
rect 4693 7044 4697 7100
rect 4697 7044 4753 7100
rect 4753 7044 4757 7100
rect 4693 7040 4757 7044
rect 4773 7100 4837 7104
rect 4773 7044 4777 7100
rect 4777 7044 4833 7100
rect 4833 7044 4837 7100
rect 4773 7040 4837 7044
rect 4853 7100 4917 7104
rect 4853 7044 4857 7100
rect 4857 7044 4913 7100
rect 4913 7044 4917 7100
rect 4853 7040 4917 7044
rect 4933 7100 4997 7104
rect 4933 7044 4937 7100
rect 4937 7044 4993 7100
rect 4993 7044 4997 7100
rect 4933 7040 4997 7044
rect 8434 7100 8498 7104
rect 8434 7044 8438 7100
rect 8438 7044 8494 7100
rect 8494 7044 8498 7100
rect 8434 7040 8498 7044
rect 8514 7100 8578 7104
rect 8514 7044 8518 7100
rect 8518 7044 8574 7100
rect 8574 7044 8578 7100
rect 8514 7040 8578 7044
rect 8594 7100 8658 7104
rect 8594 7044 8598 7100
rect 8598 7044 8654 7100
rect 8654 7044 8658 7100
rect 8594 7040 8658 7044
rect 8674 7100 8738 7104
rect 8674 7044 8678 7100
rect 8678 7044 8734 7100
rect 8734 7044 8738 7100
rect 8674 7040 8738 7044
rect 2452 6836 2516 6900
rect 2636 6700 2700 6764
rect 7420 6700 7484 6764
rect 5212 6564 5276 6628
rect 2822 6556 2886 6560
rect 2822 6500 2826 6556
rect 2826 6500 2882 6556
rect 2882 6500 2886 6556
rect 2822 6496 2886 6500
rect 2902 6556 2966 6560
rect 2902 6500 2906 6556
rect 2906 6500 2962 6556
rect 2962 6500 2966 6556
rect 2902 6496 2966 6500
rect 2982 6556 3046 6560
rect 2982 6500 2986 6556
rect 2986 6500 3042 6556
rect 3042 6500 3046 6556
rect 2982 6496 3046 6500
rect 3062 6556 3126 6560
rect 3062 6500 3066 6556
rect 3066 6500 3122 6556
rect 3122 6500 3126 6556
rect 3062 6496 3126 6500
rect 6564 6556 6628 6560
rect 6564 6500 6568 6556
rect 6568 6500 6624 6556
rect 6624 6500 6628 6556
rect 6564 6496 6628 6500
rect 6644 6556 6708 6560
rect 6644 6500 6648 6556
rect 6648 6500 6704 6556
rect 6704 6500 6708 6556
rect 6644 6496 6708 6500
rect 6724 6556 6788 6560
rect 6724 6500 6728 6556
rect 6728 6500 6784 6556
rect 6784 6500 6788 6556
rect 6724 6496 6788 6500
rect 6804 6556 6868 6560
rect 6804 6500 6808 6556
rect 6808 6500 6864 6556
rect 6864 6500 6868 6556
rect 6804 6496 6868 6500
rect 10305 6556 10369 6560
rect 10305 6500 10309 6556
rect 10309 6500 10365 6556
rect 10365 6500 10369 6556
rect 10305 6496 10369 6500
rect 10385 6556 10449 6560
rect 10385 6500 10389 6556
rect 10389 6500 10445 6556
rect 10445 6500 10449 6556
rect 10385 6496 10449 6500
rect 10465 6556 10529 6560
rect 10465 6500 10469 6556
rect 10469 6500 10525 6556
rect 10525 6500 10529 6556
rect 10465 6496 10529 6500
rect 10545 6556 10609 6560
rect 10545 6500 10549 6556
rect 10549 6500 10605 6556
rect 10605 6500 10609 6556
rect 10545 6496 10609 6500
rect 5580 6428 5644 6492
rect 5580 6292 5644 6356
rect 6316 6156 6380 6220
rect 4108 6020 4172 6084
rect 4693 6012 4757 6016
rect 4693 5956 4697 6012
rect 4697 5956 4753 6012
rect 4753 5956 4757 6012
rect 4693 5952 4757 5956
rect 4773 6012 4837 6016
rect 4773 5956 4777 6012
rect 4777 5956 4833 6012
rect 4833 5956 4837 6012
rect 4773 5952 4837 5956
rect 4853 6012 4917 6016
rect 4853 5956 4857 6012
rect 4857 5956 4913 6012
rect 4913 5956 4917 6012
rect 4853 5952 4917 5956
rect 4933 6012 4997 6016
rect 4933 5956 4937 6012
rect 4937 5956 4993 6012
rect 4993 5956 4997 6012
rect 4933 5952 4997 5956
rect 8434 6012 8498 6016
rect 8434 5956 8438 6012
rect 8438 5956 8494 6012
rect 8494 5956 8498 6012
rect 8434 5952 8498 5956
rect 8514 6012 8578 6016
rect 8514 5956 8518 6012
rect 8518 5956 8574 6012
rect 8574 5956 8578 6012
rect 8514 5952 8578 5956
rect 8594 6012 8658 6016
rect 8594 5956 8598 6012
rect 8598 5956 8654 6012
rect 8654 5956 8658 6012
rect 8594 5952 8658 5956
rect 8674 6012 8738 6016
rect 8674 5956 8678 6012
rect 8678 5956 8734 6012
rect 8734 5956 8738 6012
rect 8674 5952 8738 5956
rect 4108 5884 4172 5948
rect 1532 5612 1596 5676
rect 2822 5468 2886 5472
rect 2822 5412 2826 5468
rect 2826 5412 2882 5468
rect 2882 5412 2886 5468
rect 2822 5408 2886 5412
rect 2902 5468 2966 5472
rect 2902 5412 2906 5468
rect 2906 5412 2962 5468
rect 2962 5412 2966 5468
rect 2902 5408 2966 5412
rect 2982 5468 3046 5472
rect 2982 5412 2986 5468
rect 2986 5412 3042 5468
rect 3042 5412 3046 5468
rect 2982 5408 3046 5412
rect 3062 5468 3126 5472
rect 3062 5412 3066 5468
rect 3066 5412 3122 5468
rect 3122 5412 3126 5468
rect 3062 5408 3126 5412
rect 6564 5468 6628 5472
rect 6564 5412 6568 5468
rect 6568 5412 6624 5468
rect 6624 5412 6628 5468
rect 6564 5408 6628 5412
rect 6644 5468 6708 5472
rect 6644 5412 6648 5468
rect 6648 5412 6704 5468
rect 6704 5412 6708 5468
rect 6644 5408 6708 5412
rect 6724 5468 6788 5472
rect 6724 5412 6728 5468
rect 6728 5412 6784 5468
rect 6784 5412 6788 5468
rect 6724 5408 6788 5412
rect 6804 5468 6868 5472
rect 6804 5412 6808 5468
rect 6808 5412 6864 5468
rect 6864 5412 6868 5468
rect 6804 5408 6868 5412
rect 10305 5468 10369 5472
rect 10305 5412 10309 5468
rect 10309 5412 10365 5468
rect 10365 5412 10369 5468
rect 10305 5408 10369 5412
rect 10385 5468 10449 5472
rect 10385 5412 10389 5468
rect 10389 5412 10445 5468
rect 10445 5412 10449 5468
rect 10385 5408 10449 5412
rect 10465 5468 10529 5472
rect 10465 5412 10469 5468
rect 10469 5412 10525 5468
rect 10525 5412 10529 5468
rect 10465 5408 10529 5412
rect 10545 5468 10609 5472
rect 10545 5412 10549 5468
rect 10549 5412 10605 5468
rect 10605 5412 10609 5468
rect 10545 5408 10609 5412
rect 8156 5204 8220 5268
rect 2452 4796 2516 4860
rect 6132 5068 6196 5132
rect 7972 4932 8036 4996
rect 10732 4932 10796 4996
rect 4693 4924 4757 4928
rect 4693 4868 4697 4924
rect 4697 4868 4753 4924
rect 4753 4868 4757 4924
rect 4693 4864 4757 4868
rect 4773 4924 4837 4928
rect 4773 4868 4777 4924
rect 4777 4868 4833 4924
rect 4833 4868 4837 4924
rect 4773 4864 4837 4868
rect 4853 4924 4917 4928
rect 4853 4868 4857 4924
rect 4857 4868 4913 4924
rect 4913 4868 4917 4924
rect 4853 4864 4917 4868
rect 4933 4924 4997 4928
rect 4933 4868 4937 4924
rect 4937 4868 4993 4924
rect 4993 4868 4997 4924
rect 4933 4864 4997 4868
rect 8434 4924 8498 4928
rect 8434 4868 8438 4924
rect 8438 4868 8494 4924
rect 8494 4868 8498 4924
rect 8434 4864 8498 4868
rect 8514 4924 8578 4928
rect 8514 4868 8518 4924
rect 8518 4868 8574 4924
rect 8574 4868 8578 4924
rect 8514 4864 8578 4868
rect 8594 4924 8658 4928
rect 8594 4868 8598 4924
rect 8598 4868 8654 4924
rect 8654 4868 8658 4924
rect 8594 4864 8658 4868
rect 8674 4924 8738 4928
rect 8674 4868 8678 4924
rect 8678 4868 8734 4924
rect 8734 4868 8738 4924
rect 8674 4864 8738 4868
rect 4476 4660 4540 4724
rect 2452 4524 2516 4588
rect 2822 4380 2886 4384
rect 2822 4324 2826 4380
rect 2826 4324 2882 4380
rect 2882 4324 2886 4380
rect 2822 4320 2886 4324
rect 2902 4380 2966 4384
rect 2902 4324 2906 4380
rect 2906 4324 2962 4380
rect 2962 4324 2966 4380
rect 2902 4320 2966 4324
rect 2982 4380 3046 4384
rect 2982 4324 2986 4380
rect 2986 4324 3042 4380
rect 3042 4324 3046 4380
rect 2982 4320 3046 4324
rect 3062 4380 3126 4384
rect 3062 4324 3066 4380
rect 3066 4324 3122 4380
rect 3122 4324 3126 4380
rect 3062 4320 3126 4324
rect 1164 3980 1228 4044
rect 4476 3844 4540 3908
rect 4693 3836 4757 3840
rect 4693 3780 4697 3836
rect 4697 3780 4753 3836
rect 4753 3780 4757 3836
rect 4693 3776 4757 3780
rect 4773 3836 4837 3840
rect 4773 3780 4777 3836
rect 4777 3780 4833 3836
rect 4833 3780 4837 3836
rect 4773 3776 4837 3780
rect 4853 3836 4917 3840
rect 4853 3780 4857 3836
rect 4857 3780 4913 3836
rect 4913 3780 4917 3836
rect 4853 3776 4917 3780
rect 4933 3836 4997 3840
rect 4933 3780 4937 3836
rect 4937 3780 4993 3836
rect 4993 3780 4997 3836
rect 4933 3776 4997 3780
rect 2268 3496 2332 3500
rect 2268 3440 2318 3496
rect 2318 3440 2332 3496
rect 2268 3436 2332 3440
rect 5396 3436 5460 3500
rect 2822 3292 2886 3296
rect 2822 3236 2826 3292
rect 2826 3236 2882 3292
rect 2882 3236 2886 3292
rect 2822 3232 2886 3236
rect 2902 3292 2966 3296
rect 2902 3236 2906 3292
rect 2906 3236 2962 3292
rect 2962 3236 2966 3292
rect 2902 3232 2966 3236
rect 2982 3292 3046 3296
rect 2982 3236 2986 3292
rect 2986 3236 3042 3292
rect 3042 3236 3046 3292
rect 2982 3232 3046 3236
rect 3062 3292 3126 3296
rect 3062 3236 3066 3292
rect 3066 3236 3122 3292
rect 3122 3236 3126 3292
rect 3062 3232 3126 3236
rect 5396 3164 5460 3228
rect 3740 3028 3804 3092
rect 4476 3028 4540 3092
rect 9076 4524 9140 4588
rect 6564 4380 6628 4384
rect 6564 4324 6568 4380
rect 6568 4324 6624 4380
rect 6624 4324 6628 4380
rect 6564 4320 6628 4324
rect 6644 4380 6708 4384
rect 6644 4324 6648 4380
rect 6648 4324 6704 4380
rect 6704 4324 6708 4380
rect 6644 4320 6708 4324
rect 6724 4380 6788 4384
rect 6724 4324 6728 4380
rect 6728 4324 6784 4380
rect 6784 4324 6788 4380
rect 6724 4320 6788 4324
rect 6804 4380 6868 4384
rect 6804 4324 6808 4380
rect 6808 4324 6864 4380
rect 6864 4324 6868 4380
rect 6804 4320 6868 4324
rect 10305 4380 10369 4384
rect 10305 4324 10309 4380
rect 10309 4324 10365 4380
rect 10365 4324 10369 4380
rect 10305 4320 10369 4324
rect 10385 4380 10449 4384
rect 10385 4324 10389 4380
rect 10389 4324 10445 4380
rect 10445 4324 10449 4380
rect 10385 4320 10449 4324
rect 10465 4380 10529 4384
rect 10465 4324 10469 4380
rect 10469 4324 10525 4380
rect 10525 4324 10529 4380
rect 10465 4320 10529 4324
rect 10545 4380 10609 4384
rect 10545 4324 10549 4380
rect 10549 4324 10605 4380
rect 10605 4324 10609 4380
rect 10545 4320 10609 4324
rect 8434 3836 8498 3840
rect 8434 3780 8438 3836
rect 8438 3780 8494 3836
rect 8494 3780 8498 3836
rect 8434 3776 8498 3780
rect 8514 3836 8578 3840
rect 8514 3780 8518 3836
rect 8518 3780 8574 3836
rect 8574 3780 8578 3836
rect 8514 3776 8578 3780
rect 8594 3836 8658 3840
rect 8594 3780 8598 3836
rect 8598 3780 8654 3836
rect 8654 3780 8658 3836
rect 8594 3776 8658 3780
rect 8674 3836 8738 3840
rect 8674 3780 8678 3836
rect 8678 3780 8734 3836
rect 8734 3780 8738 3836
rect 8674 3776 8738 3780
rect 9812 3708 9876 3772
rect 9628 3300 9692 3364
rect 6564 3292 6628 3296
rect 6564 3236 6568 3292
rect 6568 3236 6624 3292
rect 6624 3236 6628 3292
rect 6564 3232 6628 3236
rect 6644 3292 6708 3296
rect 6644 3236 6648 3292
rect 6648 3236 6704 3292
rect 6704 3236 6708 3292
rect 6644 3232 6708 3236
rect 6724 3292 6788 3296
rect 6724 3236 6728 3292
rect 6728 3236 6784 3292
rect 6784 3236 6788 3292
rect 6724 3232 6788 3236
rect 6804 3292 6868 3296
rect 6804 3236 6808 3292
rect 6808 3236 6864 3292
rect 6864 3236 6868 3292
rect 6804 3232 6868 3236
rect 10305 3292 10369 3296
rect 10305 3236 10309 3292
rect 10309 3236 10365 3292
rect 10365 3236 10369 3292
rect 10305 3232 10369 3236
rect 10385 3292 10449 3296
rect 10385 3236 10389 3292
rect 10389 3236 10445 3292
rect 10445 3236 10449 3292
rect 10385 3232 10449 3236
rect 10465 3292 10529 3296
rect 10465 3236 10469 3292
rect 10469 3236 10525 3292
rect 10525 3236 10529 3292
rect 10465 3232 10529 3236
rect 10545 3292 10609 3296
rect 10545 3236 10549 3292
rect 10549 3236 10605 3292
rect 10605 3236 10609 3292
rect 10545 3232 10609 3236
rect 2452 2892 2516 2956
rect 4292 2892 4356 2956
rect 5212 2952 5276 2956
rect 5212 2896 5262 2952
rect 5262 2896 5276 2952
rect 5212 2892 5276 2896
rect 8156 2892 8220 2956
rect 4693 2748 4757 2752
rect 4693 2692 4697 2748
rect 4697 2692 4753 2748
rect 4753 2692 4757 2748
rect 4693 2688 4757 2692
rect 4773 2748 4837 2752
rect 4773 2692 4777 2748
rect 4777 2692 4833 2748
rect 4833 2692 4837 2748
rect 4773 2688 4837 2692
rect 4853 2748 4917 2752
rect 4853 2692 4857 2748
rect 4857 2692 4913 2748
rect 4913 2692 4917 2748
rect 4853 2688 4917 2692
rect 4933 2748 4997 2752
rect 4933 2692 4937 2748
rect 4937 2692 4993 2748
rect 4993 2692 4997 2748
rect 4933 2688 4997 2692
rect 3372 2544 3436 2548
rect 3372 2488 3386 2544
rect 3386 2488 3436 2544
rect 3372 2484 3436 2488
rect 7052 2756 7116 2820
rect 9076 2892 9140 2956
rect 9996 2892 10060 2956
rect 8434 2748 8498 2752
rect 8434 2692 8438 2748
rect 8438 2692 8494 2748
rect 8494 2692 8498 2748
rect 8434 2688 8498 2692
rect 8514 2748 8578 2752
rect 8514 2692 8518 2748
rect 8518 2692 8574 2748
rect 8574 2692 8578 2748
rect 8514 2688 8578 2692
rect 8594 2748 8658 2752
rect 8594 2692 8598 2748
rect 8598 2692 8654 2748
rect 8654 2692 8658 2748
rect 8594 2688 8658 2692
rect 8674 2748 8738 2752
rect 8674 2692 8678 2748
rect 8678 2692 8734 2748
rect 8734 2692 8738 2748
rect 8674 2688 8738 2692
rect 5580 2544 5644 2548
rect 5580 2488 5630 2544
rect 5630 2488 5644 2544
rect 5580 2484 5644 2488
rect 8892 2484 8956 2548
rect 5396 2348 5460 2412
rect 7972 2348 8036 2412
rect 5764 2212 5828 2276
rect 7420 2212 7484 2276
rect 2822 2204 2886 2208
rect 2822 2148 2826 2204
rect 2826 2148 2882 2204
rect 2882 2148 2886 2204
rect 2822 2144 2886 2148
rect 2902 2204 2966 2208
rect 2902 2148 2906 2204
rect 2906 2148 2962 2204
rect 2962 2148 2966 2204
rect 2902 2144 2966 2148
rect 2982 2204 3046 2208
rect 2982 2148 2986 2204
rect 2986 2148 3042 2204
rect 3042 2148 3046 2204
rect 2982 2144 3046 2148
rect 3062 2204 3126 2208
rect 3062 2148 3066 2204
rect 3066 2148 3122 2204
rect 3122 2148 3126 2204
rect 3062 2144 3126 2148
rect 6564 2204 6628 2208
rect 6564 2148 6568 2204
rect 6568 2148 6624 2204
rect 6624 2148 6628 2204
rect 6564 2144 6628 2148
rect 6644 2204 6708 2208
rect 6644 2148 6648 2204
rect 6648 2148 6704 2204
rect 6704 2148 6708 2204
rect 6644 2144 6708 2148
rect 6724 2204 6788 2208
rect 6724 2148 6728 2204
rect 6728 2148 6784 2204
rect 6784 2148 6788 2204
rect 6724 2144 6788 2148
rect 6804 2204 6868 2208
rect 6804 2148 6808 2204
rect 6808 2148 6864 2204
rect 6864 2148 6868 2204
rect 6804 2144 6868 2148
rect 10305 2204 10369 2208
rect 10305 2148 10309 2204
rect 10309 2148 10365 2204
rect 10365 2148 10369 2204
rect 10305 2144 10369 2148
rect 10385 2204 10449 2208
rect 10385 2148 10389 2204
rect 10389 2148 10445 2204
rect 10445 2148 10449 2204
rect 10385 2144 10449 2148
rect 10465 2204 10529 2208
rect 10465 2148 10469 2204
rect 10469 2148 10525 2204
rect 10525 2148 10529 2204
rect 10465 2144 10529 2148
rect 10545 2204 10609 2208
rect 10545 2148 10549 2204
rect 10549 2148 10605 2204
rect 10605 2148 10609 2204
rect 10545 2144 10609 2148
rect 5948 1940 6012 2004
rect 4108 1804 4172 1868
rect 7604 1668 7668 1732
rect 2636 1532 2700 1596
rect 6316 1532 6380 1596
rect 7236 1396 7300 1460
rect 6132 1260 6196 1324
rect 3556 1124 3620 1188
rect 9812 1124 9876 1188
rect 7788 988 7852 1052
rect 3924 852 3988 916
<< metal4 >>
rect 2814 13088 3135 13104
rect 2814 13024 2822 13088
rect 2886 13024 2902 13088
rect 2966 13024 2982 13088
rect 3046 13024 3062 13088
rect 3126 13024 3135 13088
rect 1163 12884 1229 12885
rect 1163 12820 1164 12884
rect 1228 12820 1229 12884
rect 1163 12819 1229 12820
rect 1166 4045 1226 12819
rect 2814 12000 3135 13024
rect 2814 11936 2822 12000
rect 2886 11936 2902 12000
rect 2966 11936 2982 12000
rect 3046 11936 3062 12000
rect 3126 11936 3135 12000
rect 2814 10912 3135 11936
rect 2814 10848 2822 10912
rect 2886 10848 2902 10912
rect 2966 10848 2982 10912
rect 3046 10848 3062 10912
rect 3126 10848 3135 10912
rect 2814 9824 3135 10848
rect 4685 12544 5005 13104
rect 4685 12480 4693 12544
rect 4757 12480 4773 12544
rect 4837 12480 4853 12544
rect 4917 12480 4933 12544
rect 4997 12480 5005 12544
rect 4685 11456 5005 12480
rect 4685 11392 4693 11456
rect 4757 11392 4773 11456
rect 4837 11392 4853 11456
rect 4917 11392 4933 11456
rect 4997 11392 5005 11456
rect 4107 10844 4173 10845
rect 4107 10780 4108 10844
rect 4172 10780 4173 10844
rect 4107 10779 4173 10780
rect 3555 9892 3621 9893
rect 3555 9828 3556 9892
rect 3620 9828 3621 9892
rect 3555 9827 3621 9828
rect 2814 9760 2822 9824
rect 2886 9760 2902 9824
rect 2966 9760 2982 9824
rect 3046 9760 3062 9824
rect 3126 9760 3135 9824
rect 1531 9212 1597 9213
rect 1531 9148 1532 9212
rect 1596 9148 1597 9212
rect 1531 9147 1597 9148
rect 1534 5677 1594 9147
rect 2814 8736 3135 9760
rect 3371 9484 3437 9485
rect 3371 9420 3372 9484
rect 3436 9420 3437 9484
rect 3371 9419 3437 9420
rect 2814 8672 2822 8736
rect 2886 8672 2902 8736
rect 2966 8672 2982 8736
rect 3046 8672 3062 8736
rect 3126 8672 3135 8736
rect 2267 8532 2333 8533
rect 2267 8468 2268 8532
rect 2332 8468 2333 8532
rect 2267 8467 2333 8468
rect 1531 5676 1597 5677
rect 1531 5612 1532 5676
rect 1596 5612 1597 5676
rect 1531 5611 1597 5612
rect 1163 4044 1229 4045
rect 1163 3980 1164 4044
rect 1228 3980 1229 4044
rect 1163 3979 1229 3980
rect 2270 3501 2330 8467
rect 2814 7648 3135 8672
rect 2814 7584 2822 7648
rect 2886 7584 2902 7648
rect 2966 7584 2982 7648
rect 3046 7584 3062 7648
rect 3126 7584 3135 7648
rect 2451 6900 2517 6901
rect 2451 6836 2452 6900
rect 2516 6836 2517 6900
rect 2451 6835 2517 6836
rect 2454 4861 2514 6835
rect 2635 6764 2701 6765
rect 2635 6700 2636 6764
rect 2700 6700 2701 6764
rect 2635 6699 2701 6700
rect 2451 4860 2517 4861
rect 2451 4796 2452 4860
rect 2516 4796 2517 4860
rect 2451 4795 2517 4796
rect 2451 4588 2517 4589
rect 2451 4524 2452 4588
rect 2516 4524 2517 4588
rect 2451 4523 2517 4524
rect 2267 3500 2333 3501
rect 2267 3436 2268 3500
rect 2332 3436 2333 3500
rect 2267 3435 2333 3436
rect 2454 2957 2514 4523
rect 2451 2956 2517 2957
rect 2451 2892 2452 2956
rect 2516 2892 2517 2956
rect 2451 2891 2517 2892
rect 2638 1597 2698 6699
rect 2814 6560 3135 7584
rect 2814 6496 2822 6560
rect 2886 6496 2902 6560
rect 2966 6496 2982 6560
rect 3046 6496 3062 6560
rect 3126 6496 3135 6560
rect 2814 5472 3135 6496
rect 2814 5408 2822 5472
rect 2886 5408 2902 5472
rect 2966 5408 2982 5472
rect 3046 5408 3062 5472
rect 3126 5408 3135 5472
rect 2814 4384 3135 5408
rect 2814 4320 2822 4384
rect 2886 4320 2902 4384
rect 2966 4320 2982 4384
rect 3046 4320 3062 4384
rect 3126 4320 3135 4384
rect 2814 3296 3135 4320
rect 2814 3232 2822 3296
rect 2886 3232 2902 3296
rect 2966 3232 2982 3296
rect 3046 3232 3062 3296
rect 3126 3232 3135 3296
rect 2814 2208 3135 3232
rect 3374 2549 3434 9419
rect 3371 2548 3437 2549
rect 3371 2484 3372 2548
rect 3436 2484 3437 2548
rect 3371 2483 3437 2484
rect 2814 2144 2822 2208
rect 2886 2144 2902 2208
rect 2966 2144 2982 2208
rect 3046 2144 3062 2208
rect 3126 2144 3135 2208
rect 2814 2128 3135 2144
rect 2635 1596 2701 1597
rect 2635 1532 2636 1596
rect 2700 1532 2701 1596
rect 2635 1531 2701 1532
rect 3558 1189 3618 9827
rect 3923 8124 3989 8125
rect 3923 8060 3924 8124
rect 3988 8060 3989 8124
rect 3923 8059 3989 8060
rect 3739 7988 3805 7989
rect 3739 7924 3740 7988
rect 3804 7924 3805 7988
rect 3739 7923 3805 7924
rect 3742 3093 3802 7923
rect 3739 3092 3805 3093
rect 3739 3028 3740 3092
rect 3804 3028 3805 3092
rect 3739 3027 3805 3028
rect 3555 1188 3621 1189
rect 3555 1124 3556 1188
rect 3620 1124 3621 1188
rect 3555 1123 3621 1124
rect 3926 917 3986 8059
rect 4110 6085 4170 10779
rect 4475 10708 4541 10709
rect 4475 10644 4476 10708
rect 4540 10644 4541 10708
rect 4475 10643 4541 10644
rect 4291 10572 4357 10573
rect 4291 10508 4292 10572
rect 4356 10508 4357 10572
rect 4291 10507 4357 10508
rect 4107 6084 4173 6085
rect 4107 6020 4108 6084
rect 4172 6020 4173 6084
rect 4107 6019 4173 6020
rect 4107 5948 4173 5949
rect 4107 5884 4108 5948
rect 4172 5884 4173 5948
rect 4107 5883 4173 5884
rect 4110 1869 4170 5883
rect 4294 2957 4354 10507
rect 4478 4725 4538 10643
rect 4685 10368 5005 11392
rect 6556 13088 6876 13104
rect 6556 13024 6564 13088
rect 6628 13024 6644 13088
rect 6708 13024 6724 13088
rect 6788 13024 6804 13088
rect 6868 13024 6876 13088
rect 6556 12000 6876 13024
rect 6556 11936 6564 12000
rect 6628 11936 6644 12000
rect 6708 11936 6724 12000
rect 6788 11936 6804 12000
rect 6868 11936 6876 12000
rect 5763 11116 5829 11117
rect 5763 11052 5764 11116
rect 5828 11052 5829 11116
rect 5763 11051 5829 11052
rect 4685 10304 4693 10368
rect 4757 10304 4773 10368
rect 4837 10304 4853 10368
rect 4917 10304 4933 10368
rect 4997 10304 5005 10368
rect 4685 9280 5005 10304
rect 4685 9216 4693 9280
rect 4757 9216 4773 9280
rect 4837 9216 4853 9280
rect 4917 9216 4933 9280
rect 4997 9216 5005 9280
rect 4685 8192 5005 9216
rect 5395 9212 5461 9213
rect 5395 9148 5396 9212
rect 5460 9148 5461 9212
rect 5395 9147 5461 9148
rect 4685 8128 4693 8192
rect 4757 8128 4773 8192
rect 4837 8128 4853 8192
rect 4917 8128 4933 8192
rect 4997 8128 5005 8192
rect 4685 7104 5005 8128
rect 4685 7040 4693 7104
rect 4757 7040 4773 7104
rect 4837 7040 4853 7104
rect 4917 7040 4933 7104
rect 4997 7040 5005 7104
rect 4685 6016 5005 7040
rect 5211 6628 5277 6629
rect 5211 6564 5212 6628
rect 5276 6564 5277 6628
rect 5211 6563 5277 6564
rect 4685 5952 4693 6016
rect 4757 5952 4773 6016
rect 4837 5952 4853 6016
rect 4917 5952 4933 6016
rect 4997 5952 5005 6016
rect 4685 4928 5005 5952
rect 4685 4864 4693 4928
rect 4757 4864 4773 4928
rect 4837 4864 4853 4928
rect 4917 4864 4933 4928
rect 4997 4864 5005 4928
rect 4475 4724 4541 4725
rect 4475 4660 4476 4724
rect 4540 4660 4541 4724
rect 4475 4659 4541 4660
rect 4475 3908 4541 3909
rect 4475 3844 4476 3908
rect 4540 3844 4541 3908
rect 4475 3843 4541 3844
rect 4478 3093 4538 3843
rect 4685 3840 5005 4864
rect 4685 3776 4693 3840
rect 4757 3776 4773 3840
rect 4837 3776 4853 3840
rect 4917 3776 4933 3840
rect 4997 3776 5005 3840
rect 4475 3092 4541 3093
rect 4475 3028 4476 3092
rect 4540 3028 4541 3092
rect 4475 3027 4541 3028
rect 4291 2956 4357 2957
rect 4291 2892 4292 2956
rect 4356 2892 4357 2956
rect 4291 2891 4357 2892
rect 4685 2752 5005 3776
rect 5214 2957 5274 6563
rect 5398 3501 5458 9147
rect 5579 8396 5645 8397
rect 5579 8332 5580 8396
rect 5644 8332 5645 8396
rect 5579 8331 5645 8332
rect 5582 6493 5642 8331
rect 5579 6492 5645 6493
rect 5579 6428 5580 6492
rect 5644 6428 5645 6492
rect 5579 6427 5645 6428
rect 5579 6356 5645 6357
rect 5579 6292 5580 6356
rect 5644 6292 5645 6356
rect 5579 6291 5645 6292
rect 5395 3500 5461 3501
rect 5395 3436 5396 3500
rect 5460 3436 5461 3500
rect 5395 3435 5461 3436
rect 5395 3228 5461 3229
rect 5395 3164 5396 3228
rect 5460 3164 5461 3228
rect 5395 3163 5461 3164
rect 5211 2956 5277 2957
rect 5211 2892 5212 2956
rect 5276 2892 5277 2956
rect 5211 2891 5277 2892
rect 4685 2688 4693 2752
rect 4757 2688 4773 2752
rect 4837 2688 4853 2752
rect 4917 2688 4933 2752
rect 4997 2688 5005 2752
rect 4685 2128 5005 2688
rect 5398 2413 5458 3163
rect 5582 2549 5642 6291
rect 5579 2548 5645 2549
rect 5579 2484 5580 2548
rect 5644 2484 5645 2548
rect 5579 2483 5645 2484
rect 5395 2412 5461 2413
rect 5395 2348 5396 2412
rect 5460 2348 5461 2412
rect 5395 2347 5461 2348
rect 5766 2277 5826 11051
rect 6556 10912 6876 11936
rect 8426 12544 8747 13104
rect 8426 12480 8434 12544
rect 8498 12480 8514 12544
rect 8578 12480 8594 12544
rect 8658 12480 8674 12544
rect 8738 12480 8747 12544
rect 8426 11456 8747 12480
rect 8426 11392 8434 11456
rect 8498 11392 8514 11456
rect 8578 11392 8594 11456
rect 8658 11392 8674 11456
rect 8738 11392 8747 11456
rect 7235 11252 7301 11253
rect 7235 11188 7236 11252
rect 7300 11188 7301 11252
rect 7235 11187 7301 11188
rect 7603 11252 7669 11253
rect 7603 11188 7604 11252
rect 7668 11188 7669 11252
rect 7603 11187 7669 11188
rect 6556 10848 6564 10912
rect 6628 10848 6644 10912
rect 6708 10848 6724 10912
rect 6788 10848 6804 10912
rect 6868 10848 6876 10912
rect 6556 9824 6876 10848
rect 7051 10164 7117 10165
rect 7051 10100 7052 10164
rect 7116 10100 7117 10164
rect 7051 10099 7117 10100
rect 6556 9760 6564 9824
rect 6628 9760 6644 9824
rect 6708 9760 6724 9824
rect 6788 9760 6804 9824
rect 6868 9760 6876 9824
rect 6556 8736 6876 9760
rect 6556 8672 6564 8736
rect 6628 8672 6644 8736
rect 6708 8672 6724 8736
rect 6788 8672 6804 8736
rect 6868 8672 6876 8736
rect 6556 7648 6876 8672
rect 6556 7584 6564 7648
rect 6628 7584 6644 7648
rect 6708 7584 6724 7648
rect 6788 7584 6804 7648
rect 6868 7584 6876 7648
rect 5947 7580 6013 7581
rect 5947 7516 5948 7580
rect 6012 7516 6013 7580
rect 5947 7515 6013 7516
rect 5763 2276 5829 2277
rect 5763 2212 5764 2276
rect 5828 2212 5829 2276
rect 5763 2211 5829 2212
rect 5950 2005 6010 7515
rect 6556 6560 6876 7584
rect 6556 6496 6564 6560
rect 6628 6496 6644 6560
rect 6708 6496 6724 6560
rect 6788 6496 6804 6560
rect 6868 6496 6876 6560
rect 6315 6220 6381 6221
rect 6315 6156 6316 6220
rect 6380 6156 6381 6220
rect 6315 6155 6381 6156
rect 6131 5132 6197 5133
rect 6131 5068 6132 5132
rect 6196 5068 6197 5132
rect 6131 5067 6197 5068
rect 5947 2004 6013 2005
rect 5947 1940 5948 2004
rect 6012 1940 6013 2004
rect 5947 1939 6013 1940
rect 4107 1868 4173 1869
rect 4107 1804 4108 1868
rect 4172 1804 4173 1868
rect 4107 1803 4173 1804
rect 6134 1325 6194 5067
rect 6318 1597 6378 6155
rect 6556 5472 6876 6496
rect 6556 5408 6564 5472
rect 6628 5408 6644 5472
rect 6708 5408 6724 5472
rect 6788 5408 6804 5472
rect 6868 5408 6876 5472
rect 6556 4384 6876 5408
rect 6556 4320 6564 4384
rect 6628 4320 6644 4384
rect 6708 4320 6724 4384
rect 6788 4320 6804 4384
rect 6868 4320 6876 4384
rect 6556 3296 6876 4320
rect 6556 3232 6564 3296
rect 6628 3232 6644 3296
rect 6708 3232 6724 3296
rect 6788 3232 6804 3296
rect 6868 3232 6876 3296
rect 6556 2208 6876 3232
rect 7054 2821 7114 10099
rect 7051 2820 7117 2821
rect 7051 2756 7052 2820
rect 7116 2756 7117 2820
rect 7051 2755 7117 2756
rect 6556 2144 6564 2208
rect 6628 2144 6644 2208
rect 6708 2144 6724 2208
rect 6788 2144 6804 2208
rect 6868 2144 6876 2208
rect 6556 2128 6876 2144
rect 6315 1596 6381 1597
rect 6315 1532 6316 1596
rect 6380 1532 6381 1596
rect 6315 1531 6381 1532
rect 7238 1461 7298 11187
rect 7419 6764 7485 6765
rect 7419 6700 7420 6764
rect 7484 6700 7485 6764
rect 7419 6699 7485 6700
rect 7422 2277 7482 6699
rect 7419 2276 7485 2277
rect 7419 2212 7420 2276
rect 7484 2212 7485 2276
rect 7419 2211 7485 2212
rect 7606 1733 7666 11187
rect 7787 11116 7853 11117
rect 7787 11052 7788 11116
rect 7852 11052 7853 11116
rect 7787 11051 7853 11052
rect 7603 1732 7669 1733
rect 7603 1668 7604 1732
rect 7668 1668 7669 1732
rect 7603 1667 7669 1668
rect 7235 1460 7301 1461
rect 7235 1396 7236 1460
rect 7300 1396 7301 1460
rect 7235 1395 7301 1396
rect 6131 1324 6197 1325
rect 6131 1260 6132 1324
rect 6196 1260 6197 1324
rect 6131 1259 6197 1260
rect 7790 1053 7850 11051
rect 8155 10572 8221 10573
rect 8155 10508 8156 10572
rect 8220 10508 8221 10572
rect 8155 10507 8221 10508
rect 7971 8940 8037 8941
rect 7971 8876 7972 8940
rect 8036 8876 8037 8940
rect 7971 8875 8037 8876
rect 7974 5130 8034 8875
rect 8158 5269 8218 10507
rect 8426 10368 8747 11392
rect 8426 10304 8434 10368
rect 8498 10304 8514 10368
rect 8578 10304 8594 10368
rect 8658 10304 8674 10368
rect 8738 10304 8747 10368
rect 8426 9280 8747 10304
rect 10297 13088 10617 13104
rect 10297 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10465 13088
rect 10529 13024 10545 13088
rect 10609 13024 10617 13088
rect 10297 12000 10617 13024
rect 10297 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10545 12000
rect 10609 11936 10617 12000
rect 10297 10912 10617 11936
rect 10297 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10545 10912
rect 10609 10848 10617 10912
rect 10297 9824 10617 10848
rect 10297 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10545 9824
rect 10609 9760 10617 9824
rect 8891 9620 8957 9621
rect 8891 9556 8892 9620
rect 8956 9556 8957 9620
rect 8891 9555 8957 9556
rect 8426 9216 8434 9280
rect 8498 9216 8514 9280
rect 8578 9216 8594 9280
rect 8658 9216 8674 9280
rect 8738 9216 8747 9280
rect 8426 8192 8747 9216
rect 8426 8128 8434 8192
rect 8498 8128 8514 8192
rect 8578 8128 8594 8192
rect 8658 8128 8674 8192
rect 8738 8128 8747 8192
rect 8426 7104 8747 8128
rect 8426 7040 8434 7104
rect 8498 7040 8514 7104
rect 8578 7040 8594 7104
rect 8658 7040 8674 7104
rect 8738 7040 8747 7104
rect 8426 6016 8747 7040
rect 8426 5952 8434 6016
rect 8498 5952 8514 6016
rect 8578 5952 8594 6016
rect 8658 5952 8674 6016
rect 8738 5952 8747 6016
rect 8155 5268 8221 5269
rect 8155 5204 8156 5268
rect 8220 5204 8221 5268
rect 8155 5203 8221 5204
rect 7974 5070 8218 5130
rect 7971 4996 8037 4997
rect 7971 4932 7972 4996
rect 8036 4932 8037 4996
rect 7971 4931 8037 4932
rect 7974 2413 8034 4931
rect 8158 2957 8218 5070
rect 8426 4928 8747 5952
rect 8426 4864 8434 4928
rect 8498 4864 8514 4928
rect 8578 4864 8594 4928
rect 8658 4864 8674 4928
rect 8738 4864 8747 4928
rect 8426 3840 8747 4864
rect 8426 3776 8434 3840
rect 8498 3776 8514 3840
rect 8578 3776 8594 3840
rect 8658 3776 8674 3840
rect 8738 3776 8747 3840
rect 8155 2956 8221 2957
rect 8155 2892 8156 2956
rect 8220 2892 8221 2956
rect 8155 2891 8221 2892
rect 8426 2752 8747 3776
rect 8426 2688 8434 2752
rect 8498 2688 8514 2752
rect 8578 2688 8594 2752
rect 8658 2688 8674 2752
rect 8738 2688 8747 2752
rect 7971 2412 8037 2413
rect 7971 2348 7972 2412
rect 8036 2348 8037 2412
rect 7971 2347 8037 2348
rect 8426 2128 8747 2688
rect 8894 2549 8954 9555
rect 10297 8736 10617 9760
rect 10297 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10545 8736
rect 10609 8672 10617 8736
rect 9995 8124 10061 8125
rect 9995 8060 9996 8124
rect 10060 8060 10061 8124
rect 9995 8059 10061 8060
rect 9627 7988 9693 7989
rect 9627 7924 9628 7988
rect 9692 7924 9693 7988
rect 9627 7923 9693 7924
rect 9075 4588 9141 4589
rect 9075 4524 9076 4588
rect 9140 4524 9141 4588
rect 9075 4523 9141 4524
rect 9078 2957 9138 4523
rect 9630 3365 9690 7923
rect 9811 3772 9877 3773
rect 9811 3708 9812 3772
rect 9876 3708 9877 3772
rect 9811 3707 9877 3708
rect 9627 3364 9693 3365
rect 9627 3300 9628 3364
rect 9692 3300 9693 3364
rect 9627 3299 9693 3300
rect 9075 2956 9141 2957
rect 9075 2892 9076 2956
rect 9140 2892 9141 2956
rect 9075 2891 9141 2892
rect 8891 2548 8957 2549
rect 8891 2484 8892 2548
rect 8956 2484 8957 2548
rect 8891 2483 8957 2484
rect 9814 1189 9874 3707
rect 9998 2957 10058 8059
rect 10297 7648 10617 8672
rect 10731 8124 10797 8125
rect 10731 8060 10732 8124
rect 10796 8060 10797 8124
rect 10731 8059 10797 8060
rect 10297 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10465 7648
rect 10529 7584 10545 7648
rect 10609 7584 10617 7648
rect 10297 6560 10617 7584
rect 10297 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10465 6560
rect 10529 6496 10545 6560
rect 10609 6496 10617 6560
rect 10297 5472 10617 6496
rect 10297 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10545 5472
rect 10609 5408 10617 5472
rect 10297 4384 10617 5408
rect 10734 4997 10794 8059
rect 10731 4996 10797 4997
rect 10731 4932 10732 4996
rect 10796 4932 10797 4996
rect 10731 4931 10797 4932
rect 10297 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10545 4384
rect 10609 4320 10617 4384
rect 10297 3296 10617 4320
rect 10297 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10545 3296
rect 10609 3232 10617 3296
rect 9995 2956 10061 2957
rect 9995 2892 9996 2956
rect 10060 2892 10061 2956
rect 9995 2891 10061 2892
rect 10297 2208 10617 3232
rect 10297 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10545 2208
rect 10609 2144 10617 2208
rect 10297 2128 10617 2144
rect 9811 1188 9877 1189
rect 9811 1124 9812 1188
rect 9876 1124 9877 1188
rect 9811 1123 9877 1124
rect 7787 1052 7853 1053
rect 7787 988 7788 1052
rect 7852 988 7853 1052
rect 7787 987 7853 988
rect 3923 916 3989 917
rect 3923 852 3924 916
rect 3988 852 3989 916
rect 3923 851 3989 852
use sky130_fd_sc_hd__nand3_4  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__a31oi_4  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1621208567
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1621208567
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1621208567
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3864 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1621208567
transform 1 0 4784 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 4692 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 6164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1621208567
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1621208567
transform 1 0 6440 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1621208567
transform 1 0 6532 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1621208567
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1621208567
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1621208567
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1621208567
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1621208567
transform 1 0 7544 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output103 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1621208567
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1621208567
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1621208567
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1621208567
transform 1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1621208567
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1621208567
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1621208567
transform 1 0 10304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1621208567
transform 1 0 10212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1621208567
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1621208567
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1621208567
transform 1 0 11040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1621208567
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1621208567
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1621208567
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1621208567
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1621208567
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1621208567
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1621208567
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1621208567
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1621208567
transform -1 0 12328 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1621208567
transform -1 0 12328 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _265_
timestamp 1621208567
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1621208567
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1621208567
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _255_
timestamp 1621208567
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1621208567
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1621208567
transform 1 0 3220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1621208567
transform 1 0 4140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1621208567
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1621208567
transform 1 0 4508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1621208567
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1621208567
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1621208567
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _251_
timestamp 1621208567
transform 1 0 6164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1621208567
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1621208567
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _315_
timestamp 1621208567
transform 1 0 6808 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _317_
timestamp 1621208567
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_50
timestamp 1621208567
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _241_
timestamp 1621208567
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _314_
timestamp 1621208567
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1621208567
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1621208567
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp 1621208567
transform 1 0 8556 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1621208567
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1621208567
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1621208567
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1621208567
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1621208567
transform 1 0 9476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1621208567
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1621208567
transform -1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1621208567
transform 1 0 11316 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1621208567
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1621208567
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1621208567
transform 1 0 2208 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1621208567
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1621208567
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1621208567
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1621208567
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _258_
timestamp 1621208567
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp 1621208567
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1621208567
transform 1 0 3680 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _247_
timestamp 1621208567
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _248_
timestamp 1621208567
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _319_
timestamp 1621208567
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _323_
timestamp 1621208567
transform 1 0 5796 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1621208567
transform 1 0 5520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _328_
timestamp 1621208567
transform 1 0 5244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1621208567
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_44
timestamp 1621208567
transform 1 0 5152 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1621208567
transform 1 0 7912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1621208567
transform 1 0 7452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _316_
timestamp 1621208567
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1621208567
transform 1 0 8556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1621208567
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1621208567
transform 1 0 7084 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1621208567
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _238_
timestamp 1621208567
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1621208567
transform 1 0 9292 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1621208567
transform -1 0 12328 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1621208567
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1621208567
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1621208567
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1621208567
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_105
timestamp 1621208567
transform 1 0 10764 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1621208567
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1621208567
transform 1 0 2760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _268_
timestamp 1621208567
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1621208567
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1621208567
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1621208567
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp 1621208567
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 1621208567
transform 1 0 3956 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _271_
timestamp 1621208567
transform 1 0 4232 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _338_
timestamp 1621208567
transform 1 0 4508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1621208567
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1621208567
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1621208567
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1621208567
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1621208567
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _236_
timestamp 1621208567
transform 1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1621208567
transform 1 0 5152 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1621208567
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1621208567
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1621208567
transform 1 0 7268 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1621208567
transform 1 0 9108 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1621208567
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1621208567
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1621208567
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1621208567
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1621208567
transform -1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1621208567
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1621208567
transform 1 0 11316 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1621208567
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1621208567
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1621208567
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1621208567
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _263_
timestamp 1621208567
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1621208567
transform 1 0 3128 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_41
timestamp 1621208567
transform 1 0 4876 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1621208567
transform 1 0 4968 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1621208567
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _246_
timestamp 1621208567
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _334_
timestamp 1621208567
transform 1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1621208567
transform 1 0 6532 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1621208567
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1621208567
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _229_
timestamp 1621208567
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 1621208567
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1621208567
transform 1 0 7360 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1621208567
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1621208567
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1621208567
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1621208567
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1621208567
transform 1 0 10120 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1621208567
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1621208567
transform -1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1621208567
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1621208567
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1621208567
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1621208567
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1621208567
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1621208567
transform 1 0 1748 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _278_
timestamp 1621208567
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1621208567
transform 1 0 1656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1621208567
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1621208567
transform 1 0 2852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1621208567
transform 1 0 2024 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _277_
timestamp 1621208567
transform 1 0 2576 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _272_
timestamp 1621208567
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_24
timestamp 1621208567
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1621208567
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1621208567
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1621208567
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1621208567
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1621208567
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1621208567
transform 1 0 3864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1621208567
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1621208567
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1621208567
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1621208567
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1621208567
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1621208567
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1621208567
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1621208567
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _322_
timestamp 1621208567
transform 1 0 5428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1621208567
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1621208567
transform 1 0 4968 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1621208567
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1621208567
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1621208567
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1621208567
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1621208567
transform 1 0 6532 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _212_
timestamp 1621208567
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _213_
timestamp 1621208567
transform 1 0 8004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 1621208567
transform 1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _234_
timestamp 1621208567
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1621208567
transform 1 0 7176 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1621208567
transform 1 0 8464 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1621208567
transform 1 0 8280 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1621208567
transform 1 0 7084 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1621208567
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _227_
timestamp 1621208567
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _230_
timestamp 1621208567
transform 1 0 9568 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _231_
timestamp 1621208567
transform 1 0 9844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1621208567
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1621208567
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1621208567
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1621208567
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1621208567
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1621208567
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1621208567
transform 1 0 10764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _318_
timestamp 1621208567
transform 1 0 11132 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _320_
timestamp 1621208567
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1621208567
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1621208567
transform 1 0 11960 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1621208567
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _321_
timestamp 1621208567
transform 1 0 11684 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _226_
timestamp 1621208567
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1621208567
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1621208567
transform -1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1621208567
transform 1 0 2852 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1621208567
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1621208567
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1621208567
transform 1 0 3864 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1621208567
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1621208567
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1621208567
transform 1 0 6808 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1621208567
transform 1 0 5336 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1621208567
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _219_
timestamp 1621208567
transform 1 0 8372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1621208567
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1621208567
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1621208567
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1621208567
transform 1 0 9384 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1621208567
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1621208567
transform 1 0 11040 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1621208567
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1621208567
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1621208567
transform -1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1621208567
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1621208567
transform 1 0 2576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1621208567
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1621208567
transform 1 0 2300 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1621208567
transform 1 0 2024 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1621208567
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1621208567
transform 1 0 1472 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1621208567
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1621208567
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _275_
timestamp 1621208567
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _280_
timestamp 1621208567
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1621208567
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1621208567
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1621208567
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1621208567
transform 1 0 3036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 1621208567
transform 1 0 3312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1621208567
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1621208567
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _208_
timestamp 1621208567
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _209_
timestamp 1621208567
transform 1 0 5060 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1621208567
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1621208567
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 6440 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 1621208567
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1621208567
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1621208567
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1621208567
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _224_
timestamp 1621208567
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 1621208567
transform 1 0 10120 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _223_
timestamp 1621208567
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1621208567
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1621208567
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1621208567
transform -1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1621208567
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1621208567
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_118
timestamp 1621208567
transform 1 0 11960 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _282_
timestamp 1621208567
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1621208567
transform 1 0 2392 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1621208567
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1621208567
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1621208567
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1621208567
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1621208567
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp 1621208567
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1621208567
transform 1 0 3220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1621208567
transform 1 0 4692 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1621208567
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1621208567
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_22
timestamp 1621208567
transform 1 0 3128 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_34
timestamp 1621208567
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1621208567
transform 1 0 6256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp 1621208567
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1621208567
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1621208567
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _217_
timestamp 1621208567
transform 1 0 6900 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _337_
timestamp 1621208567
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1621208567
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1621208567
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1621208567
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp 1621208567
transform 1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _221_
timestamp 1621208567
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _333_
timestamp 1621208567
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _336_
timestamp 1621208567
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1621208567
transform 1 0 10304 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1621208567
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1621208567
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _331_
timestamp 1621208567
transform 1 0 11776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1621208567
transform -1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _284_
timestamp 1621208567
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1621208567
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1621208567
transform 1 0 2852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1621208567
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1621208567
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1621208567
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1621208567
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1621208567
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1621208567
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1621208567
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _203_
timestamp 1621208567
transform 1 0 6624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _206_
timestamp 1621208567
transform 1 0 5336 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1621208567
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_50
timestamp 1621208567
transform 1 0 5704 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1621208567
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_58
timestamp 1621208567
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1621208567
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1621208567
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1621208567
transform 1 0 8740 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp 1621208567
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1621208567
transform 1 0 8832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1621208567
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9844 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1621208567
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_91
timestamp 1621208567
transform 1 0 9476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _332_
timestamp 1621208567
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1621208567
transform -1 0 12328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1621208567
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_118
timestamp 1621208567
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1621208567
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1621208567
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1621208567
transform 1 0 2852 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1621208567
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1621208567
transform 1 0 3864 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1621208567
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1621208567
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1621208567
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1621208567
transform 1 0 6164 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1621208567
transform 1 0 8556 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1621208567
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1621208567
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1621208567
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1621208567
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1621208567
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9936 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 10396 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1621208567
transform 1 0 9108 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1621208567
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1621208567
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 1621208567
transform 1 0 10856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _335_
timestamp 1621208567
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1621208567
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1621208567
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1621208567
transform -1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1621208567
transform 1 0 11960 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1621208567
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _289_
timestamp 1621208567
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1621208567
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1621208567
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1621208567
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1621208567
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1621208567
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1621208567
transform 1 0 1656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1621208567
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1621208567
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1621208567
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1621208567
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1621208567
transform 1 0 3404 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1621208567
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1621208567
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1621208567
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_38
timestamp 1621208567
transform 1 0 4600 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1621208567
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1621208567
transform 1 0 4232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _300_
timestamp 1621208567
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _297_
timestamp 1621208567
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1621208567
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1621208567
transform 1 0 5428 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_52
timestamp 1621208567
transform 1 0 5888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1621208567
transform 1 0 5520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1621208567
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1621208567
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 1621208567
transform 1 0 5612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 1621208567
transform 1 0 5244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1621208567
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1621208567
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1621208567
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1621208567
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1621208567
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 1621208567
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1621208567
transform 1 0 5520 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1621208567
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1621208567
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _304_
timestamp 1621208567
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1621208567
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1621208567
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1621208567
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1621208567
transform 1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1621208567
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _308_
timestamp 1621208567
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1621208567
transform 1 0 7084 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3_4  _162_
timestamp 1621208567
transform 1 0 8648 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1621208567
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 1621208567
transform 1 0 10212 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _172_
timestamp 1621208567
transform 1 0 9936 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1621208567
transform 1 0 10396 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9108 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1621208567
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1621208567
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_97
timestamp 1621208567
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1621208567
transform 1 0 10488 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1621208567
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1621208567
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1621208567
transform -1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1621208567
transform -1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1621208567
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1621208567
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1621208567
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_118
timestamp 1621208567
transform 1 0 11960 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1621208567
transform 1 0 2300 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1621208567
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1621208567
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1621208567
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1621208567
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_12
timestamp 1621208567
transform 1 0 2208 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1621208567
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1621208567
transform 1 0 3956 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _188_
timestamp 1621208567
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1621208567
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _192_
timestamp 1621208567
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _194_
timestamp 1621208567
transform 1 0 5428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1621208567
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1621208567
transform 1 0 6716 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1621208567
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _421_
timestamp 1621208567
transform 1 0 7268 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1621208567
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9476 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8832 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1621208567
transform 1 0 10120 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_90
timestamp 1621208567
transform 1 0 9384 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1621208567
transform -1 0 12328 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1621208567
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1621208567
transform 1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_118
timestamp 1621208567
transform 1 0 11960 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1621208567
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _291_
timestamp 1621208567
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _292_
timestamp 1621208567
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _295_
timestamp 1621208567
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1621208567
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1621208567
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_10
timestamp 1621208567
transform 1 0 2024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1621208567
transform 1 0 2392 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _294_
timestamp 1621208567
transform 1 0 3312 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _298_
timestamp 1621208567
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1621208567
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1621208567
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1621208567
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1621208567
transform 1 0 4508 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1621208567
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1621208567
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_40
timestamp 1621208567
transform 1 0 4784 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1621208567
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _197_
timestamp 1621208567
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1621208567
transform 1 0 6072 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1621208567
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1621208567
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1621208567
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1621208567
transform 1 0 8464 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1621208567
transform 1 0 7728 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1621208567
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_79
timestamp 1621208567
transform 1 0 8372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1621208567
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9568 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 10304 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1621208567
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1621208567
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1621208567
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1621208567
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _167_
timestamp 1621208567
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1621208567
transform -1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1621208567
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1621208567
transform 1 0 11960 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1621208567
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1621208567
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1621208567
transform 1 0 2484 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1621208567
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _195_
timestamp 1621208567
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1621208567
transform 1 0 4416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1621208567
transform 1 0 3956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1621208567
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1621208567
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1621208567
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _189_
timestamp 1621208567
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1621208567
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1621208567
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1621208567
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1621208567
transform 1 0 5796 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1621208567
transform 1 0 6072 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1621208567
transform 1 0 7728 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1621208567
transform 1 0 7452 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1621208567
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1621208567
transform 1 0 7084 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _161_
timestamp 1621208567
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _164_
timestamp 1621208567
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9292 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1621208567
transform 1 0 10672 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1621208567
transform 1 0 9200 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1621208567
transform -1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1621208567
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1621208567
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1621208567
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1621208567
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1621208567
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1621208567
transform 1 0 1380 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1621208567
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1621208567
transform 1 0 3864 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1621208567
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1621208567
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1621208567
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1621208567
transform 1 0 5336 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1621208567
transform 1 0 6808 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__o21bai_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8280 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _165_
timestamp 1621208567
transform 1 0 9844 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9108 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1621208567
transform 1 0 10120 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1621208567
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1621208567
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1621208567
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _345_
timestamp 1621208567
transform 1 0 11592 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1621208567
transform -1 0 12328 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_118
timestamp 1621208567
transform 1 0 11960 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1621208567
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1621208567
transform -1 0 2208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1621208567
transform -1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1621208567
transform -1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform -1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1621208567
transform -1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1621208567
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_12
timestamp 1621208567
transform 1 0 2208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _198_
timestamp 1621208567
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1621208567
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1621208567
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1621208567
transform 1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1621208567
transform -1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1621208567
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1621208567
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1621208567
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_30
timestamp 1621208567
transform 1 0 3864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _347_
timestamp 1621208567
transform 1 0 4968 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp 1621208567
transform 1 0 5612 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp 1621208567
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1621208567
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1621208567
transform 1 0 5336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1621208567
transform 1 0 6532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1621208567
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1621208567
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _312_
timestamp 1621208567
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _350_
timestamp 1621208567
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1621208567
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1621208567
transform 1 0 7544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1621208567
transform 1 0 8188 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1621208567
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1621208567
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1621208567
transform 1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1621208567
transform 1 0 10028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1621208567
transform 1 0 9660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1621208567
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_88
timestamp 1621208567
transform 1 0 9200 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1621208567
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1621208567
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1621208567
transform -1 0 12328 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1621208567
transform 1 0 11776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1621208567
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1621208567
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1621208567
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1621208567
transform 1 0 11868 0 1 12512
box -38 -48 222 592
<< labels >>
rlabel metal2 s 11150 14818 11206 15618 6 cfg_bit_out
port 0 nsew signal tristate
rlabel metal2 s 12622 14818 12678 15618 6 cfg_bit_out_valid
port 1 nsew signal tristate
rlabel metal2 s 9678 14818 9734 15618 6 cfg_out_start
port 2 nsew signal tristate
rlabel metal2 s 3698 14818 3754 15618 6 col_sel[0]
port 3 nsew signal tristate
rlabel metal2 s 5170 14818 5226 15618 6 col_sel[1]
port 4 nsew signal tristate
rlabel metal2 s 6642 14818 6698 15618 6 col_sel[2]
port 5 nsew signal tristate
rlabel metal2 s 8206 14818 8262 15618 6 col_sel[3]
port 6 nsew signal tristate
rlabel metal2 s 754 14818 810 15618 6 wb_clk_i
port 7 nsew signal input
rlabel metal2 s 2226 14818 2282 15618 6 wb_rst_i
port 8 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_ack_o
port 9 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[0]
port 10 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[10]
port 11 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[11]
port 12 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[12]
port 13 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[13]
port 14 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[14]
port 15 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[15]
port 16 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[16]
port 17 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[17]
port 18 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[18]
port 19 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[19]
port 20 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[1]
port 21 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[20]
port 22 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[21]
port 23 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[22]
port 24 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[23]
port 25 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[24]
port 26 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[25]
port 27 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[26]
port 28 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[27]
port 29 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[28]
port 30 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[29]
port 31 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[2]
port 32 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[30]
port 33 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[31]
port 34 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[3]
port 35 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[4]
port 36 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[5]
port 37 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[6]
port 38 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[7]
port 39 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_adr_i[8]
port 40 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[9]
port 41 nsew signal input
rlabel metal2 s 110 0 166 800 6 wbs_cyc_i
port 42 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_dat_i[0]
port 43 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[10]
port 44 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[11]
port 45 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[12]
port 46 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[13]
port 47 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[14]
port 48 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[15]
port 49 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[16]
port 50 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[17]
port 51 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[18]
port 52 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[19]
port 53 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 54 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[20]
port 55 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[21]
port 56 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[22]
port 57 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[23]
port 58 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[24]
port 59 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[25]
port 60 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[26]
port 61 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[27]
port 62 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[28]
port 63 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[29]
port 64 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_dat_i[2]
port 65 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[30]
port 66 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[31]
port 67 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_dat_i[3]
port 68 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[4]
port 69 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[5]
port 70 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[6]
port 71 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[7]
port 72 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[8]
port 73 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_i[9]
port 74 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[0]
port 75 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[10]
port 76 nsew signal tristate
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[11]
port 77 nsew signal tristate
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[12]
port 78 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[13]
port 79 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 80 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[15]
port 81 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[16]
port 82 nsew signal tristate
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[17]
port 83 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[18]
port 84 nsew signal tristate
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[19]
port 85 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[1]
port 86 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[20]
port 87 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[21]
port 88 nsew signal tristate
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[22]
port 89 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[23]
port 90 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[24]
port 91 nsew signal tristate
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[25]
port 92 nsew signal tristate
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[26]
port 93 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[27]
port 94 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[28]
port 95 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[29]
port 96 nsew signal tristate
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[2]
port 97 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[30]
port 98 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[31]
port 99 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[3]
port 100 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[4]
port 101 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 102 nsew signal tristate
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[6]
port 103 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[7]
port 104 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[8]
port 105 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[9]
port 106 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 wbs_sel_i[0]
port 107 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_sel_i[1]
port 108 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_sel_i[2]
port 109 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_sel_i[3]
port 110 nsew signal input
rlabel metal2 s 18 0 74 800 6 wbs_stb_i
port 111 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_we_i
port 112 nsew signal input
rlabel metal4 s 10297 2128 10617 13104 6 VPWR
port 113 nsew power bidirectional
rlabel metal4 s 6556 2128 6876 13104 6 VPWR
port 114 nsew power bidirectional
rlabel metal4 s 2815 2128 3135 13104 6 VPWR
port 115 nsew power bidirectional
rlabel metal4 s 8427 2128 8747 13104 6 VGND
port 116 nsew ground bidirectional
rlabel metal4 s 4685 2128 5005 13104 6 VGND
port 117 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 13474 15618
<< end >>
