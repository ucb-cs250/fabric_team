VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 274.470 BY 285.190 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 281.190 255.210 285.190 ;
    END
  END COUT
  PIN cb_e_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 2.760 274.470 3.360 ;
    END
  END cb_e_clb1_input[0]
  PIN cb_e_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 8.880 274.470 9.480 ;
    END
  END cb_e_clb1_input[1]
  PIN cb_e_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 15.000 274.470 15.600 ;
    END
  END cb_e_clb1_input[2]
  PIN cb_e_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 21.120 274.470 21.720 ;
    END
  END cb_e_clb1_input[3]
  PIN cb_e_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 27.240 274.470 27.840 ;
    END
  END cb_e_clb1_input[4]
  PIN cb_e_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 33.360 274.470 33.960 ;
    END
  END cb_e_clb1_input[5]
  PIN cb_e_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 39.480 274.470 40.080 ;
    END
  END cb_e_clb1_input[6]
  PIN cb_e_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 45.600 274.470 46.200 ;
    END
  END cb_e_clb1_input[7]
  PIN cb_e_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 51.720 274.470 52.320 ;
    END
  END cb_e_clb1_input[8]
  PIN cb_e_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 57.840 274.470 58.440 ;
    END
  END cb_e_clb1_input[9]
  PIN cb_e_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 64.640 274.470 65.240 ;
    END
  END cb_e_clb1_output[0]
  PIN cb_e_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 70.760 274.470 71.360 ;
    END
  END cb_e_clb1_output[1]
  PIN cb_e_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 76.880 274.470 77.480 ;
    END
  END cb_e_clb1_output[2]
  PIN cb_e_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 83.000 274.470 83.600 ;
    END
  END cb_e_clb1_output[3]
  PIN cb_e_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END cb_e_single1_in[0]
  PIN cb_e_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END cb_e_single1_in[10]
  PIN cb_e_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END cb_e_single1_in[11]
  PIN cb_e_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END cb_e_single1_in[12]
  PIN cb_e_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END cb_e_single1_in[13]
  PIN cb_e_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END cb_e_single1_in[14]
  PIN cb_e_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END cb_e_single1_in[15]
  PIN cb_e_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END cb_e_single1_in[1]
  PIN cb_e_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END cb_e_single1_in[2]
  PIN cb_e_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END cb_e_single1_in[3]
  PIN cb_e_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END cb_e_single1_in[4]
  PIN cb_e_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END cb_e_single1_in[5]
  PIN cb_e_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END cb_e_single1_in[6]
  PIN cb_e_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END cb_e_single1_in[7]
  PIN cb_e_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END cb_e_single1_in[8]
  PIN cb_e_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cb_e_single1_in[9]
  PIN cb_e_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END cb_e_single1_out[0]
  PIN cb_e_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END cb_e_single1_out[10]
  PIN cb_e_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END cb_e_single1_out[11]
  PIN cb_e_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END cb_e_single1_out[12]
  PIN cb_e_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END cb_e_single1_out[13]
  PIN cb_e_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END cb_e_single1_out[14]
  PIN cb_e_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END cb_e_single1_out[15]
  PIN cb_e_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END cb_e_single1_out[1]
  PIN cb_e_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END cb_e_single1_out[2]
  PIN cb_e_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END cb_e_single1_out[3]
  PIN cb_e_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END cb_e_single1_out[4]
  PIN cb_e_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END cb_e_single1_out[5]
  PIN cb_e_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END cb_e_single1_out[6]
  PIN cb_e_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END cb_e_single1_out[7]
  PIN cb_e_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END cb_e_single1_out[8]
  PIN cb_e_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END cb_e_single1_out[9]
  PIN cb_n_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 281.190 2.670 285.190 ;
    END
  END cb_n_clb1_input[0]
  PIN cb_n_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 281.190 7.730 285.190 ;
    END
  END cb_n_clb1_input[1]
  PIN cb_n_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 281.190 13.250 285.190 ;
    END
  END cb_n_clb1_input[2]
  PIN cb_n_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 281.190 18.770 285.190 ;
    END
  END cb_n_clb1_input[3]
  PIN cb_n_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 281.190 24.290 285.190 ;
    END
  END cb_n_clb1_input[4]
  PIN cb_n_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 281.190 29.810 285.190 ;
    END
  END cb_n_clb1_input[5]
  PIN cb_n_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 281.190 35.330 285.190 ;
    END
  END cb_n_clb1_input[6]
  PIN cb_n_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 281.190 40.850 285.190 ;
    END
  END cb_n_clb1_input[7]
  PIN cb_n_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 281.190 46.370 285.190 ;
    END
  END cb_n_clb1_input[8]
  PIN cb_n_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 281.190 51.890 285.190 ;
    END
  END cb_n_clb1_input[9]
  PIN cb_n_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 281.190 57.410 285.190 ;
    END
  END cb_n_clb1_output[0]
  PIN cb_n_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 281.190 62.930 285.190 ;
    END
  END cb_n_clb1_output[1]
  PIN cb_n_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 281.190 68.450 285.190 ;
    END
  END cb_n_clb1_output[2]
  PIN cb_n_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 281.190 73.970 285.190 ;
    END
  END cb_n_clb1_output[3]
  PIN cb_n_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END cb_n_single1_in[0]
  PIN cb_n_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END cb_n_single1_in[10]
  PIN cb_n_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END cb_n_single1_in[11]
  PIN cb_n_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END cb_n_single1_in[12]
  PIN cb_n_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END cb_n_single1_in[13]
  PIN cb_n_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END cb_n_single1_in[14]
  PIN cb_n_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END cb_n_single1_in[15]
  PIN cb_n_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END cb_n_single1_in[1]
  PIN cb_n_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END cb_n_single1_in[2]
  PIN cb_n_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END cb_n_single1_in[3]
  PIN cb_n_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END cb_n_single1_in[4]
  PIN cb_n_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END cb_n_single1_in[5]
  PIN cb_n_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END cb_n_single1_in[6]
  PIN cb_n_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END cb_n_single1_in[7]
  PIN cb_n_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END cb_n_single1_in[8]
  PIN cb_n_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END cb_n_single1_in[9]
  PIN cb_n_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END cb_n_single1_out[0]
  PIN cb_n_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END cb_n_single1_out[10]
  PIN cb_n_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END cb_n_single1_out[11]
  PIN cb_n_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END cb_n_single1_out[12]
  PIN cb_n_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END cb_n_single1_out[13]
  PIN cb_n_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END cb_n_single1_out[14]
  PIN cb_n_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END cb_n_single1_out[15]
  PIN cb_n_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END cb_n_single1_out[1]
  PIN cb_n_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END cb_n_single1_out[2]
  PIN cb_n_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END cb_n_single1_out[3]
  PIN cb_n_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END cb_n_single1_out[4]
  PIN cb_n_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END cb_n_single1_out[5]
  PIN cb_n_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END cb_n_single1_out[6]
  PIN cb_n_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END cb_n_single1_out[7]
  PIN cb_n_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END cb_n_single1_out[8]
  PIN cb_n_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END cb_n_single1_out[9]
  PIN cfg_bit_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END cfg_bit_in
  PIN cfg_bit_in_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END cfg_bit_in_valid
  PIN cfg_bit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 281.190 266.250 285.190 ;
    END
  END cfg_bit_out
  PIN cfg_bit_out_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 281.190 271.770 285.190 ;
    END
  END cfg_bit_out_valid
  PIN cfg_in_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END cfg_in_start
  PIN cfg_out_start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 281.190 260.730 285.190 ;
    END
  END cfg_out_start
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END clb_south_out[3]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END clb_west_out[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END clk
  PIN crst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END crst
  PIN sb_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 89.120 274.470 89.720 ;
    END
  END sb_east_in[0]
  PIN sb_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 151.000 274.470 151.600 ;
    END
  END sb_east_in[10]
  PIN sb_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 157.120 274.470 157.720 ;
    END
  END sb_east_in[11]
  PIN sb_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 163.240 274.470 163.840 ;
    END
  END sb_east_in[12]
  PIN sb_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 169.360 274.470 169.960 ;
    END
  END sb_east_in[13]
  PIN sb_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 176.160 274.470 176.760 ;
    END
  END sb_east_in[14]
  PIN sb_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 182.280 274.470 182.880 ;
    END
  END sb_east_in[15]
  PIN sb_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 95.240 274.470 95.840 ;
    END
  END sb_east_in[1]
  PIN sb_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 101.360 274.470 101.960 ;
    END
  END sb_east_in[2]
  PIN sb_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 107.480 274.470 108.080 ;
    END
  END sb_east_in[3]
  PIN sb_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 113.600 274.470 114.200 ;
    END
  END sb_east_in[4]
  PIN sb_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 120.400 274.470 121.000 ;
    END
  END sb_east_in[5]
  PIN sb_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 126.520 274.470 127.120 ;
    END
  END sb_east_in[6]
  PIN sb_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 132.640 274.470 133.240 ;
    END
  END sb_east_in[7]
  PIN sb_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 138.760 274.470 139.360 ;
    END
  END sb_east_in[8]
  PIN sb_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 144.880 274.470 145.480 ;
    END
  END sb_east_in[9]
  PIN sb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 188.400 274.470 189.000 ;
    END
  END sb_east_out[0]
  PIN sb_east_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 250.280 274.470 250.880 ;
    END
  END sb_east_out[10]
  PIN sb_east_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 256.400 274.470 257.000 ;
    END
  END sb_east_out[11]
  PIN sb_east_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 262.520 274.470 263.120 ;
    END
  END sb_east_out[12]
  PIN sb_east_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 268.640 274.470 269.240 ;
    END
  END sb_east_out[13]
  PIN sb_east_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 274.760 274.470 275.360 ;
    END
  END sb_east_out[14]
  PIN sb_east_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 280.880 274.470 281.480 ;
    END
  END sb_east_out[15]
  PIN sb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 194.520 274.470 195.120 ;
    END
  END sb_east_out[1]
  PIN sb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 200.640 274.470 201.240 ;
    END
  END sb_east_out[2]
  PIN sb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 206.760 274.470 207.360 ;
    END
  END sb_east_out[3]
  PIN sb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 212.880 274.470 213.480 ;
    END
  END sb_east_out[4]
  PIN sb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 219.000 274.470 219.600 ;
    END
  END sb_east_out[5]
  PIN sb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 225.120 274.470 225.720 ;
    END
  END sb_east_out[6]
  PIN sb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 231.920 274.470 232.520 ;
    END
  END sb_east_out[7]
  PIN sb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 238.040 274.470 238.640 ;
    END
  END sb_east_out[8]
  PIN sb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 270.470 244.160 274.470 244.760 ;
    END
  END sb_east_out[9]
  PIN sb_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 281.190 79.490 285.190 ;
    END
  END sb_north_in[0]
  PIN sb_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 281.190 134.230 285.190 ;
    END
  END sb_north_in[10]
  PIN sb_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 281.190 139.750 285.190 ;
    END
  END sb_north_in[11]
  PIN sb_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 281.190 145.270 285.190 ;
    END
  END sb_north_in[12]
  PIN sb_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 281.190 150.790 285.190 ;
    END
  END sb_north_in[13]
  PIN sb_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 281.190 156.310 285.190 ;
    END
  END sb_north_in[14]
  PIN sb_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 281.190 161.830 285.190 ;
    END
  END sb_north_in[15]
  PIN sb_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 281.190 85.010 285.190 ;
    END
  END sb_north_in[1]
  PIN sb_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 281.190 90.530 285.190 ;
    END
  END sb_north_in[2]
  PIN sb_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 281.190 95.590 285.190 ;
    END
  END sb_north_in[3]
  PIN sb_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 281.190 101.110 285.190 ;
    END
  END sb_north_in[4]
  PIN sb_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 281.190 106.630 285.190 ;
    END
  END sb_north_in[5]
  PIN sb_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 281.190 112.150 285.190 ;
    END
  END sb_north_in[6]
  PIN sb_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 281.190 117.670 285.190 ;
    END
  END sb_north_in[7]
  PIN sb_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 281.190 123.190 285.190 ;
    END
  END sb_north_in[8]
  PIN sb_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 281.190 128.710 285.190 ;
    END
  END sb_north_in[9]
  PIN sb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 281.190 167.350 285.190 ;
    END
  END sb_north_out[0]
  PIN sb_north_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 281.190 222.090 285.190 ;
    END
  END sb_north_out[10]
  PIN sb_north_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 281.190 227.610 285.190 ;
    END
  END sb_north_out[11]
  PIN sb_north_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 281.190 233.130 285.190 ;
    END
  END sb_north_out[12]
  PIN sb_north_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 281.190 238.650 285.190 ;
    END
  END sb_north_out[13]
  PIN sb_north_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 281.190 244.170 285.190 ;
    END
  END sb_north_out[14]
  PIN sb_north_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 281.190 249.690 285.190 ;
    END
  END sb_north_out[15]
  PIN sb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 281.190 172.870 285.190 ;
    END
  END sb_north_out[1]
  PIN sb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 281.190 178.390 285.190 ;
    END
  END sb_north_out[2]
  PIN sb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 281.190 183.910 285.190 ;
    END
  END sb_north_out[3]
  PIN sb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 281.190 188.970 285.190 ;
    END
  END sb_north_out[4]
  PIN sb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 281.190 194.490 285.190 ;
    END
  END sb_north_out[5]
  PIN sb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 281.190 200.010 285.190 ;
    END
  END sb_north_out[6]
  PIN sb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 281.190 205.530 285.190 ;
    END
  END sb_north_out[7]
  PIN sb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 281.190 211.050 285.190 ;
    END
  END sb_north_out[8]
  PIN sb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 281.190 216.570 285.190 ;
    END
  END sb_north_out[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 272.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 272.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 272.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 272.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 7.905 269.415 272.085 ;
      LAYER met1 ;
        RECT 2.370 6.840 271.790 275.360 ;
      LAYER met2 ;
        RECT 2.950 280.910 7.170 281.365 ;
        RECT 8.010 280.910 12.690 281.365 ;
        RECT 13.530 280.910 18.210 281.365 ;
        RECT 19.050 280.910 23.730 281.365 ;
        RECT 24.570 280.910 29.250 281.365 ;
        RECT 30.090 280.910 34.770 281.365 ;
        RECT 35.610 280.910 40.290 281.365 ;
        RECT 41.130 280.910 45.810 281.365 ;
        RECT 46.650 280.910 51.330 281.365 ;
        RECT 52.170 280.910 56.850 281.365 ;
        RECT 57.690 280.910 62.370 281.365 ;
        RECT 63.210 280.910 67.890 281.365 ;
        RECT 68.730 280.910 73.410 281.365 ;
        RECT 74.250 280.910 78.930 281.365 ;
        RECT 79.770 280.910 84.450 281.365 ;
        RECT 85.290 280.910 89.970 281.365 ;
        RECT 90.810 280.910 95.030 281.365 ;
        RECT 95.870 280.910 100.550 281.365 ;
        RECT 101.390 280.910 106.070 281.365 ;
        RECT 106.910 280.910 111.590 281.365 ;
        RECT 112.430 280.910 117.110 281.365 ;
        RECT 117.950 280.910 122.630 281.365 ;
        RECT 123.470 280.910 128.150 281.365 ;
        RECT 128.990 280.910 133.670 281.365 ;
        RECT 134.510 280.910 139.190 281.365 ;
        RECT 140.030 280.910 144.710 281.365 ;
        RECT 145.550 280.910 150.230 281.365 ;
        RECT 151.070 280.910 155.750 281.365 ;
        RECT 156.590 280.910 161.270 281.365 ;
        RECT 162.110 280.910 166.790 281.365 ;
        RECT 167.630 280.910 172.310 281.365 ;
        RECT 173.150 280.910 177.830 281.365 ;
        RECT 178.670 280.910 183.350 281.365 ;
        RECT 184.190 280.910 188.410 281.365 ;
        RECT 189.250 280.910 193.930 281.365 ;
        RECT 194.770 280.910 199.450 281.365 ;
        RECT 200.290 280.910 204.970 281.365 ;
        RECT 205.810 280.910 210.490 281.365 ;
        RECT 211.330 280.910 216.010 281.365 ;
        RECT 216.850 280.910 221.530 281.365 ;
        RECT 222.370 280.910 227.050 281.365 ;
        RECT 227.890 280.910 232.570 281.365 ;
        RECT 233.410 280.910 238.090 281.365 ;
        RECT 238.930 280.910 243.610 281.365 ;
        RECT 244.450 280.910 249.130 281.365 ;
        RECT 249.970 280.910 254.650 281.365 ;
        RECT 255.490 280.910 260.170 281.365 ;
        RECT 261.010 280.910 265.690 281.365 ;
        RECT 266.530 280.910 271.210 281.365 ;
        RECT 2.400 4.280 271.760 280.910 ;
        RECT 2.950 2.875 7.170 4.280 ;
        RECT 8.010 2.875 12.230 4.280 ;
        RECT 13.070 2.875 17.750 4.280 ;
        RECT 18.590 2.875 22.810 4.280 ;
        RECT 23.650 2.875 28.330 4.280 ;
        RECT 29.170 2.875 33.390 4.280 ;
        RECT 34.230 2.875 38.910 4.280 ;
        RECT 39.750 2.875 43.970 4.280 ;
        RECT 44.810 2.875 49.490 4.280 ;
        RECT 50.330 2.875 54.550 4.280 ;
        RECT 55.390 2.875 60.070 4.280 ;
        RECT 60.910 2.875 65.130 4.280 ;
        RECT 65.970 2.875 70.650 4.280 ;
        RECT 71.490 2.875 75.710 4.280 ;
        RECT 76.550 2.875 81.230 4.280 ;
        RECT 82.070 2.875 86.290 4.280 ;
        RECT 87.130 2.875 91.810 4.280 ;
        RECT 92.650 2.875 96.870 4.280 ;
        RECT 97.710 2.875 102.390 4.280 ;
        RECT 103.230 2.875 107.450 4.280 ;
        RECT 108.290 2.875 112.970 4.280 ;
        RECT 113.810 2.875 118.030 4.280 ;
        RECT 118.870 2.875 123.550 4.280 ;
        RECT 124.390 2.875 128.610 4.280 ;
        RECT 129.450 2.875 134.130 4.280 ;
        RECT 134.970 2.875 139.190 4.280 ;
        RECT 140.030 2.875 144.250 4.280 ;
        RECT 145.090 2.875 149.770 4.280 ;
        RECT 150.610 2.875 154.830 4.280 ;
        RECT 155.670 2.875 160.350 4.280 ;
        RECT 161.190 2.875 165.410 4.280 ;
        RECT 166.250 2.875 170.930 4.280 ;
        RECT 171.770 2.875 175.990 4.280 ;
        RECT 176.830 2.875 181.510 4.280 ;
        RECT 182.350 2.875 186.570 4.280 ;
        RECT 187.410 2.875 192.090 4.280 ;
        RECT 192.930 2.875 197.150 4.280 ;
        RECT 197.990 2.875 202.670 4.280 ;
        RECT 203.510 2.875 207.730 4.280 ;
        RECT 208.570 2.875 213.250 4.280 ;
        RECT 214.090 2.875 218.310 4.280 ;
        RECT 219.150 2.875 223.830 4.280 ;
        RECT 224.670 2.875 228.890 4.280 ;
        RECT 229.730 2.875 234.410 4.280 ;
        RECT 235.250 2.875 239.470 4.280 ;
        RECT 240.310 2.875 244.990 4.280 ;
        RECT 245.830 2.875 250.050 4.280 ;
        RECT 250.890 2.875 255.570 4.280 ;
        RECT 256.410 2.875 260.630 4.280 ;
        RECT 261.470 2.875 266.150 4.280 ;
        RECT 266.990 2.875 271.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 280.480 270.070 281.345 ;
        RECT 4.000 275.760 270.470 280.480 ;
        RECT 4.400 274.360 270.070 275.760 ;
        RECT 4.000 269.640 270.470 274.360 ;
        RECT 4.400 268.240 270.070 269.640 ;
        RECT 4.000 263.520 270.470 268.240 ;
        RECT 4.400 262.120 270.070 263.520 ;
        RECT 4.000 257.400 270.470 262.120 ;
        RECT 4.400 256.000 270.070 257.400 ;
        RECT 4.000 251.280 270.470 256.000 ;
        RECT 4.400 249.880 270.070 251.280 ;
        RECT 4.000 245.160 270.470 249.880 ;
        RECT 4.400 243.760 270.070 245.160 ;
        RECT 4.000 239.040 270.470 243.760 ;
        RECT 4.400 237.640 270.070 239.040 ;
        RECT 4.000 232.920 270.470 237.640 ;
        RECT 4.400 231.520 270.070 232.920 ;
        RECT 4.000 226.120 270.470 231.520 ;
        RECT 4.400 224.720 270.070 226.120 ;
        RECT 4.000 220.000 270.470 224.720 ;
        RECT 4.400 218.600 270.070 220.000 ;
        RECT 4.000 213.880 270.470 218.600 ;
        RECT 4.400 212.480 270.070 213.880 ;
        RECT 4.000 207.760 270.470 212.480 ;
        RECT 4.400 206.360 270.070 207.760 ;
        RECT 4.000 201.640 270.470 206.360 ;
        RECT 4.400 200.240 270.070 201.640 ;
        RECT 4.000 195.520 270.470 200.240 ;
        RECT 4.400 194.120 270.070 195.520 ;
        RECT 4.000 189.400 270.470 194.120 ;
        RECT 4.400 188.000 270.070 189.400 ;
        RECT 4.000 183.280 270.470 188.000 ;
        RECT 4.400 181.880 270.070 183.280 ;
        RECT 4.000 177.160 270.470 181.880 ;
        RECT 4.400 175.760 270.070 177.160 ;
        RECT 4.000 170.360 270.470 175.760 ;
        RECT 4.400 168.960 270.070 170.360 ;
        RECT 4.000 164.240 270.470 168.960 ;
        RECT 4.400 162.840 270.070 164.240 ;
        RECT 4.000 158.120 270.470 162.840 ;
        RECT 4.400 156.720 270.070 158.120 ;
        RECT 4.000 152.000 270.470 156.720 ;
        RECT 4.400 150.600 270.070 152.000 ;
        RECT 4.000 145.880 270.470 150.600 ;
        RECT 4.400 144.480 270.070 145.880 ;
        RECT 4.000 139.760 270.470 144.480 ;
        RECT 4.400 138.360 270.070 139.760 ;
        RECT 4.000 133.640 270.470 138.360 ;
        RECT 4.400 132.240 270.070 133.640 ;
        RECT 4.000 127.520 270.470 132.240 ;
        RECT 4.400 126.120 270.070 127.520 ;
        RECT 4.000 121.400 270.470 126.120 ;
        RECT 4.400 120.000 270.070 121.400 ;
        RECT 4.000 114.600 270.470 120.000 ;
        RECT 4.400 113.200 270.070 114.600 ;
        RECT 4.000 108.480 270.470 113.200 ;
        RECT 4.400 107.080 270.070 108.480 ;
        RECT 4.000 102.360 270.470 107.080 ;
        RECT 4.400 100.960 270.070 102.360 ;
        RECT 4.000 96.240 270.470 100.960 ;
        RECT 4.400 94.840 270.070 96.240 ;
        RECT 4.000 90.120 270.470 94.840 ;
        RECT 4.400 88.720 270.070 90.120 ;
        RECT 4.000 84.000 270.470 88.720 ;
        RECT 4.400 82.600 270.070 84.000 ;
        RECT 4.000 77.880 270.470 82.600 ;
        RECT 4.400 76.480 270.070 77.880 ;
        RECT 4.000 71.760 270.470 76.480 ;
        RECT 4.400 70.360 270.070 71.760 ;
        RECT 4.000 65.640 270.470 70.360 ;
        RECT 4.400 64.240 270.070 65.640 ;
        RECT 4.000 58.840 270.470 64.240 ;
        RECT 4.400 57.440 270.070 58.840 ;
        RECT 4.000 52.720 270.470 57.440 ;
        RECT 4.400 51.320 270.070 52.720 ;
        RECT 4.000 46.600 270.470 51.320 ;
        RECT 4.400 45.200 270.070 46.600 ;
        RECT 4.000 40.480 270.470 45.200 ;
        RECT 4.400 39.080 270.070 40.480 ;
        RECT 4.000 34.360 270.470 39.080 ;
        RECT 4.400 32.960 270.070 34.360 ;
        RECT 4.000 28.240 270.470 32.960 ;
        RECT 4.400 26.840 270.070 28.240 ;
        RECT 4.000 22.120 270.470 26.840 ;
        RECT 4.400 20.720 270.070 22.120 ;
        RECT 4.000 16.000 270.470 20.720 ;
        RECT 4.400 14.600 270.070 16.000 ;
        RECT 4.000 9.880 270.470 14.600 ;
        RECT 4.400 8.480 270.070 9.880 ;
        RECT 4.000 3.760 270.470 8.480 ;
        RECT 4.400 2.895 270.070 3.760 ;
      LAYER met4 ;
        RECT 7.655 11.055 20.640 269.105 ;
        RECT 23.040 11.055 97.440 269.105 ;
        RECT 99.840 11.055 174.240 269.105 ;
        RECT 176.640 11.055 251.040 269.105 ;
        RECT 253.440 11.055 260.065 269.105 ;
  END
END clb_tile
END LIBRARY

