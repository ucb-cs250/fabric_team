module clb_tile (carry_in,
    carry_out,
    cen,
    clk,
    rst,
    set_in_hard,
    set_out_hard,
    shift_in_hard,
    shift_out_hard,
    VPWR,
    VGND,
    cb_east_in,
    cb_east_out,
    cb_north_in,
    cb_north_out,
    clb_south_in,
    clb_south_out,
    clb_west_in,
    clb_west_out,
    east_double,
    east_single,
    north_double,
    north_single,
    south_double,
    south_single,
    west_double,
    west_single);
 input carry_in;
 output carry_out;
 input cen;
 input clk;
 input rst;
 input set_in_hard;
 output set_out_hard;
 input shift_in_hard;
 output shift_out_hard;
 input VPWR;
 input VGND;
 input [4:0] cb_east_in;
 output [9:0] cb_east_out;
 input [4:0] cb_north_in;
 output [9:0] cb_north_out;
 input [9:0] clb_south_in;
 output [4:0] clb_south_out;
 input [9:0] clb_west_in;
 output [4:0] clb_west_out;
 inout [7:0] east_double;
 inout [3:0] east_single;
 inout [7:0] north_double;
 inout [3:0] north_single;
 inout [7:0] south_double;
 inout [3:0] south_single;
 inout [7:0] west_double;
 inout [3:0] west_single;

 sky130_fd_sc_hd__mux2_1 _04316_ (.A0(set_in_hard),
    .A1(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ),
    .S(\slice.configuroni.input_mux ),
    .X(set_out_hard));
 sky130_fd_sc_hd__mux2_1 _04317_ (.A0(\slice.sliceluroni.cc.P[0] ),
    .A1(\slice.sliceluroni.cc.P[1] ),
    .S(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _04318_ (.A0(\slice.sliceluroni.cc.P[0] ),
    .A1(_00090_),
    .S(\slice.sliceluroni.muxes.config_state[0] ),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _04319_ (.A0(\slice.sliceluroni.cc.P[2] ),
    .A1(\slice.sliceluroni.cc.P[3] ),
    .S(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _04320_ (.A0(\slice.sliceluroni.cc.P[2] ),
    .A1(_00092_),
    .S(\slice.sliceluroni.muxes.config_state[0] ),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _04321_ (.A0(_00091_),
    .A1(_00093_),
    .S(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _04322_ (.A0(_00091_),
    .A1(_00094_),
    .S(\slice.sliceluroni.muxes.config_state[1] ),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _04323_ (.A0(_00095_),
    .A1(_00096_),
    .S(\slice.sliceluroni.use_cc ),
    .X(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ));
 sky130_fd_sc_hd__mux2_1 _04324_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(carry_in),
    .S(\slice.sliceluroni.cc.P[0] ),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _04325_ (.A0(\slice.sliceluroni.cc.P[1] ),
    .A1(_00098_),
    .S(\slice.sliceluroni.use_cc ),
    .X(clb_south_out[0]));
 sky130_fd_sc_hd__mux2_1 _04326_ (.A0(clb_south_out[1]),
    .A1(_00097_),
    .S(\slice.sliceluroni.cc.P[1] ),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _04327_ (.A0(_00093_),
    .A1(_00100_),
    .S(\slice.sliceluroni.use_cc ),
    .X(clb_west_out[0]));
 sky130_fd_sc_hd__mux2_1 _04328_ (.A0(clb_west_out[1]),
    .A1(_00099_),
    .S(\slice.sliceluroni.cc.P[2] ),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _04329_ (.A0(\slice.sliceluroni.cc.P[3] ),
    .A1(_00102_),
    .S(\slice.sliceluroni.use_cc ),
    .X(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ));
 sky130_fd_sc_hd__mux2_1 _04330_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .A1(\slice.configuroni.mem_config[6] ),
    .S(_00089_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _04331_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(\slice.configuroni.mem_config[7] ),
    .S(_00089_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _04332_ (.A0(clb_west_out[0]),
    .A1(\slice.configuroni.mem_config[4] ),
    .S(_00089_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _04333_ (.A0(clb_west_out[1]),
    .A1(\slice.configuroni.mem_config[5] ),
    .S(_00089_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _04334_ (.A0(clb_south_out[0]),
    .A1(\slice.configuroni.mem_config[2] ),
    .S(_00089_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _04335_ (.A0(clb_south_out[1]),
    .A1(\slice.configuroni.mem_config[3] ),
    .S(_00089_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _04336_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .A1(\cb_north.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .S(_00089_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _04337_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(\slice.configuroni.mem_config[1] ),
    .S(_00089_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _04338_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(_00101_),
    .S(\slice.sliceluroni.cc.P[3] ),
    .X(carry_out));
 sky130_fd_sc_hd__mux2_1 _04339_ (.A0(shift_in_hard),
    .A1(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ),
    .S(\slice.configuroni.input_mux ),
    .X(\slice.configuroni.comb_shifter.head_bit.shift_in ));
 sky130_fd_sc_hd__mux2_1 _04340_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ),
    .S(_04168_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _04341_ (.A0(clb_south_out[1]),
    .A1(clb_south_in[3]),
    .S(_04217_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _04342_ (.A0(clb_west_out[1]),
    .A1(clb_west_in[3]),
    .S(_04266_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _04343_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .A1(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ),
    .S(_04315_),
    .X(_00106_));
 sky130_fd_sc_hd__inv_2 _04344_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].singles[0].s.c ),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_2 _04345_ (.A(\slice.configuroni.mem_ctrl ),
    .Y(_00107_));
 sky130_fd_sc_hd__and2_4 _04346_ (.A(set_out_hard),
    .B(_00107_),
    .X(_00089_));
 sky130_fd_sc_hd__a21o_4 _04347_ (.A1(set_out_hard),
    .A2(_00107_),
    .B1(clb_south_in[8]),
    .X(_00000_));
 sky130_fd_sc_hd__xor2_4 _04348_ (.A(carry_in),
    .B(\slice.sliceluroni.cc.P[0] ),
    .X(_00096_));
 sky130_fd_sc_hd__xor2_4 _04349_ (.A(_00097_),
    .B(\slice.sliceluroni.cc.P[1] ),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_4 _04350_ (.A(_00099_),
    .B(\slice.sliceluroni.cc.P[2] ),
    .X(_00100_));
 sky130_fd_sc_hd__xor2_4 _04351_ (.A(_00101_),
    .B(\slice.sliceluroni.cc.P[3] ),
    .X(_00102_));
 sky130_fd_sc_hd__inv_2 _04352_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0e0.c ),
    .Y(_00040_));
 sky130_fd_sc_hd__inv_2 _04353_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1s0.c ),
    .Y(_00038_));
 sky130_fd_sc_hd__inv_2 _04354_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1w1.c ),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _04355_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0n1.c ),
    .Y(_00047_));
 sky130_fd_sc_hd__inv_2 _04356_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0s0.c ),
    .Y(_00041_));
 sky130_fd_sc_hd__inv_2 _04357_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1w1.c ),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _04358_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1n1.c ),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_2 _04359_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0e0.c ),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _04360_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.n1e1.c ),
    .Y(_00042_));
 sky130_fd_sc_hd__inv_2 _04361_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.e0s1.c ),
    .Y(_00037_));
 sky130_fd_sc_hd__inv_2 _04362_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.s0w0.c ),
    .Y(_00043_));
 sky130_fd_sc_hd__inv_2 _04363_ (.A(\sb.switcharoni.susb.switch_box_element_two[1].elem.w1n0.c ),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_2 _04364_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0e0.c ),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _04365_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1s0.c ),
    .Y(_00026_));
 sky130_fd_sc_hd__inv_2 _04366_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1w1.c ),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_2 _04367_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0n1.c ),
    .Y(_00035_));
 sky130_fd_sc_hd__inv_2 _04368_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0s0.c ),
    .Y(_00029_));
 sky130_fd_sc_hd__inv_2 _04369_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1w1.c ),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _04370_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1n1.c ),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_2 _04371_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0e0.c ),
    .Y(_00034_));
 sky130_fd_sc_hd__inv_2 _04372_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.n1e1.c ),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _04373_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.e0s1.c ),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_2 _04374_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.s0w0.c ),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _04375_ (.A(\sb.switcharoni.susb.switch_box_element_two[0].elem.w1n0.c ),
    .Y(_00036_));
 sky130_fd_sc_hd__inv_2 _04376_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0e0.c ),
    .Y(_00016_));
 sky130_fd_sc_hd__inv_2 _04377_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1s0.c ),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _04378_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1w1.c ),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _04379_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0n1.c ),
    .Y(_00023_));
 sky130_fd_sc_hd__inv_2 _04380_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0s0.c ),
    .Y(_00017_));
 sky130_fd_sc_hd__inv_2 _04381_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1w1.c ),
    .Y(_00015_));
 sky130_fd_sc_hd__inv_2 _04382_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1n1.c ),
    .Y(_00020_));
 sky130_fd_sc_hd__inv_2 _04383_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0e0.c ),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_2 _04384_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n1e1.c ),
    .Y(_00018_));
 sky130_fd_sc_hd__inv_2 _04385_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e0s1.c ),
    .Y(_00013_));
 sky130_fd_sc_hd__inv_2 _04386_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s0w0.c ),
    .Y(_00019_));
 sky130_fd_sc_hd__inv_2 _04387_ (.A(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w1n0.c ),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_2 _04388_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0e0.c ),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _04389_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1s0.c ),
    .Y(_00002_));
 sky130_fd_sc_hd__inv_2 _04390_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1w1.c ),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _04391_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0n1.c ),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _04392_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0s0.c ),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _04393_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1w1.c ),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_2 _04394_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1n1.c ),
    .Y(_00008_));
 sky130_fd_sc_hd__inv_2 _04395_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0e0.c ),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _04396_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n1e1.c ),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _04397_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e0s1.c ),
    .Y(_00001_));
 sky130_fd_sc_hd__inv_2 _04398_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s0w0.c ),
    .Y(_00007_));
 sky130_fd_sc_hd__inv_2 _04399_ (.A(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w1n0.c ),
    .Y(_00012_));
 sky130_fd_sc_hd__and2_4 _04400_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00103_),
    .X(_00108_));
 sky130_fd_sc_hd__buf_2 _04401_ (.A(_00108_),
    .X(_04151_));
 sky130_fd_sc_hd__inv_2 _04402_ (.A(_04151_),
    .Y(_00064_));
 sky130_fd_sc_hd__inv_2 _04403_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .Y(_00109_));
 sky130_fd_sc_hd__and2_4 _04404_ (.A(_00109_),
    .B(_00103_),
    .X(_04150_));
 sky130_fd_sc_hd__inv_2 _04405_ (.A(_00103_),
    .Y(_00110_));
 sky130_fd_sc_hd__or2_4 _04406_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00110_),
    .X(_00063_));
 sky130_fd_sc_hd__and2_4 _04407_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00110_),
    .X(_04149_));
 sky130_fd_sc_hd__or2_4 _04408_ (.A(_00109_),
    .B(_00103_),
    .X(_00062_));
 sky130_fd_sc_hd__or2_4 _04409_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00103_),
    .X(_00111_));
 sky130_fd_sc_hd__buf_2 _04410_ (.A(_00111_),
    .X(_00061_));
 sky130_fd_sc_hd__inv_2 _04411_ (.A(_00061_),
    .Y(_04148_));
 sky130_fd_sc_hd__and2_4 _04412_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00112_));
 sky130_fd_sc_hd__buf_2 _04413_ (.A(_00112_),
    .X(_04127_));
 sky130_fd_sc_hd__inv_2 _04414_ (.A(_04127_),
    .Y(_00060_));
 sky130_fd_sc_hd__inv_2 _04415_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .Y(_00113_));
 sky130_fd_sc_hd__and2_4 _04416_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(_00113_),
    .X(_04126_));
 sky130_fd_sc_hd__inv_2 _04417_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .Y(_00114_));
 sky130_fd_sc_hd__or2_4 _04418_ (.A(_00114_),
    .B(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00059_));
 sky130_fd_sc_hd__and2_4 _04419_ (.A(_00114_),
    .B(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_04125_));
 sky130_fd_sc_hd__or2_4 _04420_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(_00113_),
    .X(_00058_));
 sky130_fd_sc_hd__or2_4 _04421_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00115_));
 sky130_fd_sc_hd__buf_2 _04422_ (.A(_00115_),
    .X(_00057_));
 sky130_fd_sc_hd__inv_2 _04423_ (.A(_00057_),
    .Y(_04124_));
 sky130_fd_sc_hd__and2_4 _04424_ (.A(clb_south_in[2]),
    .B(_00104_),
    .X(_00116_));
 sky130_fd_sc_hd__buf_2 _04425_ (.A(_00116_),
    .X(_04200_));
 sky130_fd_sc_hd__inv_2 _04426_ (.A(_04200_),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_2 _04427_ (.A(clb_south_in[2]),
    .Y(_00117_));
 sky130_fd_sc_hd__and2_4 _04428_ (.A(_00117_),
    .B(_00104_),
    .X(_04199_));
 sky130_fd_sc_hd__inv_2 _04429_ (.A(_00104_),
    .Y(_00118_));
 sky130_fd_sc_hd__or2_4 _04430_ (.A(clb_south_in[2]),
    .B(_00118_),
    .X(_00071_));
 sky130_fd_sc_hd__and2_4 _04431_ (.A(clb_south_in[2]),
    .B(_00118_),
    .X(_04198_));
 sky130_fd_sc_hd__or2_4 _04432_ (.A(_00117_),
    .B(_00104_),
    .X(_00070_));
 sky130_fd_sc_hd__or2_4 _04433_ (.A(clb_south_in[2]),
    .B(_00104_),
    .X(_00119_));
 sky130_fd_sc_hd__buf_2 _04434_ (.A(_00119_),
    .X(_00069_));
 sky130_fd_sc_hd__inv_2 _04435_ (.A(_00069_),
    .Y(_04197_));
 sky130_fd_sc_hd__and2_4 _04436_ (.A(clb_south_in[7]),
    .B(clb_south_in[6]),
    .X(_00120_));
 sky130_fd_sc_hd__buf_2 _04437_ (.A(_00120_),
    .X(_04176_));
 sky130_fd_sc_hd__inv_2 _04438_ (.A(_04176_),
    .Y(_00068_));
 sky130_fd_sc_hd__inv_2 _04439_ (.A(clb_south_in[6]),
    .Y(_00121_));
 sky130_fd_sc_hd__and2_4 _04440_ (.A(clb_south_in[7]),
    .B(_00121_),
    .X(_04175_));
 sky130_fd_sc_hd__inv_2 _04441_ (.A(clb_south_in[7]),
    .Y(_00122_));
 sky130_fd_sc_hd__or2_4 _04442_ (.A(_00122_),
    .B(clb_south_in[6]),
    .X(_00067_));
 sky130_fd_sc_hd__and2_4 _04443_ (.A(_00122_),
    .B(clb_south_in[6]),
    .X(_04174_));
 sky130_fd_sc_hd__or2_4 _04444_ (.A(clb_south_in[7]),
    .B(_00121_),
    .X(_00066_));
 sky130_fd_sc_hd__or2_4 _04445_ (.A(clb_south_in[7]),
    .B(clb_south_in[6]),
    .X(_00123_));
 sky130_fd_sc_hd__buf_2 _04446_ (.A(_00123_),
    .X(_00065_));
 sky130_fd_sc_hd__inv_2 _04447_ (.A(_00065_),
    .Y(_04173_));
 sky130_fd_sc_hd__and2_4 _04448_ (.A(clb_west_in[2]),
    .B(_00105_),
    .X(_00124_));
 sky130_fd_sc_hd__buf_2 _04449_ (.A(_00124_),
    .X(_04249_));
 sky130_fd_sc_hd__inv_2 _04450_ (.A(_04249_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _04451_ (.A(clb_west_in[2]),
    .Y(_00125_));
 sky130_fd_sc_hd__and2_4 _04452_ (.A(_00125_),
    .B(_00105_),
    .X(_04248_));
 sky130_fd_sc_hd__inv_2 _04453_ (.A(_00105_),
    .Y(_00126_));
 sky130_fd_sc_hd__or2_4 _04454_ (.A(clb_west_in[2]),
    .B(_00126_),
    .X(_00079_));
 sky130_fd_sc_hd__and2_4 _04455_ (.A(clb_west_in[2]),
    .B(_00126_),
    .X(_04247_));
 sky130_fd_sc_hd__or2_4 _04456_ (.A(_00125_),
    .B(_00105_),
    .X(_00078_));
 sky130_fd_sc_hd__or2_4 _04457_ (.A(clb_west_in[2]),
    .B(_00105_),
    .X(_00127_));
 sky130_fd_sc_hd__buf_2 _04458_ (.A(_00127_),
    .X(_00077_));
 sky130_fd_sc_hd__inv_2 _04459_ (.A(_00077_),
    .Y(_04246_));
 sky130_fd_sc_hd__and2_4 _04460_ (.A(clb_west_in[7]),
    .B(clb_west_in[6]),
    .X(_00128_));
 sky130_fd_sc_hd__buf_2 _04461_ (.A(_00128_),
    .X(_04225_));
 sky130_fd_sc_hd__inv_2 _04462_ (.A(_04225_),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _04463_ (.A(clb_west_in[6]),
    .Y(_00129_));
 sky130_fd_sc_hd__and2_4 _04464_ (.A(clb_west_in[7]),
    .B(_00129_),
    .X(_04224_));
 sky130_fd_sc_hd__inv_2 _04465_ (.A(clb_west_in[7]),
    .Y(_00130_));
 sky130_fd_sc_hd__or2_4 _04466_ (.A(_00130_),
    .B(clb_west_in[6]),
    .X(_00075_));
 sky130_fd_sc_hd__and2_4 _04467_ (.A(_00130_),
    .B(clb_west_in[6]),
    .X(_04223_));
 sky130_fd_sc_hd__or2_4 _04468_ (.A(clb_west_in[7]),
    .B(_00129_),
    .X(_00074_));
 sky130_fd_sc_hd__or2_4 _04469_ (.A(clb_west_in[7]),
    .B(clb_west_in[6]),
    .X(_00131_));
 sky130_fd_sc_hd__buf_2 _04470_ (.A(_00131_),
    .X(_00073_));
 sky130_fd_sc_hd__inv_2 _04471_ (.A(_00073_),
    .Y(_04222_));
 sky130_fd_sc_hd__and2_4 _04472_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00106_),
    .X(_00132_));
 sky130_fd_sc_hd__buf_2 _04473_ (.A(_00132_),
    .X(_04298_));
 sky130_fd_sc_hd__inv_2 _04474_ (.A(_04298_),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_2 _04475_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .Y(_00133_));
 sky130_fd_sc_hd__and2_4 _04476_ (.A(_00133_),
    .B(_00106_),
    .X(_04297_));
 sky130_fd_sc_hd__inv_2 _04477_ (.A(_00106_),
    .Y(_00134_));
 sky130_fd_sc_hd__or2_4 _04478_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00134_),
    .X(_00087_));
 sky130_fd_sc_hd__and2_4 _04479_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00134_),
    .X(_04296_));
 sky130_fd_sc_hd__or2_4 _04480_ (.A(_00133_),
    .B(_00106_),
    .X(_00086_));
 sky130_fd_sc_hd__or2_4 _04481_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ),
    .B(_00106_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_2 _04482_ (.A(_00135_),
    .X(_00085_));
 sky130_fd_sc_hd__inv_2 _04483_ (.A(_00085_),
    .Y(_04295_));
 sky130_fd_sc_hd__and2_4 _04484_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00136_));
 sky130_fd_sc_hd__buf_2 _04485_ (.A(_00136_),
    .X(_04274_));
 sky130_fd_sc_hd__inv_2 _04486_ (.A(_04274_),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_2 _04487_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .Y(_00137_));
 sky130_fd_sc_hd__and2_4 _04488_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(_00137_),
    .X(_04273_));
 sky130_fd_sc_hd__inv_2 _04489_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .Y(_00138_));
 sky130_fd_sc_hd__or2_4 _04490_ (.A(_00138_),
    .B(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00083_));
 sky130_fd_sc_hd__and2_4 _04491_ (.A(_00138_),
    .B(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_04272_));
 sky130_fd_sc_hd__or2_4 _04492_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(_00137_),
    .X(_00082_));
 sky130_fd_sc_hd__or2_4 _04493_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ),
    .B(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ),
    .X(_00139_));
 sky130_fd_sc_hd__buf_2 _04494_ (.A(_00139_),
    .X(_00081_));
 sky130_fd_sc_hd__inv_2 _04495_ (.A(_00081_),
    .Y(_04271_));
 sky130_fd_sc_hd__inv_2 _04496_ (.A(set_in_hard),
    .Y(_00140_));
 sky130_fd_sc_hd__and2_4 _04497_ (.A(cen),
    .B(_00140_),
    .X(\slice.configuroni.comb_shifter.head_bit.shift_enable ));
 sky130_fd_sc_hd__inv_2 _04498_ (.A(set_out_hard),
    .Y(_00141_));
 sky130_fd_sc_hd__and2_4 _04499_ (.A(_00141_),
    .B(cen),
    .X(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ));
 sky130_fd_sc_hd__inv_2 _04500_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[2].s.c ),
    .Y(_00686_));
 sky130_fd_sc_hd__inv_2 _04501_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[1].s.c ),
    .Y(_00687_));
 sky130_fd_sc_hd__inv_2 _04502_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[0].s.c ),
    .Y(_00688_));
 sky130_fd_sc_hd__inv_2 _04503_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].singles[3].s.c ),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_2 _04504_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].singles[2].s.c ),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _04505_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].singles[1].s.c ),
    .Y(_00691_));
 sky130_fd_sc_hd__inv_2 _04506_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].singles[0].s.c ),
    .Y(_00692_));
 sky130_fd_sc_hd__inv_2 _04507_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[4].s.c ),
    .Y(_00693_));
 sky130_fd_sc_hd__inv_2 _04508_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[3].s.c ),
    .Y(_00694_));
 sky130_fd_sc_hd__inv_2 _04509_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[2].s.c ),
    .Y(_00695_));
 sky130_fd_sc_hd__inv_2 _04510_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[1].s.c ),
    .Y(_00696_));
 sky130_fd_sc_hd__inv_2 _04511_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.c ),
    .Y(_00697_));
 sky130_fd_sc_hd__inv_2 _04512_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[7].s.c ),
    .Y(_00698_));
 sky130_fd_sc_hd__inv_2 _04513_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[6].s.c ),
    .Y(_00699_));
 sky130_fd_sc_hd__inv_2 _04514_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[5].s.c ),
    .Y(_00700_));
 sky130_fd_sc_hd__inv_2 _04515_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[4].s.c ),
    .Y(_00701_));
 sky130_fd_sc_hd__inv_2 _04516_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[3].s.c ),
    .Y(_00702_));
 sky130_fd_sc_hd__inv_2 _04517_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[2].s.c ),
    .Y(_00703_));
 sky130_fd_sc_hd__inv_2 _04518_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[1].s.c ),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _04519_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[0].s.c ),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _04520_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].singles[3].s.c ),
    .Y(_00706_));
 sky130_fd_sc_hd__inv_2 _04521_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].singles[2].s.c ),
    .Y(_00707_));
 sky130_fd_sc_hd__inv_2 _04522_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].singles[1].s.c ),
    .Y(_00708_));
 sky130_fd_sc_hd__inv_2 _04523_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].singles[0].s.c ),
    .Y(_00709_));
 sky130_fd_sc_hd__inv_2 _04524_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[4].s.c ),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _04525_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[3].s.c ),
    .Y(_00711_));
 sky130_fd_sc_hd__inv_2 _04526_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[2].s.c ),
    .Y(_00712_));
 sky130_fd_sc_hd__inv_2 _04527_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[1].s.c ),
    .Y(_00713_));
 sky130_fd_sc_hd__inv_2 _04528_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.c ),
    .Y(_00714_));
 sky130_fd_sc_hd__inv_2 _04529_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[7].s.c ),
    .Y(_00715_));
 sky130_fd_sc_hd__inv_2 _04530_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[6].s.c ),
    .Y(_00716_));
 sky130_fd_sc_hd__inv_2 _04531_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[5].s.c ),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _04532_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[4].s.c ),
    .Y(_00718_));
 sky130_fd_sc_hd__inv_2 _04533_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[3].s.c ),
    .Y(_00719_));
 sky130_fd_sc_hd__inv_2 _04534_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[2].s.c ),
    .Y(_00720_));
 sky130_fd_sc_hd__inv_2 _04535_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[1].s.c ),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _04536_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[0].s.c ),
    .Y(_00722_));
 sky130_fd_sc_hd__inv_2 _04537_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].singles[3].s.c ),
    .Y(_00723_));
 sky130_fd_sc_hd__inv_2 _04538_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].singles[2].s.c ),
    .Y(_00724_));
 sky130_fd_sc_hd__inv_2 _04539_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].singles[1].s.c ),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _04540_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].singles[0].s.c ),
    .Y(_00726_));
 sky130_fd_sc_hd__inv_2 _04541_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[4].s.c ),
    .Y(_00727_));
 sky130_fd_sc_hd__inv_2 _04542_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[3].s.c ),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _04543_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[2].s.c ),
    .Y(_00729_));
 sky130_fd_sc_hd__inv_2 _04544_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[1].s.c ),
    .Y(_00730_));
 sky130_fd_sc_hd__inv_2 _04545_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.c ),
    .Y(_00731_));
 sky130_fd_sc_hd__inv_2 _04546_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[7].s.c ),
    .Y(_00732_));
 sky130_fd_sc_hd__inv_2 _04547_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[6].s.c ),
    .Y(_00733_));
 sky130_fd_sc_hd__inv_2 _04548_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[5].s.c ),
    .Y(_00734_));
 sky130_fd_sc_hd__inv_2 _04549_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[4].s.c ),
    .Y(_00735_));
 sky130_fd_sc_hd__inv_2 _04550_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[3].s.c ),
    .Y(_00736_));
 sky130_fd_sc_hd__inv_2 _04551_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[2].s.c ),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _04552_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[1].s.c ),
    .Y(_00738_));
 sky130_fd_sc_hd__inv_2 _04553_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[0].s.c ),
    .Y(_00739_));
 sky130_fd_sc_hd__inv_2 _04554_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].singles[3].s.c ),
    .Y(_00740_));
 sky130_fd_sc_hd__inv_2 _04555_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].singles[2].s.c ),
    .Y(_00741_));
 sky130_fd_sc_hd__inv_2 _04556_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].singles[1].s.c ),
    .Y(_00742_));
 sky130_fd_sc_hd__inv_2 _04557_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].singles[0].s.c ),
    .Y(_00743_));
 sky130_fd_sc_hd__inv_2 _04558_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[4].s.c ),
    .Y(_00744_));
 sky130_fd_sc_hd__inv_2 _04559_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[3].s.c ),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _04560_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[2].s.c ),
    .Y(_00746_));
 sky130_fd_sc_hd__inv_2 _04561_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[1].s.c ),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _04562_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.c ),
    .Y(_00748_));
 sky130_fd_sc_hd__inv_2 _04563_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[7].s.c ),
    .Y(_00749_));
 sky130_fd_sc_hd__inv_2 _04564_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[6].s.c ),
    .Y(_00750_));
 sky130_fd_sc_hd__inv_2 _04565_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[5].s.c ),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_2 _04566_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[4].s.c ),
    .Y(_00752_));
 sky130_fd_sc_hd__inv_2 _04567_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[3].s.c ),
    .Y(_00753_));
 sky130_fd_sc_hd__inv_2 _04568_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[2].s.c ),
    .Y(_00754_));
 sky130_fd_sc_hd__inv_2 _04569_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[1].s.c ),
    .Y(_00755_));
 sky130_fd_sc_hd__inv_2 _04570_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[0].s.c ),
    .Y(_00756_));
 sky130_fd_sc_hd__inv_2 _04571_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].singles[3].s.c ),
    .Y(_00757_));
 sky130_fd_sc_hd__inv_2 _04572_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].singles[2].s.c ),
    .Y(_00758_));
 sky130_fd_sc_hd__inv_2 _04573_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].singles[1].s.c ),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_2 _04574_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].singles[0].s.c ),
    .Y(_00760_));
 sky130_fd_sc_hd__inv_2 _04575_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[4].s.c ),
    .Y(_00761_));
 sky130_fd_sc_hd__inv_2 _04576_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[3].s.c ),
    .Y(_00762_));
 sky130_fd_sc_hd__inv_2 _04577_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[2].s.c ),
    .Y(_00763_));
 sky130_fd_sc_hd__inv_2 _04578_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[1].s.c ),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_2 _04579_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.c ),
    .Y(_00765_));
 sky130_fd_sc_hd__inv_2 _04580_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[7].s.c ),
    .Y(_00766_));
 sky130_fd_sc_hd__inv_2 _04581_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[6].s.c ),
    .Y(_00767_));
 sky130_fd_sc_hd__inv_2 _04582_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[5].s.c ),
    .Y(_00768_));
 sky130_fd_sc_hd__inv_2 _04583_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[4].s.c ),
    .Y(_00769_));
 sky130_fd_sc_hd__inv_2 _04584_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[3].s.c ),
    .Y(_00770_));
 sky130_fd_sc_hd__inv_2 _04585_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[2].s.c ),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_2 _04586_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[1].s.c ),
    .Y(_00772_));
 sky130_fd_sc_hd__inv_2 _04587_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[0].s.c ),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _04588_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].singles[3].s.c ),
    .Y(_00774_));
 sky130_fd_sc_hd__inv_2 _04589_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].singles[2].s.c ),
    .Y(_00775_));
 sky130_fd_sc_hd__inv_2 _04590_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].singles[1].s.c ),
    .Y(_00776_));
 sky130_fd_sc_hd__inv_2 _04591_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].singles[0].s.c ),
    .Y(_00777_));
 sky130_fd_sc_hd__inv_2 _04592_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[4].s.c ),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _04593_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[3].s.c ),
    .Y(_00779_));
 sky130_fd_sc_hd__inv_2 _04594_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[2].s.c ),
    .Y(_00780_));
 sky130_fd_sc_hd__inv_2 _04595_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[1].s.c ),
    .Y(_00781_));
 sky130_fd_sc_hd__inv_2 _04596_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.c ),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _04597_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[7].s.c ),
    .Y(_00783_));
 sky130_fd_sc_hd__inv_2 _04598_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[6].s.c ),
    .Y(_00784_));
 sky130_fd_sc_hd__inv_2 _04599_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[5].s.c ),
    .Y(_00785_));
 sky130_fd_sc_hd__inv_2 _04600_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[4].s.c ),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _04601_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[3].s.c ),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _04602_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[2].s.c ),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _04603_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[1].s.c ),
    .Y(_00789_));
 sky130_fd_sc_hd__inv_2 _04604_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[0].s.c ),
    .Y(_00790_));
 sky130_fd_sc_hd__inv_2 _04605_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].singles[3].s.c ),
    .Y(_00791_));
 sky130_fd_sc_hd__inv_2 _04606_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].singles[2].s.c ),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_2 _04607_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].singles[1].s.c ),
    .Y(_00793_));
 sky130_fd_sc_hd__inv_2 _04608_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].singles[0].s.c ),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _04609_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[4].s.c ),
    .Y(_00795_));
 sky130_fd_sc_hd__inv_2 _04610_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[3].s.c ),
    .Y(_00796_));
 sky130_fd_sc_hd__inv_2 _04611_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[2].s.c ),
    .Y(_00797_));
 sky130_fd_sc_hd__inv_2 _04612_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[1].s.c ),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _04613_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.c ),
    .Y(_00799_));
 sky130_fd_sc_hd__inv_2 _04614_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[7].s.c ),
    .Y(_00800_));
 sky130_fd_sc_hd__inv_2 _04615_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[6].s.c ),
    .Y(_00801_));
 sky130_fd_sc_hd__inv_2 _04616_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[5].s.c ),
    .Y(_00802_));
 sky130_fd_sc_hd__inv_2 _04617_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[4].s.c ),
    .Y(_00803_));
 sky130_fd_sc_hd__inv_2 _04618_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[3].s.c ),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _04619_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[2].s.c ),
    .Y(_00805_));
 sky130_fd_sc_hd__inv_2 _04620_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[1].s.c ),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _04621_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[0].s.c ),
    .Y(_00807_));
 sky130_fd_sc_hd__inv_2 _04622_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].singles[3].s.c ),
    .Y(_00808_));
 sky130_fd_sc_hd__inv_2 _04623_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].singles[2].s.c ),
    .Y(_00809_));
 sky130_fd_sc_hd__inv_2 _04624_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].singles[1].s.c ),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_2 _04625_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[4].s.c ),
    .Y(_00610_));
 sky130_fd_sc_hd__inv_2 _04626_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[3].s.c ),
    .Y(_00616_));
 sky130_fd_sc_hd__inv_2 _04627_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[2].s.c ),
    .Y(_00622_));
 sky130_fd_sc_hd__inv_2 _04628_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[1].s.c ),
    .Y(_00628_));
 sky130_fd_sc_hd__inv_2 _04629_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[0].s.c ),
    .Y(_00634_));
 sky130_fd_sc_hd__inv_2 _04630_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].singles[3].s.c ),
    .Y(_00640_));
 sky130_fd_sc_hd__inv_2 _04631_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].singles[2].s.c ),
    .Y(_00646_));
 sky130_fd_sc_hd__inv_2 _04632_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].singles[1].s.c ),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_2 _04633_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[3].s.c ),
    .Y(_00611_));
 sky130_fd_sc_hd__inv_2 _04634_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[2].s.c ),
    .Y(_00617_));
 sky130_fd_sc_hd__inv_2 _04635_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[1].s.c ),
    .Y(_00623_));
 sky130_fd_sc_hd__inv_2 _04636_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[0].s.c ),
    .Y(_00629_));
 sky130_fd_sc_hd__inv_2 _04637_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].singles[3].s.c ),
    .Y(_00635_));
 sky130_fd_sc_hd__inv_2 _04638_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].singles[2].s.c ),
    .Y(_00641_));
 sky130_fd_sc_hd__inv_2 _04639_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].singles[1].s.c ),
    .Y(_00647_));
 sky130_fd_sc_hd__inv_2 _04640_ (.A(\cb_east.inst.connectaroni.clb0_outputs[4].singles[0].s.c ),
    .Y(_00653_));
 sky130_fd_sc_hd__inv_2 _04641_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[3].s.c ),
    .Y(_00612_));
 sky130_fd_sc_hd__inv_2 _04642_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[2].s.c ),
    .Y(_00618_));
 sky130_fd_sc_hd__inv_2 _04643_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[1].s.c ),
    .Y(_00624_));
 sky130_fd_sc_hd__inv_2 _04644_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.c ),
    .Y(_00630_));
 sky130_fd_sc_hd__inv_2 _04645_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].singles[3].s.c ),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _04646_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].singles[2].s.c ),
    .Y(_00642_));
 sky130_fd_sc_hd__inv_2 _04647_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].singles[1].s.c ),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _04648_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].singles[0].s.c ),
    .Y(_00654_));
 sky130_fd_sc_hd__inv_2 _04649_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[3].s.c ),
    .Y(_00613_));
 sky130_fd_sc_hd__inv_2 _04650_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[2].s.c ),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _04651_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[1].s.c ),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _04652_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.c ),
    .Y(_00631_));
 sky130_fd_sc_hd__inv_2 _04653_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].singles[3].s.c ),
    .Y(_00637_));
 sky130_fd_sc_hd__inv_2 _04654_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].singles[2].s.c ),
    .Y(_00643_));
 sky130_fd_sc_hd__inv_2 _04655_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].singles[1].s.c ),
    .Y(_00649_));
 sky130_fd_sc_hd__inv_2 _04656_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].singles[0].s.c ),
    .Y(_00655_));
 sky130_fd_sc_hd__inv_2 _04657_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[3].s.c ),
    .Y(_00614_));
 sky130_fd_sc_hd__inv_2 _04658_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[2].s.c ),
    .Y(_00620_));
 sky130_fd_sc_hd__inv_2 _04659_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[1].s.c ),
    .Y(_00626_));
 sky130_fd_sc_hd__inv_2 _04660_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.c ),
    .Y(_00632_));
 sky130_fd_sc_hd__inv_2 _04661_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].singles[3].s.c ),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _04662_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].singles[2].s.c ),
    .Y(_00644_));
 sky130_fd_sc_hd__inv_2 _04663_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].singles[1].s.c ),
    .Y(_00650_));
 sky130_fd_sc_hd__inv_2 _04664_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].singles[0].s.c ),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_2 _04665_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].singles[0].s.c ),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _04666_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].directs[4].s.c ),
    .Y(_00812_));
 sky130_fd_sc_hd__inv_2 _04667_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].directs[3].s.c ),
    .Y(_00813_));
 sky130_fd_sc_hd__inv_2 _04668_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].directs[2].s.c ),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _04669_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].directs[1].s.c ),
    .Y(_00815_));
 sky130_fd_sc_hd__inv_2 _04670_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.c ),
    .Y(_00816_));
 sky130_fd_sc_hd__inv_2 _04671_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[7].s.c ),
    .Y(_00817_));
 sky130_fd_sc_hd__inv_2 _04672_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[6].s.c ),
    .Y(_00818_));
 sky130_fd_sc_hd__inv_2 _04673_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[5].s.c ),
    .Y(_00819_));
 sky130_fd_sc_hd__inv_2 _04674_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[4].s.c ),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _04675_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[3].s.c ),
    .Y(_00821_));
 sky130_fd_sc_hd__inv_2 _04676_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[2].s.c ),
    .Y(_00822_));
 sky130_fd_sc_hd__inv_2 _04677_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[1].s.c ),
    .Y(_00823_));
 sky130_fd_sc_hd__inv_2 _04678_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[0].s.c ),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _04679_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].singles[3].s.c ),
    .Y(_00825_));
 sky130_fd_sc_hd__inv_2 _04680_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].singles[2].s.c ),
    .Y(_00826_));
 sky130_fd_sc_hd__inv_2 _04681_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].singles[1].s.c ),
    .Y(_00827_));
 sky130_fd_sc_hd__inv_2 _04682_ (.A(\cb_east.inst.connectaroni.clb0_inputs[9].singles[0].s.c ),
    .Y(_00828_));
 sky130_fd_sc_hd__inv_2 _04683_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].directs[4].s.c ),
    .Y(_00829_));
 sky130_fd_sc_hd__inv_2 _04684_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].directs[3].s.c ),
    .Y(_00830_));
 sky130_fd_sc_hd__inv_2 _04685_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].directs[2].s.c ),
    .Y(_00831_));
 sky130_fd_sc_hd__inv_2 _04686_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].directs[1].s.c ),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _04687_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.c ),
    .Y(_00833_));
 sky130_fd_sc_hd__inv_2 _04688_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[7].s.c ),
    .Y(_00834_));
 sky130_fd_sc_hd__inv_2 _04689_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[6].s.c ),
    .Y(_00835_));
 sky130_fd_sc_hd__inv_2 _04690_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[5].s.c ),
    .Y(_00836_));
 sky130_fd_sc_hd__inv_2 _04691_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[4].s.c ),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _04692_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[3].s.c ),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _04693_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[2].s.c ),
    .Y(_00839_));
 sky130_fd_sc_hd__inv_2 _04694_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[1].s.c ),
    .Y(_00840_));
 sky130_fd_sc_hd__inv_2 _04695_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[0].s.c ),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _04696_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].singles[3].s.c ),
    .Y(_00842_));
 sky130_fd_sc_hd__inv_2 _04697_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].singles[2].s.c ),
    .Y(_00843_));
 sky130_fd_sc_hd__inv_2 _04698_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].singles[1].s.c ),
    .Y(_00844_));
 sky130_fd_sc_hd__inv_2 _04699_ (.A(\cb_east.inst.connectaroni.clb0_inputs[8].singles[0].s.c ),
    .Y(_00845_));
 sky130_fd_sc_hd__inv_2 _04700_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[4].s.c ),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _04701_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[3].s.c ),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _04702_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[2].s.c ),
    .Y(_00848_));
 sky130_fd_sc_hd__inv_2 _04703_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[1].s.c ),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _04704_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.c ),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _04705_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[7].s.c ),
    .Y(_00851_));
 sky130_fd_sc_hd__inv_2 _04706_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[6].s.c ),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _04707_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[5].s.c ),
    .Y(_00853_));
 sky130_fd_sc_hd__inv_2 _04708_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[4].s.c ),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _04709_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[3].s.c ),
    .Y(_00855_));
 sky130_fd_sc_hd__inv_2 _04710_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[2].s.c ),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _04711_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[1].s.c ),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _04712_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[0].s.c ),
    .Y(_00858_));
 sky130_fd_sc_hd__inv_2 _04713_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].singles[3].s.c ),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _04714_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].singles[2].s.c ),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _04715_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].singles[1].s.c ),
    .Y(_00861_));
 sky130_fd_sc_hd__inv_2 _04716_ (.A(\cb_east.inst.connectaroni.clb0_inputs[7].singles[0].s.c ),
    .Y(_00862_));
 sky130_fd_sc_hd__inv_2 _04717_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[4].s.c ),
    .Y(_00863_));
 sky130_fd_sc_hd__inv_2 _04718_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[3].s.c ),
    .Y(_00864_));
 sky130_fd_sc_hd__inv_2 _04719_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[2].s.c ),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _04720_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[1].s.c ),
    .Y(_00866_));
 sky130_fd_sc_hd__inv_2 _04721_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.c ),
    .Y(_00867_));
 sky130_fd_sc_hd__inv_2 _04722_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[7].s.c ),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_2 _04723_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[6].s.c ),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _04724_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[5].s.c ),
    .Y(_00870_));
 sky130_fd_sc_hd__inv_2 _04725_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[4].s.c ),
    .Y(_00871_));
 sky130_fd_sc_hd__inv_2 _04726_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[3].s.c ),
    .Y(_00872_));
 sky130_fd_sc_hd__inv_2 _04727_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[2].s.c ),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _04728_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[1].s.c ),
    .Y(_00874_));
 sky130_fd_sc_hd__inv_2 _04729_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[0].s.c ),
    .Y(_00875_));
 sky130_fd_sc_hd__inv_2 _04730_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].singles[3].s.c ),
    .Y(_00876_));
 sky130_fd_sc_hd__inv_2 _04731_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].singles[2].s.c ),
    .Y(_00877_));
 sky130_fd_sc_hd__inv_2 _04732_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].singles[1].s.c ),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_2 _04733_ (.A(\cb_east.inst.connectaroni.clb0_inputs[6].singles[0].s.c ),
    .Y(_00879_));
 sky130_fd_sc_hd__inv_2 _04734_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].directs[4].s.c ),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _04735_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].directs[3].s.c ),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _04736_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].directs[2].s.c ),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _04737_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].directs[1].s.c ),
    .Y(_00883_));
 sky130_fd_sc_hd__inv_2 _04738_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.c ),
    .Y(_00884_));
 sky130_fd_sc_hd__inv_2 _04739_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[7].s.c ),
    .Y(_00885_));
 sky130_fd_sc_hd__inv_2 _04740_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[6].s.c ),
    .Y(_00886_));
 sky130_fd_sc_hd__inv_2 _04741_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[5].s.c ),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _04742_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[4].s.c ),
    .Y(_00888_));
 sky130_fd_sc_hd__inv_2 _04743_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[3].s.c ),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _04744_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[2].s.c ),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _04745_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[1].s.c ),
    .Y(_00891_));
 sky130_fd_sc_hd__inv_2 _04746_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[0].s.c ),
    .Y(_00892_));
 sky130_fd_sc_hd__inv_2 _04747_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].singles[3].s.c ),
    .Y(_00893_));
 sky130_fd_sc_hd__inv_2 _04748_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].singles[2].s.c ),
    .Y(_00894_));
 sky130_fd_sc_hd__inv_2 _04749_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].singles[1].s.c ),
    .Y(_00895_));
 sky130_fd_sc_hd__inv_2 _04750_ (.A(\cb_east.inst.connectaroni.clb0_inputs[5].singles[0].s.c ),
    .Y(_00896_));
 sky130_fd_sc_hd__inv_2 _04751_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].directs[4].s.c ),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _04752_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].directs[3].s.c ),
    .Y(_00898_));
 sky130_fd_sc_hd__inv_2 _04753_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].directs[2].s.c ),
    .Y(_00899_));
 sky130_fd_sc_hd__inv_2 _04754_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].directs[1].s.c ),
    .Y(_00900_));
 sky130_fd_sc_hd__inv_2 _04755_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.c ),
    .Y(_00901_));
 sky130_fd_sc_hd__inv_2 _04756_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[7].s.c ),
    .Y(_00902_));
 sky130_fd_sc_hd__inv_2 _04757_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[6].s.c ),
    .Y(_00903_));
 sky130_fd_sc_hd__inv_2 _04758_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[5].s.c ),
    .Y(_00904_));
 sky130_fd_sc_hd__inv_2 _04759_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[4].s.c ),
    .Y(_00905_));
 sky130_fd_sc_hd__inv_2 _04760_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[3].s.c ),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_2 _04761_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[2].s.c ),
    .Y(_00907_));
 sky130_fd_sc_hd__inv_2 _04762_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[1].s.c ),
    .Y(_00908_));
 sky130_fd_sc_hd__inv_2 _04763_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[0].s.c ),
    .Y(_00909_));
 sky130_fd_sc_hd__inv_2 _04764_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].singles[3].s.c ),
    .Y(_00910_));
 sky130_fd_sc_hd__inv_2 _04765_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].singles[2].s.c ),
    .Y(_00911_));
 sky130_fd_sc_hd__inv_2 _04766_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].singles[1].s.c ),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _04767_ (.A(\cb_east.inst.connectaroni.clb0_inputs[4].singles[0].s.c ),
    .Y(_00913_));
 sky130_fd_sc_hd__inv_2 _04768_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].directs[4].s.c ),
    .Y(_00914_));
 sky130_fd_sc_hd__inv_2 _04769_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].directs[3].s.c ),
    .Y(_00915_));
 sky130_fd_sc_hd__inv_2 _04770_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].directs[2].s.c ),
    .Y(_00916_));
 sky130_fd_sc_hd__inv_2 _04771_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].directs[1].s.c ),
    .Y(_00917_));
 sky130_fd_sc_hd__inv_2 _04772_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.c ),
    .Y(_00918_));
 sky130_fd_sc_hd__inv_2 _04773_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[7].s.c ),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _04774_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[6].s.c ),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_2 _04775_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[5].s.c ),
    .Y(_00921_));
 sky130_fd_sc_hd__inv_2 _04776_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[4].s.c ),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _04777_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[3].s.c ),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _04778_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[2].s.c ),
    .Y(_00924_));
 sky130_fd_sc_hd__inv_2 _04779_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[1].s.c ),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _04780_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[0].s.c ),
    .Y(_00926_));
 sky130_fd_sc_hd__inv_2 _04781_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].singles[3].s.c ),
    .Y(_00927_));
 sky130_fd_sc_hd__inv_2 _04782_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].singles[2].s.c ),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _04783_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].singles[1].s.c ),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _04784_ (.A(\cb_east.inst.connectaroni.clb0_inputs[3].singles[0].s.c ),
    .Y(_00930_));
 sky130_fd_sc_hd__inv_2 _04785_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[4].s.c ),
    .Y(_00931_));
 sky130_fd_sc_hd__inv_2 _04786_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[3].s.c ),
    .Y(_00932_));
 sky130_fd_sc_hd__inv_2 _04787_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[2].s.c ),
    .Y(_00933_));
 sky130_fd_sc_hd__inv_2 _04788_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[1].s.c ),
    .Y(_00934_));
 sky130_fd_sc_hd__inv_2 _04789_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.c ),
    .Y(_00935_));
 sky130_fd_sc_hd__inv_2 _04790_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[7].s.c ),
    .Y(_00936_));
 sky130_fd_sc_hd__inv_2 _04791_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[6].s.c ),
    .Y(_00937_));
 sky130_fd_sc_hd__inv_2 _04792_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[5].s.c ),
    .Y(_00938_));
 sky130_fd_sc_hd__inv_2 _04793_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[4].s.c ),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _04794_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[3].s.c ),
    .Y(_00940_));
 sky130_fd_sc_hd__inv_2 _04795_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[2].s.c ),
    .Y(_00941_));
 sky130_fd_sc_hd__inv_2 _04796_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[1].s.c ),
    .Y(_00942_));
 sky130_fd_sc_hd__inv_2 _04797_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[0].s.c ),
    .Y(_00943_));
 sky130_fd_sc_hd__inv_2 _04798_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].singles[3].s.c ),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _04799_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].singles[2].s.c ),
    .Y(_00945_));
 sky130_fd_sc_hd__inv_2 _04800_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].singles[1].s.c ),
    .Y(_00946_));
 sky130_fd_sc_hd__inv_2 _04801_ (.A(\cb_east.inst.connectaroni.clb0_inputs[2].singles[0].s.c ),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _04802_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].directs[4].s.c ),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _04803_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].directs[3].s.c ),
    .Y(_00949_));
 sky130_fd_sc_hd__inv_2 _04804_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].directs[2].s.c ),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_2 _04805_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].directs[1].s.c ),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _04806_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.c ),
    .Y(_00952_));
 sky130_fd_sc_hd__inv_2 _04807_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[7].s.c ),
    .Y(_00953_));
 sky130_fd_sc_hd__inv_2 _04808_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[6].s.c ),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _04809_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[5].s.c ),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _04810_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[4].s.c ),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _04811_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[3].s.c ),
    .Y(_00957_));
 sky130_fd_sc_hd__inv_2 _04812_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[2].s.c ),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _04813_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[1].s.c ),
    .Y(_00959_));
 sky130_fd_sc_hd__inv_2 _04814_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[0].s.c ),
    .Y(_00960_));
 sky130_fd_sc_hd__inv_2 _04815_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].singles[3].s.c ),
    .Y(_00961_));
 sky130_fd_sc_hd__inv_2 _04816_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].singles[2].s.c ),
    .Y(_00962_));
 sky130_fd_sc_hd__inv_2 _04817_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].singles[1].s.c ),
    .Y(_00963_));
 sky130_fd_sc_hd__inv_2 _04818_ (.A(\cb_east.inst.connectaroni.clb0_inputs[1].singles[0].s.c ),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _04819_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].directs[4].s.c ),
    .Y(_00965_));
 sky130_fd_sc_hd__inv_2 _04820_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].directs[3].s.c ),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _04821_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].directs[2].s.c ),
    .Y(_00967_));
 sky130_fd_sc_hd__inv_2 _04822_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].directs[1].s.c ),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _04823_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.c ),
    .Y(_00969_));
 sky130_fd_sc_hd__inv_2 _04824_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[7].s.c ),
    .Y(_00970_));
 sky130_fd_sc_hd__inv_2 _04825_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[6].s.c ),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _04826_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[5].s.c ),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _04827_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[4].s.c ),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _04828_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[3].s.c ),
    .Y(_00974_));
 sky130_fd_sc_hd__inv_2 _04829_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[2].s.c ),
    .Y(_00975_));
 sky130_fd_sc_hd__inv_2 _04830_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[1].s.c ),
    .Y(_00976_));
 sky130_fd_sc_hd__inv_2 _04831_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[0].s.c ),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_2 _04832_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].singles[3].s.c ),
    .Y(_00978_));
 sky130_fd_sc_hd__inv_2 _04833_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].singles[2].s.c ),
    .Y(_00979_));
 sky130_fd_sc_hd__inv_2 _04834_ (.A(\cb_east.inst.connectaroni.clb0_inputs[0].singles[1].s.c ),
    .Y(_00980_));
 sky130_fd_sc_hd__inv_2 _04835_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[3].s.c ),
    .Y(_00142_));
 sky130_fd_sc_hd__inv_2 _04836_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[2].s.c ),
    .Y(_00143_));
 sky130_fd_sc_hd__inv_2 _04837_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[1].s.c ),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _04838_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[0].s.c ),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _04839_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].singles[3].s.c ),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _04840_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].singles[2].s.c ),
    .Y(_00147_));
 sky130_fd_sc_hd__inv_2 _04841_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].singles[1].s.c ),
    .Y(_00148_));
 sky130_fd_sc_hd__inv_2 _04842_ (.A(\cb_north.inst.connectaroni.clb1_outputs[4].singles[0].s.c ),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _04843_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[3].s.c ),
    .Y(_00150_));
 sky130_fd_sc_hd__inv_2 _04844_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[2].s.c ),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _04845_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[1].s.c ),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _04846_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[0].s.c ),
    .Y(_00153_));
 sky130_fd_sc_hd__inv_2 _04847_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].singles[3].s.c ),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _04848_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].singles[2].s.c ),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _04849_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].singles[1].s.c ),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _04850_ (.A(\cb_north.inst.connectaroni.clb1_outputs[3].singles[0].s.c ),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _04851_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[3].s.c ),
    .Y(_00158_));
 sky130_fd_sc_hd__inv_2 _04852_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[2].s.c ),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _04853_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[1].s.c ),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _04854_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[0].s.c ),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _04855_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].singles[3].s.c ),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _04856_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].singles[2].s.c ),
    .Y(_00163_));
 sky130_fd_sc_hd__inv_2 _04857_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].singles[1].s.c ),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _04858_ (.A(\cb_north.inst.connectaroni.clb1_outputs[2].singles[0].s.c ),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_2 _04859_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[3].s.c ),
    .Y(_00166_));
 sky130_fd_sc_hd__inv_2 _04860_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[2].s.c ),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _04861_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[1].s.c ),
    .Y(_00168_));
 sky130_fd_sc_hd__inv_2 _04862_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[0].s.c ),
    .Y(_00169_));
 sky130_fd_sc_hd__inv_2 _04863_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].singles[3].s.c ),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_2 _04864_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].singles[2].s.c ),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _04865_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].singles[1].s.c ),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _04866_ (.A(\cb_north.inst.connectaroni.clb1_outputs[1].singles[0].s.c ),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _04867_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[3].s.c ),
    .Y(_00174_));
 sky130_fd_sc_hd__inv_2 _04868_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[2].s.c ),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _04869_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[1].s.c ),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_2 _04870_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[0].s.c ),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _04871_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].singles[3].s.c ),
    .Y(_00178_));
 sky130_fd_sc_hd__inv_2 _04872_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].singles[2].s.c ),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _04873_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].singles[1].s.c ),
    .Y(_00180_));
 sky130_fd_sc_hd__inv_2 _04874_ (.A(\cb_north.inst.connectaroni.clb1_outputs[0].singles[0].s.c ),
    .Y(_00181_));
 sky130_fd_sc_hd__inv_2 _04875_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[4].s.c ),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _04876_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[3].s.c ),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _04877_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[2].s.c ),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _04878_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[1].s.c ),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _04879_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.c ),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _04880_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[7].s.c ),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _04881_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[6].s.c ),
    .Y(_00188_));
 sky130_fd_sc_hd__inv_2 _04882_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[5].s.c ),
    .Y(_00189_));
 sky130_fd_sc_hd__inv_2 _04883_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[3].s.c ),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _04884_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[2].s.c ),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _04885_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[1].s.c ),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _04886_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.c ),
    .Y(_00213_));
 sky130_fd_sc_hd__inv_2 _04887_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].singles[3].s.c ),
    .Y(_00219_));
 sky130_fd_sc_hd__inv_2 _04888_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].singles[2].s.c ),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _04889_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].singles[1].s.c ),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_2 _04890_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].singles[0].s.c ),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _04891_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].singles[0].s.c ),
    .Y(_00238_));
 sky130_fd_sc_hd__inv_2 _04892_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[4].s.c ),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _04893_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[3].s.c ),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _04894_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[2].s.c ),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _04895_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[1].s.c ),
    .Y(_00242_));
 sky130_fd_sc_hd__inv_2 _04896_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.c ),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _04897_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[7].s.c ),
    .Y(_00244_));
 sky130_fd_sc_hd__inv_2 _04898_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[6].s.c ),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _04899_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[5].s.c ),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _04900_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[4].s.c ),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _04901_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[3].s.c ),
    .Y(_00248_));
 sky130_fd_sc_hd__inv_2 _04902_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[2].s.c ),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _04903_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[1].s.c ),
    .Y(_00250_));
 sky130_fd_sc_hd__inv_2 _04904_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[0].s.c ),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _04905_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].singles[3].s.c ),
    .Y(_00252_));
 sky130_fd_sc_hd__inv_2 _04906_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].singles[2].s.c ),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _04907_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].singles[1].s.c ),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _04908_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].singles[0].s.c ),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_2 _04909_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[4].s.c ),
    .Y(_00256_));
 sky130_fd_sc_hd__inv_2 _04910_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[3].s.c ),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _04911_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[2].s.c ),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _04912_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[1].s.c ),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _04913_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.c ),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _04914_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[7].s.c ),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _04915_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[6].s.c ),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _04916_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[5].s.c ),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _04917_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[4].s.c ),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _04918_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[3].s.c ),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _04919_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[2].s.c ),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _04920_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[1].s.c ),
    .Y(_00267_));
 sky130_fd_sc_hd__inv_2 _04921_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[0].s.c ),
    .Y(_00268_));
 sky130_fd_sc_hd__inv_2 _04922_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].singles[3].s.c ),
    .Y(_00269_));
 sky130_fd_sc_hd__inv_2 _04923_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].singles[2].s.c ),
    .Y(_00270_));
 sky130_fd_sc_hd__inv_2 _04924_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].singles[1].s.c ),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _04925_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].singles[0].s.c ),
    .Y(_00272_));
 sky130_fd_sc_hd__inv_2 _04926_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[4].s.c ),
    .Y(_00273_));
 sky130_fd_sc_hd__inv_2 _04927_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[3].s.c ),
    .Y(_00274_));
 sky130_fd_sc_hd__inv_2 _04928_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[2].s.c ),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _04929_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[1].s.c ),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _04930_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.c ),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_2 _04931_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[7].s.c ),
    .Y(_00278_));
 sky130_fd_sc_hd__inv_2 _04932_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[6].s.c ),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _04933_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[5].s.c ),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _04934_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[4].s.c ),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _04935_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[3].s.c ),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _04936_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[2].s.c ),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _04937_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[1].s.c ),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _04938_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[0].s.c ),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _04939_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].singles[3].s.c ),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _04940_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].singles[2].s.c ),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _04941_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].singles[1].s.c ),
    .Y(_00288_));
 sky130_fd_sc_hd__inv_2 _04942_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].singles[0].s.c ),
    .Y(_00289_));
 sky130_fd_sc_hd__inv_2 _04943_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[4].s.c ),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _04944_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[3].s.c ),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _04945_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[2].s.c ),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _04946_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[1].s.c ),
    .Y(_00293_));
 sky130_fd_sc_hd__inv_2 _04947_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.c ),
    .Y(_00294_));
 sky130_fd_sc_hd__inv_2 _04948_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[7].s.c ),
    .Y(_00295_));
 sky130_fd_sc_hd__inv_2 _04949_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[6].s.c ),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _04950_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[5].s.c ),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _04951_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[4].s.c ),
    .Y(_00298_));
 sky130_fd_sc_hd__inv_2 _04952_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[3].s.c ),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_2 _04953_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[2].s.c ),
    .Y(_00300_));
 sky130_fd_sc_hd__inv_2 _04954_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[1].s.c ),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _04955_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[0].s.c ),
    .Y(_00302_));
 sky130_fd_sc_hd__inv_2 _04956_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].singles[3].s.c ),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _04957_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].singles[2].s.c ),
    .Y(_00304_));
 sky130_fd_sc_hd__inv_2 _04958_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].singles[1].s.c ),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _04959_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].singles[0].s.c ),
    .Y(_00306_));
 sky130_fd_sc_hd__inv_2 _04960_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[4].s.c ),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _04961_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[3].s.c ),
    .Y(_00308_));
 sky130_fd_sc_hd__inv_2 _04962_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[2].s.c ),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _04963_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[1].s.c ),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _04964_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.c ),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _04965_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[7].s.c ),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _04966_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[6].s.c ),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _04967_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[5].s.c ),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _04968_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[4].s.c ),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _04969_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[3].s.c ),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _04970_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[2].s.c ),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _04971_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[1].s.c ),
    .Y(_00318_));
 sky130_fd_sc_hd__inv_2 _04972_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[0].s.c ),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _04973_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].singles[3].s.c ),
    .Y(_00320_));
 sky130_fd_sc_hd__inv_2 _04974_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].singles[2].s.c ),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _04975_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].singles[1].s.c ),
    .Y(_00322_));
 sky130_fd_sc_hd__inv_2 _04976_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].singles[0].s.c ),
    .Y(_00323_));
 sky130_fd_sc_hd__inv_2 _04977_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[4].s.c ),
    .Y(_00324_));
 sky130_fd_sc_hd__inv_2 _04978_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[3].s.c ),
    .Y(_00325_));
 sky130_fd_sc_hd__inv_2 _04979_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[2].s.c ),
    .Y(_00326_));
 sky130_fd_sc_hd__inv_2 _04980_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[1].s.c ),
    .Y(_00327_));
 sky130_fd_sc_hd__inv_2 _04981_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.c ),
    .Y(_00328_));
 sky130_fd_sc_hd__inv_2 _04982_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[7].s.c ),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _04983_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[6].s.c ),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_2 _04984_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[5].s.c ),
    .Y(_00331_));
 sky130_fd_sc_hd__inv_2 _04985_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[4].s.c ),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _04986_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[3].s.c ),
    .Y(_00333_));
 sky130_fd_sc_hd__inv_2 _04987_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[2].s.c ),
    .Y(_00334_));
 sky130_fd_sc_hd__inv_2 _04988_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[1].s.c ),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _04989_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[0].s.c ),
    .Y(_00336_));
 sky130_fd_sc_hd__inv_2 _04990_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].singles[3].s.c ),
    .Y(_00337_));
 sky130_fd_sc_hd__inv_2 _04991_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].singles[2].s.c ),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _04992_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].singles[1].s.c ),
    .Y(_00339_));
 sky130_fd_sc_hd__inv_2 _04993_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].singles[0].s.c ),
    .Y(_00340_));
 sky130_fd_sc_hd__inv_2 _04994_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[4].s.c ),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _04995_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[3].s.c ),
    .Y(_00342_));
 sky130_fd_sc_hd__inv_2 _04996_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[2].s.c ),
    .Y(_00343_));
 sky130_fd_sc_hd__inv_2 _04997_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[1].s.c ),
    .Y(_00344_));
 sky130_fd_sc_hd__inv_2 _04998_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.c ),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _04999_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[7].s.c ),
    .Y(_00346_));
 sky130_fd_sc_hd__inv_2 _05000_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[6].s.c ),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _05001_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[5].s.c ),
    .Y(_00348_));
 sky130_fd_sc_hd__inv_2 _05002_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[4].s.c ),
    .Y(_00349_));
 sky130_fd_sc_hd__inv_2 _05003_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[3].s.c ),
    .Y(_00350_));
 sky130_fd_sc_hd__inv_2 _05004_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[2].s.c ),
    .Y(_00351_));
 sky130_fd_sc_hd__inv_2 _05005_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[1].s.c ),
    .Y(_00352_));
 sky130_fd_sc_hd__inv_2 _05006_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[0].s.c ),
    .Y(_00353_));
 sky130_fd_sc_hd__inv_2 _05007_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].singles[3].s.c ),
    .Y(_00354_));
 sky130_fd_sc_hd__inv_2 _05008_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].singles[2].s.c ),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_2 _05009_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].singles[1].s.c ),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_2 _05010_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].singles[0].s.c ),
    .Y(_00357_));
 sky130_fd_sc_hd__inv_2 _05011_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[4].s.c ),
    .Y(_00358_));
 sky130_fd_sc_hd__inv_2 _05012_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[3].s.c ),
    .Y(_00359_));
 sky130_fd_sc_hd__inv_2 _05013_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[2].s.c ),
    .Y(_00360_));
 sky130_fd_sc_hd__inv_2 _05014_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[1].s.c ),
    .Y(_00361_));
 sky130_fd_sc_hd__inv_2 _05015_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.c ),
    .Y(_00362_));
 sky130_fd_sc_hd__inv_2 _05016_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[7].s.c ),
    .Y(_00363_));
 sky130_fd_sc_hd__inv_2 _05017_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[6].s.c ),
    .Y(_00364_));
 sky130_fd_sc_hd__inv_2 _05018_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[5].s.c ),
    .Y(_00365_));
 sky130_fd_sc_hd__inv_2 _05019_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[4].s.c ),
    .Y(_00366_));
 sky130_fd_sc_hd__inv_2 _05020_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[3].s.c ),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_2 _05021_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[2].s.c ),
    .Y(_00368_));
 sky130_fd_sc_hd__inv_2 _05022_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[1].s.c ),
    .Y(_00369_));
 sky130_fd_sc_hd__inv_2 _05023_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[0].s.c ),
    .Y(_00370_));
 sky130_fd_sc_hd__inv_2 _05024_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].singles[3].s.c ),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _05025_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].singles[2].s.c ),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _05026_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].singles[1].s.c ),
    .Y(_00373_));
 sky130_fd_sc_hd__inv_2 _05027_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].singles[0].s.c ),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_2 _05028_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[4].s.c ),
    .Y(_00375_));
 sky130_fd_sc_hd__inv_2 _05029_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[3].s.c ),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _05030_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[2].s.c ),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _05031_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[1].s.c ),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _05032_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.c ),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _05033_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[7].s.c ),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_2 _05034_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[6].s.c ),
    .Y(_00381_));
 sky130_fd_sc_hd__inv_2 _05035_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[5].s.c ),
    .Y(_00382_));
 sky130_fd_sc_hd__inv_2 _05036_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[4].s.c ),
    .Y(_00383_));
 sky130_fd_sc_hd__inv_2 _05037_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[3].s.c ),
    .Y(_00384_));
 sky130_fd_sc_hd__inv_2 _05038_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[2].s.c ),
    .Y(_00385_));
 sky130_fd_sc_hd__inv_2 _05039_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[1].s.c ),
    .Y(_00386_));
 sky130_fd_sc_hd__inv_2 _05040_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[0].s.c ),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _05041_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].singles[3].s.c ),
    .Y(_00388_));
 sky130_fd_sc_hd__inv_2 _05042_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].singles[2].s.c ),
    .Y(_00389_));
 sky130_fd_sc_hd__inv_2 _05043_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].singles[1].s.c ),
    .Y(_00390_));
 sky130_fd_sc_hd__inv_2 _05044_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[4].s.c ),
    .Y(_00190_));
 sky130_fd_sc_hd__inv_2 _05045_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[3].s.c ),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _05046_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[2].s.c ),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _05047_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[1].s.c ),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_2 _05048_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[0].s.c ),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _05049_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].singles[3].s.c ),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _05050_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].singles[2].s.c ),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _05051_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].singles[1].s.c ),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _05052_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[3].s.c ),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _05053_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[2].s.c ),
    .Y(_00197_));
 sky130_fd_sc_hd__inv_2 _05054_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[1].s.c ),
    .Y(_00203_));
 sky130_fd_sc_hd__inv_2 _05055_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[0].s.c ),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _05056_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].singles[3].s.c ),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _05057_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].singles[2].s.c ),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _05058_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].singles[1].s.c ),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _05059_ (.A(\cb_north.inst.connectaroni.clb0_outputs[4].singles[0].s.c ),
    .Y(_00233_));
 sky130_fd_sc_hd__inv_2 _05060_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[3].s.c ),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _05061_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[2].s.c ),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_2 _05062_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[1].s.c ),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _05063_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.c ),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _05064_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].singles[3].s.c ),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _05065_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].singles[2].s.c ),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _05066_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].singles[1].s.c ),
    .Y(_00228_));
 sky130_fd_sc_hd__inv_2 _05067_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].singles[0].s.c ),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_2 _05068_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[3].s.c ),
    .Y(_00193_));
 sky130_fd_sc_hd__inv_2 _05069_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[2].s.c ),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _05070_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[1].s.c ),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _05071_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.c ),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _05072_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].singles[3].s.c ),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _05073_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].singles[2].s.c ),
    .Y(_00223_));
 sky130_fd_sc_hd__inv_2 _05074_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].singles[1].s.c ),
    .Y(_00229_));
 sky130_fd_sc_hd__inv_2 _05075_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].singles[0].s.c ),
    .Y(_00235_));
 sky130_fd_sc_hd__inv_2 _05076_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[3].s.c ),
    .Y(_00194_));
 sky130_fd_sc_hd__inv_2 _05077_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[2].s.c ),
    .Y(_00200_));
 sky130_fd_sc_hd__inv_2 _05078_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[1].s.c ),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _05079_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.c ),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _05080_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].singles[3].s.c ),
    .Y(_00218_));
 sky130_fd_sc_hd__inv_2 _05081_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].singles[2].s.c ),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _05082_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].singles[1].s.c ),
    .Y(_00230_));
 sky130_fd_sc_hd__inv_2 _05083_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].singles[0].s.c ),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _05084_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].singles[0].s.c ),
    .Y(_00391_));
 sky130_fd_sc_hd__inv_2 _05085_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].directs[4].s.c ),
    .Y(_00392_));
 sky130_fd_sc_hd__inv_2 _05086_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].directs[3].s.c ),
    .Y(_00393_));
 sky130_fd_sc_hd__inv_2 _05087_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].directs[2].s.c ),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _05088_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].directs[1].s.c ),
    .Y(_00395_));
 sky130_fd_sc_hd__inv_2 _05089_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.c ),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _05090_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[7].s.c ),
    .Y(_00397_));
 sky130_fd_sc_hd__inv_2 _05091_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[6].s.c ),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _05092_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[5].s.c ),
    .Y(_00399_));
 sky130_fd_sc_hd__inv_2 _05093_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[4].s.c ),
    .Y(_00400_));
 sky130_fd_sc_hd__inv_2 _05094_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[3].s.c ),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_2 _05095_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[2].s.c ),
    .Y(_00402_));
 sky130_fd_sc_hd__inv_2 _05096_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[1].s.c ),
    .Y(_00403_));
 sky130_fd_sc_hd__inv_2 _05097_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[0].s.c ),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_2 _05098_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].singles[3].s.c ),
    .Y(_00405_));
 sky130_fd_sc_hd__inv_2 _05099_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].singles[2].s.c ),
    .Y(_00406_));
 sky130_fd_sc_hd__inv_2 _05100_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].singles[1].s.c ),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_2 _05101_ (.A(\cb_north.inst.connectaroni.clb0_inputs[9].singles[0].s.c ),
    .Y(_00408_));
 sky130_fd_sc_hd__inv_2 _05102_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].directs[4].s.c ),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _05103_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].directs[3].s.c ),
    .Y(_00410_));
 sky130_fd_sc_hd__inv_2 _05104_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].directs[2].s.c ),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _05105_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].directs[1].s.c ),
    .Y(_00412_));
 sky130_fd_sc_hd__inv_2 _05106_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.c ),
    .Y(_00413_));
 sky130_fd_sc_hd__inv_2 _05107_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[7].s.c ),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _05108_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[6].s.c ),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _05109_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[5].s.c ),
    .Y(_00416_));
 sky130_fd_sc_hd__inv_2 _05110_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[4].s.c ),
    .Y(_00417_));
 sky130_fd_sc_hd__inv_2 _05111_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[3].s.c ),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_2 _05112_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[2].s.c ),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _05113_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[1].s.c ),
    .Y(_00420_));
 sky130_fd_sc_hd__inv_2 _05114_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[0].s.c ),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _05115_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].singles[3].s.c ),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _05116_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].singles[2].s.c ),
    .Y(_00423_));
 sky130_fd_sc_hd__inv_2 _05117_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].singles[1].s.c ),
    .Y(_00424_));
 sky130_fd_sc_hd__inv_2 _05118_ (.A(\cb_north.inst.connectaroni.clb0_inputs[8].singles[0].s.c ),
    .Y(_00425_));
 sky130_fd_sc_hd__inv_2 _05119_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[4].s.c ),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _05120_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[3].s.c ),
    .Y(_00427_));
 sky130_fd_sc_hd__inv_2 _05121_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[2].s.c ),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _05122_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[1].s.c ),
    .Y(_00429_));
 sky130_fd_sc_hd__inv_2 _05123_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.c ),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_2 _05124_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[7].s.c ),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _05125_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[6].s.c ),
    .Y(_00432_));
 sky130_fd_sc_hd__inv_2 _05126_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[5].s.c ),
    .Y(_00433_));
 sky130_fd_sc_hd__inv_2 _05127_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[4].s.c ),
    .Y(_00434_));
 sky130_fd_sc_hd__inv_2 _05128_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[3].s.c ),
    .Y(_00435_));
 sky130_fd_sc_hd__inv_2 _05129_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[2].s.c ),
    .Y(_00436_));
 sky130_fd_sc_hd__inv_2 _05130_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[1].s.c ),
    .Y(_00437_));
 sky130_fd_sc_hd__inv_2 _05131_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[0].s.c ),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _05132_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].singles[3].s.c ),
    .Y(_00439_));
 sky130_fd_sc_hd__inv_2 _05133_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].singles[2].s.c ),
    .Y(_00440_));
 sky130_fd_sc_hd__inv_2 _05134_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].singles[1].s.c ),
    .Y(_00441_));
 sky130_fd_sc_hd__inv_2 _05135_ (.A(\cb_north.inst.connectaroni.clb0_inputs[7].singles[0].s.c ),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _05136_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[4].s.c ),
    .Y(_00443_));
 sky130_fd_sc_hd__inv_2 _05137_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[3].s.c ),
    .Y(_00444_));
 sky130_fd_sc_hd__inv_2 _05138_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[2].s.c ),
    .Y(_00445_));
 sky130_fd_sc_hd__inv_2 _05139_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[1].s.c ),
    .Y(_00446_));
 sky130_fd_sc_hd__inv_2 _05140_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.c ),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _05141_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[7].s.c ),
    .Y(_00448_));
 sky130_fd_sc_hd__inv_2 _05142_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[6].s.c ),
    .Y(_00449_));
 sky130_fd_sc_hd__inv_2 _05143_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[5].s.c ),
    .Y(_00450_));
 sky130_fd_sc_hd__inv_2 _05144_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[4].s.c ),
    .Y(_00451_));
 sky130_fd_sc_hd__inv_2 _05145_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[3].s.c ),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _05146_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[2].s.c ),
    .Y(_00453_));
 sky130_fd_sc_hd__inv_2 _05147_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[1].s.c ),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _05148_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[0].s.c ),
    .Y(_00455_));
 sky130_fd_sc_hd__inv_2 _05149_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].singles[3].s.c ),
    .Y(_00456_));
 sky130_fd_sc_hd__inv_2 _05150_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].singles[2].s.c ),
    .Y(_00457_));
 sky130_fd_sc_hd__inv_2 _05151_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].singles[1].s.c ),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _05152_ (.A(\cb_north.inst.connectaroni.clb0_inputs[6].singles[0].s.c ),
    .Y(_00459_));
 sky130_fd_sc_hd__inv_2 _05153_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].directs[4].s.c ),
    .Y(_00460_));
 sky130_fd_sc_hd__inv_2 _05154_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].directs[3].s.c ),
    .Y(_00461_));
 sky130_fd_sc_hd__inv_2 _05155_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].directs[2].s.c ),
    .Y(_00462_));
 sky130_fd_sc_hd__inv_2 _05156_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].directs[1].s.c ),
    .Y(_00463_));
 sky130_fd_sc_hd__inv_2 _05157_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.c ),
    .Y(_00464_));
 sky130_fd_sc_hd__inv_2 _05158_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[7].s.c ),
    .Y(_00465_));
 sky130_fd_sc_hd__inv_2 _05159_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[6].s.c ),
    .Y(_00466_));
 sky130_fd_sc_hd__inv_2 _05160_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[5].s.c ),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _05161_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[4].s.c ),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _05162_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[3].s.c ),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _05163_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[2].s.c ),
    .Y(_00470_));
 sky130_fd_sc_hd__inv_2 _05164_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[1].s.c ),
    .Y(_00471_));
 sky130_fd_sc_hd__inv_2 _05165_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[0].s.c ),
    .Y(_00472_));
 sky130_fd_sc_hd__inv_2 _05166_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].singles[3].s.c ),
    .Y(_00473_));
 sky130_fd_sc_hd__inv_2 _05167_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].singles[2].s.c ),
    .Y(_00474_));
 sky130_fd_sc_hd__inv_2 _05168_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].singles[1].s.c ),
    .Y(_00475_));
 sky130_fd_sc_hd__inv_2 _05169_ (.A(\cb_north.inst.connectaroni.clb0_inputs[5].singles[0].s.c ),
    .Y(_00476_));
 sky130_fd_sc_hd__inv_2 _05170_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].directs[4].s.c ),
    .Y(_00477_));
 sky130_fd_sc_hd__inv_2 _05171_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].directs[3].s.c ),
    .Y(_00478_));
 sky130_fd_sc_hd__inv_2 _05172_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].directs[2].s.c ),
    .Y(_00479_));
 sky130_fd_sc_hd__inv_2 _05173_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].directs[1].s.c ),
    .Y(_00480_));
 sky130_fd_sc_hd__inv_2 _05174_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.c ),
    .Y(_00481_));
 sky130_fd_sc_hd__inv_2 _05175_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[7].s.c ),
    .Y(_00482_));
 sky130_fd_sc_hd__inv_2 _05176_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[6].s.c ),
    .Y(_00483_));
 sky130_fd_sc_hd__inv_2 _05177_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[5].s.c ),
    .Y(_00484_));
 sky130_fd_sc_hd__inv_2 _05178_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[4].s.c ),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _05179_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[3].s.c ),
    .Y(_00486_));
 sky130_fd_sc_hd__inv_2 _05180_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[2].s.c ),
    .Y(_00487_));
 sky130_fd_sc_hd__inv_2 _05181_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[1].s.c ),
    .Y(_00488_));
 sky130_fd_sc_hd__inv_2 _05182_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[0].s.c ),
    .Y(_00489_));
 sky130_fd_sc_hd__inv_2 _05183_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].singles[3].s.c ),
    .Y(_00490_));
 sky130_fd_sc_hd__inv_2 _05184_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].singles[2].s.c ),
    .Y(_00491_));
 sky130_fd_sc_hd__inv_2 _05185_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].singles[1].s.c ),
    .Y(_00492_));
 sky130_fd_sc_hd__inv_2 _05186_ (.A(\cb_north.inst.connectaroni.clb0_inputs[4].singles[0].s.c ),
    .Y(_00493_));
 sky130_fd_sc_hd__inv_2 _05187_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].directs[4].s.c ),
    .Y(_00494_));
 sky130_fd_sc_hd__inv_2 _05188_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].directs[3].s.c ),
    .Y(_00495_));
 sky130_fd_sc_hd__inv_2 _05189_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].directs[2].s.c ),
    .Y(_00496_));
 sky130_fd_sc_hd__inv_2 _05190_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].directs[1].s.c ),
    .Y(_00497_));
 sky130_fd_sc_hd__inv_2 _05191_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.c ),
    .Y(_00498_));
 sky130_fd_sc_hd__inv_2 _05192_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[7].s.c ),
    .Y(_00499_));
 sky130_fd_sc_hd__inv_2 _05193_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[6].s.c ),
    .Y(_00500_));
 sky130_fd_sc_hd__inv_2 _05194_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[5].s.c ),
    .Y(_00501_));
 sky130_fd_sc_hd__inv_2 _05195_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[4].s.c ),
    .Y(_00502_));
 sky130_fd_sc_hd__inv_2 _05196_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[3].s.c ),
    .Y(_00503_));
 sky130_fd_sc_hd__inv_2 _05197_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[2].s.c ),
    .Y(_00504_));
 sky130_fd_sc_hd__inv_2 _05198_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[1].s.c ),
    .Y(_00505_));
 sky130_fd_sc_hd__inv_2 _05199_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[0].s.c ),
    .Y(_00506_));
 sky130_fd_sc_hd__inv_2 _05200_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].singles[3].s.c ),
    .Y(_00507_));
 sky130_fd_sc_hd__inv_2 _05201_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].singles[2].s.c ),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _05202_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].singles[1].s.c ),
    .Y(_00509_));
 sky130_fd_sc_hd__inv_2 _05203_ (.A(\cb_north.inst.connectaroni.clb0_inputs[3].singles[0].s.c ),
    .Y(_00510_));
 sky130_fd_sc_hd__inv_2 _05204_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[4].s.c ),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _05205_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[3].s.c ),
    .Y(_00512_));
 sky130_fd_sc_hd__inv_2 _05206_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[2].s.c ),
    .Y(_00513_));
 sky130_fd_sc_hd__inv_2 _05207_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[1].s.c ),
    .Y(_00514_));
 sky130_fd_sc_hd__inv_2 _05208_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.c ),
    .Y(_00515_));
 sky130_fd_sc_hd__inv_2 _05209_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[7].s.c ),
    .Y(_00516_));
 sky130_fd_sc_hd__inv_2 _05210_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[6].s.c ),
    .Y(_00517_));
 sky130_fd_sc_hd__inv_2 _05211_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[5].s.c ),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _05212_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[4].s.c ),
    .Y(_00519_));
 sky130_fd_sc_hd__inv_2 _05213_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[3].s.c ),
    .Y(_00520_));
 sky130_fd_sc_hd__inv_2 _05214_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[2].s.c ),
    .Y(_00521_));
 sky130_fd_sc_hd__inv_2 _05215_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[1].s.c ),
    .Y(_00522_));
 sky130_fd_sc_hd__inv_2 _05216_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[0].s.c ),
    .Y(_00523_));
 sky130_fd_sc_hd__inv_2 _05217_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].singles[3].s.c ),
    .Y(_00524_));
 sky130_fd_sc_hd__inv_2 _05218_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].singles[2].s.c ),
    .Y(_00525_));
 sky130_fd_sc_hd__inv_2 _05219_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].singles[1].s.c ),
    .Y(_00526_));
 sky130_fd_sc_hd__inv_2 _05220_ (.A(\cb_north.inst.connectaroni.clb0_inputs[2].singles[0].s.c ),
    .Y(_00527_));
 sky130_fd_sc_hd__inv_2 _05221_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].directs[4].s.c ),
    .Y(_00528_));
 sky130_fd_sc_hd__inv_2 _05222_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].directs[3].s.c ),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_2 _05223_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].directs[2].s.c ),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _05224_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].directs[1].s.c ),
    .Y(_00531_));
 sky130_fd_sc_hd__inv_2 _05225_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.c ),
    .Y(_00532_));
 sky130_fd_sc_hd__inv_2 _05226_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[7].s.c ),
    .Y(_00533_));
 sky130_fd_sc_hd__inv_2 _05227_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[6].s.c ),
    .Y(_00534_));
 sky130_fd_sc_hd__inv_2 _05228_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[5].s.c ),
    .Y(_00535_));
 sky130_fd_sc_hd__inv_2 _05229_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[4].s.c ),
    .Y(_00536_));
 sky130_fd_sc_hd__inv_2 _05230_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[3].s.c ),
    .Y(_00537_));
 sky130_fd_sc_hd__inv_2 _05231_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[2].s.c ),
    .Y(_00538_));
 sky130_fd_sc_hd__inv_2 _05232_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[1].s.c ),
    .Y(_00539_));
 sky130_fd_sc_hd__inv_2 _05233_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[0].s.c ),
    .Y(_00540_));
 sky130_fd_sc_hd__inv_2 _05234_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].singles[3].s.c ),
    .Y(_00541_));
 sky130_fd_sc_hd__inv_2 _05235_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].singles[2].s.c ),
    .Y(_00542_));
 sky130_fd_sc_hd__inv_2 _05236_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].singles[1].s.c ),
    .Y(_00543_));
 sky130_fd_sc_hd__inv_2 _05237_ (.A(\cb_north.inst.connectaroni.clb0_inputs[1].singles[0].s.c ),
    .Y(_00544_));
 sky130_fd_sc_hd__inv_2 _05238_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].directs[4].s.c ),
    .Y(_00545_));
 sky130_fd_sc_hd__inv_2 _05239_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].directs[3].s.c ),
    .Y(_00546_));
 sky130_fd_sc_hd__inv_2 _05240_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].directs[2].s.c ),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _05241_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].directs[1].s.c ),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _05242_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.c ),
    .Y(_00549_));
 sky130_fd_sc_hd__inv_2 _05243_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[7].s.c ),
    .Y(_00550_));
 sky130_fd_sc_hd__inv_2 _05244_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[6].s.c ),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_2 _05245_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[5].s.c ),
    .Y(_00552_));
 sky130_fd_sc_hd__inv_2 _05246_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[4].s.c ),
    .Y(_00553_));
 sky130_fd_sc_hd__inv_2 _05247_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[3].s.c ),
    .Y(_00554_));
 sky130_fd_sc_hd__inv_2 _05248_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[2].s.c ),
    .Y(_00555_));
 sky130_fd_sc_hd__inv_2 _05249_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[1].s.c ),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _05250_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[0].s.c ),
    .Y(_00557_));
 sky130_fd_sc_hd__inv_2 _05251_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].singles[3].s.c ),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_2 _05252_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].singles[2].s.c ),
    .Y(_00559_));
 sky130_fd_sc_hd__inv_2 _05253_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].singles[1].s.c ),
    .Y(_00560_));
 sky130_fd_sc_hd__inv_2 _05254_ (.A(\cb_north.inst.connectaroni.clb0_inputs[0].singles[0].s.c ),
    .Y(_00561_));
 sky130_fd_sc_hd__inv_2 _05255_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[3].s.c ),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _05256_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[2].s.c ),
    .Y(_00563_));
 sky130_fd_sc_hd__inv_2 _05257_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[1].s.c ),
    .Y(_00564_));
 sky130_fd_sc_hd__inv_2 _05258_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[0].s.c ),
    .Y(_00565_));
 sky130_fd_sc_hd__inv_2 _05259_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].singles[3].s.c ),
    .Y(_00566_));
 sky130_fd_sc_hd__inv_2 _05260_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].singles[2].s.c ),
    .Y(_00567_));
 sky130_fd_sc_hd__inv_2 _05261_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].singles[1].s.c ),
    .Y(_00568_));
 sky130_fd_sc_hd__inv_2 _05262_ (.A(\cb_east.inst.connectaroni.clb1_outputs[4].singles[0].s.c ),
    .Y(_00569_));
 sky130_fd_sc_hd__inv_2 _05263_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[3].s.c ),
    .Y(_00570_));
 sky130_fd_sc_hd__inv_2 _05264_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[2].s.c ),
    .Y(_00571_));
 sky130_fd_sc_hd__inv_2 _05265_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[1].s.c ),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _05266_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[0].s.c ),
    .Y(_00573_));
 sky130_fd_sc_hd__inv_2 _05267_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].singles[3].s.c ),
    .Y(_00574_));
 sky130_fd_sc_hd__inv_2 _05268_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].singles[2].s.c ),
    .Y(_00575_));
 sky130_fd_sc_hd__inv_2 _05269_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].singles[1].s.c ),
    .Y(_00576_));
 sky130_fd_sc_hd__inv_2 _05270_ (.A(\cb_east.inst.connectaroni.clb1_outputs[3].singles[0].s.c ),
    .Y(_00577_));
 sky130_fd_sc_hd__inv_2 _05271_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[3].s.c ),
    .Y(_00578_));
 sky130_fd_sc_hd__inv_2 _05272_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[2].s.c ),
    .Y(_00579_));
 sky130_fd_sc_hd__inv_2 _05273_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[1].s.c ),
    .Y(_00580_));
 sky130_fd_sc_hd__inv_2 _05274_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[0].s.c ),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _05275_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].singles[3].s.c ),
    .Y(_00582_));
 sky130_fd_sc_hd__inv_2 _05276_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].singles[2].s.c ),
    .Y(_00583_));
 sky130_fd_sc_hd__inv_2 _05277_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].singles[1].s.c ),
    .Y(_00584_));
 sky130_fd_sc_hd__inv_2 _05278_ (.A(\cb_east.inst.connectaroni.clb1_outputs[2].singles[0].s.c ),
    .Y(_00585_));
 sky130_fd_sc_hd__inv_2 _05279_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[3].s.c ),
    .Y(_00586_));
 sky130_fd_sc_hd__inv_2 _05280_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[2].s.c ),
    .Y(_00587_));
 sky130_fd_sc_hd__inv_2 _05281_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[1].s.c ),
    .Y(_00588_));
 sky130_fd_sc_hd__inv_2 _05282_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[0].s.c ),
    .Y(_00589_));
 sky130_fd_sc_hd__inv_2 _05283_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].singles[3].s.c ),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_2 _05284_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].singles[2].s.c ),
    .Y(_00591_));
 sky130_fd_sc_hd__inv_2 _05285_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].singles[1].s.c ),
    .Y(_00592_));
 sky130_fd_sc_hd__inv_2 _05286_ (.A(\cb_east.inst.connectaroni.clb1_outputs[1].singles[0].s.c ),
    .Y(_00593_));
 sky130_fd_sc_hd__inv_2 _05287_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[3].s.c ),
    .Y(_00594_));
 sky130_fd_sc_hd__inv_2 _05288_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[2].s.c ),
    .Y(_00595_));
 sky130_fd_sc_hd__inv_2 _05289_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[1].s.c ),
    .Y(_00596_));
 sky130_fd_sc_hd__inv_2 _05290_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[0].s.c ),
    .Y(_00597_));
 sky130_fd_sc_hd__inv_2 _05291_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].singles[3].s.c ),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _05292_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].singles[2].s.c ),
    .Y(_00599_));
 sky130_fd_sc_hd__inv_2 _05293_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].singles[1].s.c ),
    .Y(_00600_));
 sky130_fd_sc_hd__inv_2 _05294_ (.A(\cb_east.inst.connectaroni.clb1_outputs[0].singles[0].s.c ),
    .Y(_00601_));
 sky130_fd_sc_hd__inv_2 _05295_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[4].s.c ),
    .Y(_00602_));
 sky130_fd_sc_hd__inv_2 _05296_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[3].s.c ),
    .Y(_00603_));
 sky130_fd_sc_hd__inv_2 _05297_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[2].s.c ),
    .Y(_00604_));
 sky130_fd_sc_hd__inv_2 _05298_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[1].s.c ),
    .Y(_00605_));
 sky130_fd_sc_hd__inv_2 _05299_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.c ),
    .Y(_00606_));
 sky130_fd_sc_hd__inv_2 _05300_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[7].s.c ),
    .Y(_00607_));
 sky130_fd_sc_hd__inv_2 _05301_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[6].s.c ),
    .Y(_00608_));
 sky130_fd_sc_hd__inv_2 _05302_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[5].s.c ),
    .Y(_00609_));
 sky130_fd_sc_hd__inv_2 _05303_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[3].s.c ),
    .Y(_00615_));
 sky130_fd_sc_hd__inv_2 _05304_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[2].s.c ),
    .Y(_00621_));
 sky130_fd_sc_hd__inv_2 _05305_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[1].s.c ),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _05306_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.c ),
    .Y(_00633_));
 sky130_fd_sc_hd__inv_2 _05307_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].singles[3].s.c ),
    .Y(_00639_));
 sky130_fd_sc_hd__inv_2 _05308_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].singles[2].s.c ),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _05309_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].singles[1].s.c ),
    .Y(_00651_));
 sky130_fd_sc_hd__inv_2 _05310_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].singles[0].s.c ),
    .Y(_00657_));
 sky130_fd_sc_hd__inv_2 _05311_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].singles[0].s.c ),
    .Y(_00658_));
 sky130_fd_sc_hd__inv_2 _05312_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[4].s.c ),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_2 _05313_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[3].s.c ),
    .Y(_00660_));
 sky130_fd_sc_hd__inv_2 _05314_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[2].s.c ),
    .Y(_00661_));
 sky130_fd_sc_hd__inv_2 _05315_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[1].s.c ),
    .Y(_00662_));
 sky130_fd_sc_hd__inv_2 _05316_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.c ),
    .Y(_00663_));
 sky130_fd_sc_hd__inv_2 _05317_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[7].s.c ),
    .Y(_00664_));
 sky130_fd_sc_hd__inv_2 _05318_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[6].s.c ),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_2 _05319_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[5].s.c ),
    .Y(_00666_));
 sky130_fd_sc_hd__inv_2 _05320_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[4].s.c ),
    .Y(_00667_));
 sky130_fd_sc_hd__inv_2 _05321_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[3].s.c ),
    .Y(_00668_));
 sky130_fd_sc_hd__inv_2 _05322_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[2].s.c ),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_2 _05323_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[1].s.c ),
    .Y(_00670_));
 sky130_fd_sc_hd__inv_2 _05324_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[0].s.c ),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _05325_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].singles[3].s.c ),
    .Y(_00672_));
 sky130_fd_sc_hd__inv_2 _05326_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].singles[2].s.c ),
    .Y(_00673_));
 sky130_fd_sc_hd__inv_2 _05327_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].singles[1].s.c ),
    .Y(_00674_));
 sky130_fd_sc_hd__inv_2 _05328_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].singles[0].s.c ),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _05329_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[4].s.c ),
    .Y(_00676_));
 sky130_fd_sc_hd__inv_2 _05330_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[3].s.c ),
    .Y(_00677_));
 sky130_fd_sc_hd__inv_2 _05331_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[2].s.c ),
    .Y(_00678_));
 sky130_fd_sc_hd__inv_2 _05332_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[1].s.c ),
    .Y(_00679_));
 sky130_fd_sc_hd__inv_2 _05333_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.c ),
    .Y(_00680_));
 sky130_fd_sc_hd__inv_2 _05334_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[7].s.c ),
    .Y(_00681_));
 sky130_fd_sc_hd__inv_2 _05335_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[6].s.c ),
    .Y(_00682_));
 sky130_fd_sc_hd__inv_2 _05336_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[5].s.c ),
    .Y(_00683_));
 sky130_fd_sc_hd__inv_2 _05337_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[4].s.c ),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _05338_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[3].s.c ),
    .Y(_00685_));
 sky130_fd_sc_hd__mux2_1 _05339_ (.A0(_04315_),
    .A1(\slice.configuroni.comb_config[131] ),
    .S(set_out_hard),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _05340_ (.A0(\slice.sliceluroni.muxes.config_state[0] ),
    .A1(\slice.configuroni.comb_config[132] ),
    .S(set_out_hard),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _05341_ (.A0(\slice.sliceluroni.muxes.config_state[1] ),
    .A1(\slice.configuroni.comb_config[133] ),
    .S(set_out_hard),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _05342_ (.A0(\slice.sliceluroni.use_cc ),
    .A1(\slice.configuroni.comb_config[134] ),
    .S(set_out_hard),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _05343_ (.A0(_04168_),
    .A1(\slice.configuroni.comb_config[32] ),
    .S(set_out_hard),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _05344_ (.A0(_04217_),
    .A1(\slice.configuroni.comb_config[65] ),
    .S(set_out_hard),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _05345_ (.A0(_04266_),
    .A1(\slice.configuroni.comb_config[98] ),
    .S(set_out_hard),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _05346_ (.A0(clb_west_out[2]),
    .A1(_00053_),
    .S(_00000_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _05347_ (.A0(clb_west_out[3]),
    .A1(_00054_),
    .S(_00000_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _05348_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .A1(_00055_),
    .S(_00000_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _05349_ (.A0(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .A1(_00056_),
    .S(_00000_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _05350_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .A1(_00049_),
    .S(_00000_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _05351_ (.A0(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .A1(_00050_),
    .S(_00000_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _05352_ (.A0(clb_south_out[2]),
    .A1(_00051_),
    .S(_00000_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _05353_ (.A0(clb_south_out[3]),
    .A1(_00052_),
    .S(_00000_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _05354_ (.A0(\cb_east.inst.configuroni.comb_shifter.config_data[421] ),
    .A1(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .S(psn_net_14),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _05355_ (.A0(shift_out_hard),
    .A1(\cb_east.inst.cb_conf_bus[1] ),
    .S(psn_net_14),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _05356_ (.A0(\cb_east.inst.cb_conf_bus[1] ),
    .A1(\cb_east.inst.cb_conf_bus[2] ),
    .S(psn_net_18),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _05357_ (.A0(\cb_east.inst.cb_conf_bus[2] ),
    .A1(\cb_east.inst.cb_conf_bus[3] ),
    .S(psn_net_18),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _05358_ (.A0(\cb_east.inst.cb_conf_bus[3] ),
    .A1(\cb_east.inst.cb_conf_bus[4] ),
    .S(psn_net_18),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _05359_ (.A0(\cb_east.inst.cb_conf_bus[4] ),
    .A1(\cb_east.inst.cb_conf_bus[5] ),
    .S(psn_net_18),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _05360_ (.A0(\cb_east.inst.cb_conf_bus[5] ),
    .A1(\cb_east.inst.cb_conf_bus[6] ),
    .S(psn_net_18),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _05361_ (.A0(\cb_east.inst.cb_conf_bus[6] ),
    .A1(\cb_east.inst.cb_conf_bus[7] ),
    .S(psn_net_18),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _05362_ (.A0(\cb_east.inst.cb_conf_bus[7] ),
    .A1(\cb_east.inst.cb_conf_bus[8] ),
    .S(psn_net_18),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _05363_ (.A0(\cb_east.inst.cb_conf_bus[8] ),
    .A1(\cb_east.inst.cb_conf_bus[9] ),
    .S(psn_net_21),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _05364_ (.A0(\cb_east.inst.cb_conf_bus[9] ),
    .A1(\cb_east.inst.cb_conf_bus[10] ),
    .S(psn_net_21),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _05365_ (.A0(\cb_east.inst.cb_conf_bus[10] ),
    .A1(\cb_east.inst.cb_conf_bus[11] ),
    .S(psn_net_21),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _05366_ (.A0(\cb_east.inst.cb_conf_bus[11] ),
    .A1(\cb_east.inst.cb_conf_bus[12] ),
    .S(psn_net_21),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _05367_ (.A0(\cb_east.inst.cb_conf_bus[12] ),
    .A1(\cb_east.inst.cb_conf_bus[13] ),
    .S(psn_net_21),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _05368_ (.A0(\cb_east.inst.cb_conf_bus[13] ),
    .A1(\cb_east.inst.cb_conf_bus[14] ),
    .S(psn_net_21),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _05369_ (.A0(\cb_east.inst.cb_conf_bus[14] ),
    .A1(\cb_east.inst.cb_conf_bus[15] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _05370_ (.A0(\cb_east.inst.cb_conf_bus[15] ),
    .A1(\cb_east.inst.cb_conf_bus[16] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _05371_ (.A0(\cb_east.inst.cb_conf_bus[16] ),
    .A1(\cb_east.inst.cb_conf_bus[17] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _05372_ (.A0(\cb_east.inst.cb_conf_bus[17] ),
    .A1(\cb_east.inst.cb_conf_bus[18] ),
    .S(psn_net_20),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _05373_ (.A0(\cb_east.inst.cb_conf_bus[18] ),
    .A1(\cb_east.inst.cb_conf_bus[19] ),
    .S(psn_net_20),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _05374_ (.A0(\cb_east.inst.cb_conf_bus[19] ),
    .A1(\cb_east.inst.cb_conf_bus[20] ),
    .S(psn_net_20),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_1 _05375_ (.A0(\cb_east.inst.cb_conf_bus[20] ),
    .A1(\cb_east.inst.cb_conf_bus[21] ),
    .S(psn_net_20),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_1 _05376_ (.A0(\cb_east.inst.cb_conf_bus[21] ),
    .A1(\cb_east.inst.cb_conf_bus[22] ),
    .S(psn_net_20),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _05377_ (.A0(\cb_east.inst.cb_conf_bus[22] ),
    .A1(\cb_east.inst.cb_conf_bus[23] ),
    .S(psn_net_20),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _05378_ (.A0(\cb_east.inst.cb_conf_bus[23] ),
    .A1(\cb_east.inst.cb_conf_bus[24] ),
    .S(psn_net_20),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_1 _05379_ (.A0(\cb_east.inst.cb_conf_bus[24] ),
    .A1(\cb_east.inst.cb_conf_bus[25] ),
    .S(psn_net_20),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _05380_ (.A0(\cb_east.inst.cb_conf_bus[25] ),
    .A1(\cb_east.inst.cb_conf_bus[26] ),
    .S(psn_net_20),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _05381_ (.A0(\cb_east.inst.cb_conf_bus[26] ),
    .A1(\cb_east.inst.cb_conf_bus[27] ),
    .S(psn_net_20),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _05382_ (.A0(\cb_east.inst.cb_conf_bus[27] ),
    .A1(\cb_east.inst.cb_conf_bus[28] ),
    .S(psn_net_20),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _05383_ (.A0(\cb_east.inst.cb_conf_bus[28] ),
    .A1(\cb_east.inst.cb_conf_bus[29] ),
    .S(psn_net_20),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _05384_ (.A0(\cb_east.inst.cb_conf_bus[29] ),
    .A1(\cb_east.inst.cb_conf_bus[30] ),
    .S(psn_net_20),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _05385_ (.A0(\cb_east.inst.cb_conf_bus[30] ),
    .A1(\cb_east.inst.cb_conf_bus[31] ),
    .S(psn_net_20),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _05386_ (.A0(\cb_east.inst.cb_conf_bus[31] ),
    .A1(\cb_east.inst.cb_conf_bus[32] ),
    .S(psn_net_20),
    .X(_02102_));
 sky130_fd_sc_hd__mux2_1 _05387_ (.A0(\cb_east.inst.cb_conf_bus[32] ),
    .A1(\cb_east.inst.cb_conf_bus[33] ),
    .S(psn_net_20),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _05388_ (.A0(\cb_east.inst.cb_conf_bus[33] ),
    .A1(\cb_east.inst.cb_conf_bus[34] ),
    .S(psn_net_20),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _05389_ (.A0(\cb_east.inst.cb_conf_bus[34] ),
    .A1(\cb_east.inst.cb_conf_bus[35] ),
    .S(psn_net_20),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _05390_ (.A0(\cb_east.inst.cb_conf_bus[35] ),
    .A1(\cb_east.inst.cb_conf_bus[36] ),
    .S(psn_net_20),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _05391_ (.A0(\cb_east.inst.cb_conf_bus[36] ),
    .A1(\cb_east.inst.cb_conf_bus[37] ),
    .S(psn_net_20),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _05392_ (.A0(\cb_east.inst.cb_conf_bus[37] ),
    .A1(\cb_east.inst.cb_conf_bus[38] ),
    .S(psn_net_20),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _05393_ (.A0(\cb_east.inst.cb_conf_bus[38] ),
    .A1(\cb_east.inst.cb_conf_bus[39] ),
    .S(psn_net_20),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _05394_ (.A0(\cb_east.inst.cb_conf_bus[39] ),
    .A1(\cb_east.inst.cb_conf_bus[40] ),
    .S(psn_net_20),
    .X(_02118_));
 sky130_fd_sc_hd__mux2_1 _05395_ (.A0(\cb_east.inst.cb_conf_bus[40] ),
    .A1(\cb_east.inst.cb_conf_bus[41] ),
    .S(psn_net_20),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _05396_ (.A0(\cb_east.inst.cb_conf_bus[41] ),
    .A1(\cb_east.inst.cb_conf_bus[42] ),
    .S(psn_net_20),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _05397_ (.A0(\cb_east.inst.cb_conf_bus[42] ),
    .A1(\cb_east.inst.cb_conf_bus[43] ),
    .S(psn_net_20),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _05398_ (.A0(\cb_east.inst.cb_conf_bus[43] ),
    .A1(\cb_east.inst.cb_conf_bus[44] ),
    .S(psn_net_20),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _05399_ (.A0(\cb_east.inst.cb_conf_bus[44] ),
    .A1(\cb_east.inst.cb_conf_bus[45] ),
    .S(psn_net_2),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _05400_ (.A0(\cb_east.inst.cb_conf_bus[45] ),
    .A1(\cb_east.inst.cb_conf_bus[46] ),
    .S(psn_net_2),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _05401_ (.A0(\cb_east.inst.cb_conf_bus[46] ),
    .A1(\cb_east.inst.cb_conf_bus[47] ),
    .S(psn_net_2),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _05402_ (.A0(\cb_east.inst.cb_conf_bus[47] ),
    .A1(\cb_east.inst.cb_conf_bus[48] ),
    .S(psn_net_2),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _05403_ (.A0(\cb_east.inst.cb_conf_bus[48] ),
    .A1(\cb_east.inst.cb_conf_bus[49] ),
    .S(psn_net_2),
    .X(_02136_));
 sky130_fd_sc_hd__mux2_1 _05404_ (.A0(\cb_east.inst.cb_conf_bus[49] ),
    .A1(\cb_east.inst.cb_conf_bus[50] ),
    .S(psn_net_2),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _05405_ (.A0(\cb_east.inst.cb_conf_bus[50] ),
    .A1(\cb_east.inst.cb_conf_bus[51] ),
    .S(psn_net_2),
    .X(_02140_));
 sky130_fd_sc_hd__mux2_1 _05406_ (.A0(\cb_east.inst.cb_conf_bus[51] ),
    .A1(\cb_east.inst.cb_conf_bus[52] ),
    .S(psn_net_2),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _05407_ (.A0(\cb_east.inst.cb_conf_bus[52] ),
    .A1(\cb_east.inst.cb_conf_bus[53] ),
    .S(psn_net_2),
    .X(_02144_));
 sky130_fd_sc_hd__mux2_1 _05408_ (.A0(\cb_east.inst.cb_conf_bus[53] ),
    .A1(\cb_east.inst.cb_conf_bus[54] ),
    .S(psn_net_2),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _05409_ (.A0(\cb_east.inst.cb_conf_bus[54] ),
    .A1(\cb_east.inst.cb_conf_bus[55] ),
    .S(psn_net_2),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _05410_ (.A0(\cb_east.inst.cb_conf_bus[55] ),
    .A1(\cb_east.inst.cb_conf_bus[56] ),
    .S(psn_net_23),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _05411_ (.A0(\cb_east.inst.cb_conf_bus[56] ),
    .A1(\cb_east.inst.cb_conf_bus[57] ),
    .S(psn_net_23),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _05412_ (.A0(\cb_east.inst.cb_conf_bus[57] ),
    .A1(\cb_east.inst.cb_conf_bus[58] ),
    .S(psn_net_23),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _05413_ (.A0(\cb_east.inst.cb_conf_bus[58] ),
    .A1(\cb_east.inst.cb_conf_bus[59] ),
    .S(psn_net_0),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _05414_ (.A0(\cb_east.inst.cb_conf_bus[59] ),
    .A1(\cb_east.inst.cb_conf_bus[60] ),
    .S(psn_net_0),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _05415_ (.A0(\cb_east.inst.cb_conf_bus[60] ),
    .A1(\cb_east.inst.cb_conf_bus[61] ),
    .S(psn_net_0),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _05416_ (.A0(\cb_east.inst.cb_conf_bus[61] ),
    .A1(\cb_east.inst.cb_conf_bus[62] ),
    .S(psn_net_0),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _05417_ (.A0(\cb_east.inst.cb_conf_bus[62] ),
    .A1(\cb_east.inst.cb_conf_bus[63] ),
    .S(psn_net_23),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _05418_ (.A0(\cb_east.inst.cb_conf_bus[63] ),
    .A1(\cb_east.inst.cb_conf_bus[64] ),
    .S(psn_net_23),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _05419_ (.A0(\cb_east.inst.cb_conf_bus[64] ),
    .A1(\cb_east.inst.cb_conf_bus[65] ),
    .S(psn_net_23),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _05420_ (.A0(\cb_east.inst.cb_conf_bus[65] ),
    .A1(\cb_east.inst.cb_conf_bus[66] ),
    .S(psn_net_23),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _05421_ (.A0(\cb_east.inst.cb_conf_bus[66] ),
    .A1(\cb_east.inst.cb_conf_bus[67] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _05422_ (.A0(\cb_east.inst.cb_conf_bus[67] ),
    .A1(\cb_east.inst.cb_conf_bus[68] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_1 _05423_ (.A0(\cb_east.inst.cb_conf_bus[68] ),
    .A1(\cb_east.inst.cb_conf_bus[69] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _05424_ (.A0(\cb_east.inst.cb_conf_bus[69] ),
    .A1(\cb_east.inst.cb_conf_bus[70] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _05425_ (.A0(\cb_east.inst.cb_conf_bus[70] ),
    .A1(\cb_east.inst.cb_conf_bus[71] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _05426_ (.A0(\cb_east.inst.cb_conf_bus[71] ),
    .A1(\cb_east.inst.cb_conf_bus[72] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _05427_ (.A0(\cb_east.inst.cb_conf_bus[72] ),
    .A1(\cb_east.inst.cb_conf_bus[73] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _05428_ (.A0(\cb_east.inst.cb_conf_bus[73] ),
    .A1(\cb_east.inst.cb_conf_bus[74] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _05429_ (.A0(\cb_east.inst.cb_conf_bus[74] ),
    .A1(\cb_east.inst.cb_conf_bus[75] ),
    .S(psn_net_21),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _05430_ (.A0(\cb_east.inst.cb_conf_bus[75] ),
    .A1(\cb_east.inst.cb_conf_bus[76] ),
    .S(psn_net_21),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _05431_ (.A0(\cb_east.inst.cb_conf_bus[76] ),
    .A1(\cb_east.inst.cb_conf_bus[77] ),
    .S(psn_net_21),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _05432_ (.A0(\cb_east.inst.cb_conf_bus[77] ),
    .A1(\cb_east.inst.cb_conf_bus[78] ),
    .S(psn_net_21),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _05433_ (.A0(\cb_east.inst.cb_conf_bus[78] ),
    .A1(\cb_east.inst.cb_conf_bus[79] ),
    .S(psn_net_21),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _05434_ (.A0(\cb_east.inst.cb_conf_bus[79] ),
    .A1(\cb_east.inst.cb_conf_bus[80] ),
    .S(psn_net_21),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _05435_ (.A0(\cb_east.inst.cb_conf_bus[80] ),
    .A1(\cb_east.inst.cb_conf_bus[81] ),
    .S(psn_net_21),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _05436_ (.A0(\cb_east.inst.cb_conf_bus[81] ),
    .A1(\cb_east.inst.cb_conf_bus[82] ),
    .S(psn_net_21),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _05437_ (.A0(\cb_east.inst.cb_conf_bus[82] ),
    .A1(\cb_east.inst.cb_conf_bus[83] ),
    .S(psn_net_21),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _05438_ (.A0(\cb_east.inst.cb_conf_bus[83] ),
    .A1(\cb_east.inst.cb_conf_bus[84] ),
    .S(psn_net_21),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _05439_ (.A0(\cb_east.inst.cb_conf_bus[84] ),
    .A1(\cb_east.inst.cb_conf_bus[85] ),
    .S(psn_net_21),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _05440_ (.A0(\cb_east.inst.cb_conf_bus[85] ),
    .A1(\cb_east.inst.cb_conf_bus[86] ),
    .S(psn_net_21),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _05441_ (.A0(\cb_east.inst.cb_conf_bus[86] ),
    .A1(\cb_east.inst.cb_conf_bus[87] ),
    .S(psn_net_21),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _05442_ (.A0(\cb_east.inst.cb_conf_bus[87] ),
    .A1(\cb_east.inst.cb_conf_bus[88] ),
    .S(psn_net_21),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _05443_ (.A0(\cb_east.inst.cb_conf_bus[88] ),
    .A1(\cb_east.inst.cb_conf_bus[89] ),
    .S(psn_net_14),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _05444_ (.A0(\cb_east.inst.cb_conf_bus[89] ),
    .A1(\cb_east.inst.cb_conf_bus[90] ),
    .S(psn_net_14),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _05445_ (.A0(\cb_east.inst.cb_conf_bus[90] ),
    .A1(\cb_east.inst.cb_conf_bus[91] ),
    .S(psn_net_14),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _05446_ (.A0(\cb_east.inst.cb_conf_bus[91] ),
    .A1(\cb_east.inst.cb_conf_bus[92] ),
    .S(psn_net_14),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _05447_ (.A0(\cb_east.inst.cb_conf_bus[92] ),
    .A1(\cb_east.inst.cb_conf_bus[93] ),
    .S(psn_net_14),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _05448_ (.A0(\cb_east.inst.cb_conf_bus[93] ),
    .A1(\cb_east.inst.cb_conf_bus[94] ),
    .S(psn_net_21),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _05449_ (.A0(\cb_east.inst.cb_conf_bus[94] ),
    .A1(\cb_east.inst.cb_conf_bus[95] ),
    .S(psn_net_21),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _05450_ (.A0(\cb_east.inst.cb_conf_bus[95] ),
    .A1(\cb_east.inst.cb_conf_bus[96] ),
    .S(psn_net_21),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _05451_ (.A0(\cb_east.inst.cb_conf_bus[96] ),
    .A1(\cb_east.inst.cb_conf_bus[97] ),
    .S(psn_net_21),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _05452_ (.A0(\cb_east.inst.cb_conf_bus[97] ),
    .A1(\cb_east.inst.cb_conf_bus[98] ),
    .S(psn_net_21),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _05453_ (.A0(\cb_east.inst.cb_conf_bus[98] ),
    .A1(\cb_east.inst.cb_conf_bus[99] ),
    .S(psn_net_21),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _05454_ (.A0(\cb_east.inst.cb_conf_bus[99] ),
    .A1(\cb_east.inst.cb_conf_bus[100] ),
    .S(psn_net_21),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _05455_ (.A0(\cb_east.inst.cb_conf_bus[100] ),
    .A1(\cb_east.inst.cb_conf_bus[101] ),
    .S(psn_net_21),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _05456_ (.A0(\cb_east.inst.cb_conf_bus[101] ),
    .A1(\cb_east.inst.cb_conf_bus[102] ),
    .S(psn_net_21),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _05457_ (.A0(\cb_east.inst.cb_conf_bus[102] ),
    .A1(\cb_east.inst.cb_conf_bus[103] ),
    .S(psn_net_21),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _05458_ (.A0(\cb_east.inst.cb_conf_bus[103] ),
    .A1(\cb_east.inst.cb_conf_bus[104] ),
    .S(psn_net_21),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _05459_ (.A0(\cb_east.inst.cb_conf_bus[104] ),
    .A1(\cb_east.inst.cb_conf_bus[105] ),
    .S(psn_net_21),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _05460_ (.A0(\cb_east.inst.cb_conf_bus[105] ),
    .A1(\cb_east.inst.cb_conf_bus[106] ),
    .S(psn_net_21),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _05461_ (.A0(\cb_east.inst.cb_conf_bus[106] ),
    .A1(\cb_east.inst.cb_conf_bus[107] ),
    .S(psn_net_21),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _05462_ (.A0(\cb_east.inst.cb_conf_bus[107] ),
    .A1(\cb_east.inst.cb_conf_bus[108] ),
    .S(psn_net_21),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _05463_ (.A0(\cb_east.inst.cb_conf_bus[108] ),
    .A1(\cb_east.inst.cb_conf_bus[109] ),
    .S(psn_net_21),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _05464_ (.A0(\cb_east.inst.cb_conf_bus[109] ),
    .A1(\cb_east.inst.cb_conf_bus[110] ),
    .S(psn_net_21),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _05465_ (.A0(\cb_east.inst.cb_conf_bus[110] ),
    .A1(\cb_east.inst.cb_conf_bus[111] ),
    .S(psn_net_21),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _05466_ (.A0(\cb_east.inst.cb_conf_bus[111] ),
    .A1(\cb_east.inst.cb_conf_bus[112] ),
    .S(psn_net_21),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _05467_ (.A0(\cb_east.inst.cb_conf_bus[112] ),
    .A1(\cb_east.inst.cb_conf_bus[113] ),
    .S(psn_net_21),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _05468_ (.A0(\cb_east.inst.cb_conf_bus[113] ),
    .A1(\cb_east.inst.cb_conf_bus[114] ),
    .S(psn_net_21),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _05469_ (.A0(\cb_east.inst.cb_conf_bus[114] ),
    .A1(\cb_east.inst.cb_conf_bus[115] ),
    .S(psn_net_21),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _05470_ (.A0(\cb_east.inst.cb_conf_bus[115] ),
    .A1(\cb_east.inst.cb_conf_bus[116] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _05471_ (.A0(\cb_east.inst.cb_conf_bus[116] ),
    .A1(\cb_east.inst.cb_conf_bus[117] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _05472_ (.A0(\cb_east.inst.cb_conf_bus[117] ),
    .A1(\cb_east.inst.cb_conf_bus[118] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _05473_ (.A0(\cb_east.inst.cb_conf_bus[118] ),
    .A1(\cb_east.inst.cb_conf_bus[119] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _05474_ (.A0(\cb_east.inst.cb_conf_bus[119] ),
    .A1(\cb_east.inst.cb_conf_bus[120] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _05475_ (.A0(\cb_east.inst.cb_conf_bus[120] ),
    .A1(\cb_east.inst.cb_conf_bus[121] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _05476_ (.A0(\cb_east.inst.cb_conf_bus[121] ),
    .A1(\cb_east.inst.cb_conf_bus[122] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _05477_ (.A0(\cb_east.inst.cb_conf_bus[122] ),
    .A1(\cb_east.inst.cb_conf_bus[123] ),
    .S(psn_net_0),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _05478_ (.A0(\cb_east.inst.cb_conf_bus[123] ),
    .A1(\cb_east.inst.cb_conf_bus[124] ),
    .S(psn_net_0),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _05479_ (.A0(\cb_east.inst.cb_conf_bus[124] ),
    .A1(\cb_east.inst.cb_conf_bus[125] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _05480_ (.A0(\cb_east.inst.cb_conf_bus[125] ),
    .A1(\cb_east.inst.cb_conf_bus[126] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _05481_ (.A0(\cb_east.inst.cb_conf_bus[126] ),
    .A1(\cb_east.inst.cb_conf_bus[127] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _05482_ (.A0(\cb_east.inst.cb_conf_bus[127] ),
    .A1(\cb_east.inst.cb_conf_bus[128] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _05483_ (.A0(\cb_east.inst.cb_conf_bus[128] ),
    .A1(\cb_east.inst.cb_conf_bus[129] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _05484_ (.A0(\cb_east.inst.cb_conf_bus[129] ),
    .A1(\cb_east.inst.cb_conf_bus[130] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _05485_ (.A0(\cb_east.inst.cb_conf_bus[130] ),
    .A1(\cb_east.inst.cb_conf_bus[131] ),
    .S(psn_net_22),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _05486_ (.A0(\cb_east.inst.cb_conf_bus[131] ),
    .A1(\cb_east.inst.cb_conf_bus[132] ),
    .S(psn_net_22),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _05487_ (.A0(\cb_east.inst.cb_conf_bus[132] ),
    .A1(\cb_east.inst.cb_conf_bus[133] ),
    .S(psn_net_22),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _05488_ (.A0(\cb_east.inst.cb_conf_bus[133] ),
    .A1(\cb_east.inst.cb_conf_bus[134] ),
    .S(psn_net_20),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _05489_ (.A0(\cb_east.inst.cb_conf_bus[134] ),
    .A1(\cb_east.inst.cb_conf_bus[135] ),
    .S(psn_net_20),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _05490_ (.A0(\cb_east.inst.cb_conf_bus[135] ),
    .A1(\cb_east.inst.cb_conf_bus[136] ),
    .S(psn_net_20),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _05491_ (.A0(\cb_east.inst.cb_conf_bus[136] ),
    .A1(\cb_east.inst.cb_conf_bus[137] ),
    .S(psn_net_20),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _05492_ (.A0(\cb_east.inst.cb_conf_bus[137] ),
    .A1(\cb_east.inst.cb_conf_bus[138] ),
    .S(psn_net_20),
    .X(_02314_));
 sky130_fd_sc_hd__mux2_1 _05493_ (.A0(\cb_east.inst.cb_conf_bus[138] ),
    .A1(\cb_east.inst.cb_conf_bus[139] ),
    .S(psn_net_20),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _05494_ (.A0(\cb_east.inst.cb_conf_bus[139] ),
    .A1(\cb_east.inst.cb_conf_bus[140] ),
    .S(psn_net_20),
    .X(_02318_));
 sky130_fd_sc_hd__mux2_1 _05495_ (.A0(\cb_east.inst.cb_conf_bus[140] ),
    .A1(\cb_east.inst.cb_conf_bus[141] ),
    .S(psn_net_20),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _05496_ (.A0(\cb_east.inst.cb_conf_bus[141] ),
    .A1(\cb_east.inst.cb_conf_bus[142] ),
    .S(psn_net_20),
    .X(_02322_));
 sky130_fd_sc_hd__mux2_1 _05497_ (.A0(\cb_east.inst.cb_conf_bus[142] ),
    .A1(\cb_east.inst.cb_conf_bus[143] ),
    .S(psn_net_20),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _05498_ (.A0(\cb_east.inst.cb_conf_bus[143] ),
    .A1(\cb_east.inst.cb_conf_bus[144] ),
    .S(psn_net_20),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _05499_ (.A0(\cb_east.inst.cb_conf_bus[144] ),
    .A1(\cb_east.inst.cb_conf_bus[145] ),
    .S(psn_net_20),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _05500_ (.A0(\cb_east.inst.cb_conf_bus[145] ),
    .A1(\cb_east.inst.cb_conf_bus[146] ),
    .S(psn_net_20),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _05501_ (.A0(\cb_east.inst.cb_conf_bus[146] ),
    .A1(\cb_east.inst.cb_conf_bus[147] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _05502_ (.A0(\cb_east.inst.cb_conf_bus[147] ),
    .A1(\cb_east.inst.cb_conf_bus[148] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _05503_ (.A0(\cb_east.inst.cb_conf_bus[148] ),
    .A1(\cb_east.inst.cb_conf_bus[149] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _05504_ (.A0(\cb_east.inst.cb_conf_bus[149] ),
    .A1(\cb_east.inst.cb_conf_bus[150] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _05505_ (.A0(\cb_east.inst.cb_conf_bus[150] ),
    .A1(\cb_east.inst.cb_conf_bus[151] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02340_));
 sky130_fd_sc_hd__mux2_1 _05506_ (.A0(\cb_east.inst.cb_conf_bus[151] ),
    .A1(\cb_east.inst.cb_conf_bus[152] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _05507_ (.A0(\cb_east.inst.cb_conf_bus[152] ),
    .A1(\cb_east.inst.cb_conf_bus[153] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _05508_ (.A0(\cb_east.inst.cb_conf_bus[153] ),
    .A1(\cb_east.inst.cb_conf_bus[154] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _05509_ (.A0(\cb_east.inst.cb_conf_bus[154] ),
    .A1(\cb_east.inst.cb_conf_bus[155] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_1 _05510_ (.A0(\cb_east.inst.cb_conf_bus[155] ),
    .A1(\cb_east.inst.cb_conf_bus[156] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _05511_ (.A0(\cb_east.inst.cb_conf_bus[156] ),
    .A1(\cb_east.inst.cb_conf_bus[157] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02352_));
 sky130_fd_sc_hd__mux2_1 _05512_ (.A0(\cb_east.inst.cb_conf_bus[157] ),
    .A1(\cb_east.inst.cb_conf_bus[158] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02354_));
 sky130_fd_sc_hd__mux2_1 _05513_ (.A0(\cb_east.inst.cb_conf_bus[158] ),
    .A1(\cb_east.inst.cb_conf_bus[159] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _05514_ (.A0(\cb_east.inst.cb_conf_bus[159] ),
    .A1(\cb_east.inst.cb_conf_bus[160] ),
    .S(psn_net_19),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _05515_ (.A0(\cb_east.inst.cb_conf_bus[160] ),
    .A1(\cb_east.inst.cb_conf_bus[161] ),
    .S(psn_net_19),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _05516_ (.A0(\cb_east.inst.cb_conf_bus[161] ),
    .A1(\cb_east.inst.cb_conf_bus[162] ),
    .S(psn_net_19),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _05517_ (.A0(\cb_east.inst.cb_conf_bus[162] ),
    .A1(\cb_east.inst.cb_conf_bus[163] ),
    .S(psn_net_19),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _05518_ (.A0(\cb_east.inst.cb_conf_bus[163] ),
    .A1(\cb_east.inst.cb_conf_bus[164] ),
    .S(psn_net_19),
    .X(_02366_));
 sky130_fd_sc_hd__mux2_1 _05519_ (.A0(\cb_east.inst.cb_conf_bus[164] ),
    .A1(\cb_east.inst.cb_conf_bus[165] ),
    .S(psn_net_19),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _05520_ (.A0(\cb_east.inst.cb_conf_bus[165] ),
    .A1(\cb_east.inst.cb_conf_bus[166] ),
    .S(psn_net_19),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _05521_ (.A0(\cb_east.inst.cb_conf_bus[166] ),
    .A1(\cb_east.inst.cb_conf_bus[167] ),
    .S(psn_net_19),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _05522_ (.A0(\cb_east.inst.cb_conf_bus[167] ),
    .A1(\cb_east.inst.cb_conf_bus[168] ),
    .S(psn_net_19),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _05523_ (.A0(\cb_east.inst.cb_conf_bus[168] ),
    .A1(\cb_east.inst.cb_conf_bus[169] ),
    .S(psn_net_19),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _05524_ (.A0(\cb_east.inst.cb_conf_bus[169] ),
    .A1(\cb_east.inst.cb_conf_bus[170] ),
    .S(psn_net_19),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _05525_ (.A0(\cb_east.inst.cb_conf_bus[170] ),
    .A1(\cb_east.inst.cb_conf_bus[171] ),
    .S(psn_net_19),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _05526_ (.A0(\cb_east.inst.cb_conf_bus[171] ),
    .A1(\cb_east.inst.cb_conf_bus[172] ),
    .S(psn_net_19),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _05527_ (.A0(\cb_east.inst.cb_conf_bus[172] ),
    .A1(\cb_east.inst.cb_conf_bus[173] ),
    .S(psn_net_18),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _05528_ (.A0(\cb_east.inst.cb_conf_bus[173] ),
    .A1(\cb_east.inst.cb_conf_bus[174] ),
    .S(psn_net_18),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _05529_ (.A0(\cb_east.inst.cb_conf_bus[174] ),
    .A1(\cb_east.inst.cb_conf_bus[175] ),
    .S(psn_net_18),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _05530_ (.A0(\cb_east.inst.cb_conf_bus[175] ),
    .A1(\cb_east.inst.cb_conf_bus[176] ),
    .S(psn_net_18),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _05531_ (.A0(\cb_east.inst.cb_conf_bus[176] ),
    .A1(\cb_east.inst.cb_conf_bus[177] ),
    .S(psn_net_18),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _05532_ (.A0(\cb_east.inst.cb_conf_bus[177] ),
    .A1(\cb_east.inst.cb_conf_bus[178] ),
    .S(psn_net_18),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _05533_ (.A0(\cb_east.inst.cb_conf_bus[178] ),
    .A1(\cb_east.inst.cb_conf_bus[179] ),
    .S(psn_net_18),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _05534_ (.A0(\cb_east.inst.cb_conf_bus[179] ),
    .A1(\cb_east.inst.cb_conf_bus[180] ),
    .S(psn_net_18),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _05535_ (.A0(\cb_east.inst.cb_conf_bus[180] ),
    .A1(\cb_east.inst.cb_conf_bus[181] ),
    .S(psn_net_18),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _05536_ (.A0(\cb_east.inst.cb_conf_bus[181] ),
    .A1(\cb_east.inst.cb_conf_bus[182] ),
    .S(psn_net_14),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _05537_ (.A0(\cb_east.inst.cb_conf_bus[182] ),
    .A1(\cb_east.inst.cb_conf_bus[183] ),
    .S(psn_net_14),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _05538_ (.A0(\cb_east.inst.cb_conf_bus[183] ),
    .A1(\cb_east.inst.cb_conf_bus[184] ),
    .S(psn_net_14),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _05539_ (.A0(\cb_east.inst.cb_conf_bus[184] ),
    .A1(\cb_east.inst.cb_conf_bus[185] ),
    .S(psn_net_14),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _05540_ (.A0(\cb_east.inst.cb_conf_bus[185] ),
    .A1(\cb_east.inst.cb_conf_bus[186] ),
    .S(psn_net_14),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _05541_ (.A0(\cb_east.inst.cb_conf_bus[186] ),
    .A1(\cb_east.inst.cb_conf_bus[187] ),
    .S(psn_net_14),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _05542_ (.A0(\cb_east.inst.cb_conf_bus[187] ),
    .A1(\cb_east.inst.cb_conf_bus[188] ),
    .S(psn_net_14),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _05543_ (.A0(\cb_east.inst.cb_conf_bus[188] ),
    .A1(\cb_east.inst.cb_conf_bus[189] ),
    .S(psn_net_14),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _05544_ (.A0(\cb_east.inst.cb_conf_bus[189] ),
    .A1(\cb_east.inst.cb_conf_bus[190] ),
    .S(psn_net_14),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _05545_ (.A0(\cb_east.inst.cb_conf_bus[190] ),
    .A1(\cb_east.inst.cb_conf_bus[191] ),
    .S(psn_net_14),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _05546_ (.A0(\cb_east.inst.cb_conf_bus[191] ),
    .A1(\cb_east.inst.cb_conf_bus[192] ),
    .S(psn_net_14),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _05547_ (.A0(\cb_east.inst.cb_conf_bus[192] ),
    .A1(\cb_east.inst.cb_conf_bus[193] ),
    .S(psn_net_14),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _05548_ (.A0(\cb_east.inst.cb_conf_bus[193] ),
    .A1(\cb_east.inst.cb_conf_bus[194] ),
    .S(psn_net_14),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _05549_ (.A0(\cb_east.inst.cb_conf_bus[194] ),
    .A1(\cb_east.inst.cb_conf_bus[195] ),
    .S(psn_net_14),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _05550_ (.A0(\cb_east.inst.cb_conf_bus[195] ),
    .A1(\cb_east.inst.cb_conf_bus[196] ),
    .S(psn_net_14),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _05551_ (.A0(\cb_east.inst.cb_conf_bus[196] ),
    .A1(\cb_east.inst.cb_conf_bus[197] ),
    .S(psn_net_14),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _05552_ (.A0(\cb_east.inst.cb_conf_bus[197] ),
    .A1(\cb_east.inst.cb_conf_bus[198] ),
    .S(psn_net_14),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _05553_ (.A0(\cb_east.inst.cb_conf_bus[198] ),
    .A1(\cb_east.inst.cb_conf_bus[199] ),
    .S(psn_net_14),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _05554_ (.A0(\cb_east.inst.cb_conf_bus[199] ),
    .A1(\cb_east.inst.cb_conf_bus[200] ),
    .S(psn_net_14),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _05555_ (.A0(\cb_east.inst.cb_conf_bus[200] ),
    .A1(\cb_east.inst.cb_conf_bus[201] ),
    .S(psn_net_14),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _05556_ (.A0(\cb_east.inst.cb_conf_bus[201] ),
    .A1(\cb_east.inst.cb_conf_bus[202] ),
    .S(psn_net_14),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _05557_ (.A0(\cb_east.inst.cb_conf_bus[202] ),
    .A1(\cb_east.inst.cb_conf_bus[203] ),
    .S(psn_net_14),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _05558_ (.A0(\cb_east.inst.cb_conf_bus[203] ),
    .A1(\cb_east.inst.cb_conf_bus[204] ),
    .S(psn_net_14),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _05559_ (.A0(\cb_east.inst.cb_conf_bus[204] ),
    .A1(\cb_east.inst.cb_conf_bus[205] ),
    .S(psn_net_14),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _05560_ (.A0(\cb_east.inst.cb_conf_bus[205] ),
    .A1(\cb_east.inst.cb_conf_bus[206] ),
    .S(psn_net_14),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _05561_ (.A0(\cb_east.inst.cb_conf_bus[206] ),
    .A1(\cb_east.inst.cb_conf_bus[207] ),
    .S(psn_net_14),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _05562_ (.A0(\cb_east.inst.cb_conf_bus[207] ),
    .A1(\cb_east.inst.cb_conf_bus[208] ),
    .S(psn_net_14),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _05563_ (.A0(\cb_east.inst.cb_conf_bus[208] ),
    .A1(\cb_east.inst.cb_conf_bus[209] ),
    .S(psn_net_14),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _05564_ (.A0(\cb_east.inst.cb_conf_bus[209] ),
    .A1(\cb_east.inst.cb_conf_bus[210] ),
    .S(psn_net_14),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _05565_ (.A0(\cb_east.inst.cb_conf_bus[210] ),
    .A1(\cb_east.inst.cb_conf_bus[211] ),
    .S(psn_net_14),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _05566_ (.A0(\cb_east.inst.cb_conf_bus[211] ),
    .A1(\cb_east.inst.cb_conf_bus[212] ),
    .S(psn_net_14),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _05567_ (.A0(\cb_east.inst.cb_conf_bus[212] ),
    .A1(\cb_east.inst.cb_conf_bus[213] ),
    .S(psn_net_14),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _05568_ (.A0(\cb_east.inst.cb_conf_bus[213] ),
    .A1(\cb_east.inst.cb_conf_bus[214] ),
    .S(psn_net_14),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _05569_ (.A0(\cb_east.inst.cb_conf_bus[214] ),
    .A1(\cb_east.inst.cb_conf_bus[215] ),
    .S(psn_net_14),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _05570_ (.A0(\cb_east.inst.cb_conf_bus[215] ),
    .A1(\cb_east.inst.cb_conf_bus[216] ),
    .S(psn_net_14),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _05571_ (.A0(\cb_east.inst.cb_conf_bus[216] ),
    .A1(\cb_east.inst.cb_conf_bus[217] ),
    .S(psn_net_14),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _05572_ (.A0(\cb_east.inst.cb_conf_bus[217] ),
    .A1(\cb_east.inst.cb_conf_bus[218] ),
    .S(psn_net_14),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _05573_ (.A0(\cb_east.inst.cb_conf_bus[218] ),
    .A1(\cb_east.inst.cb_conf_bus[219] ),
    .S(psn_net_14),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _05574_ (.A0(\cb_east.inst.cb_conf_bus[219] ),
    .A1(\cb_east.inst.cb_conf_bus[220] ),
    .S(psn_net_14),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _05575_ (.A0(\cb_east.inst.cb_conf_bus[220] ),
    .A1(\cb_east.inst.cb_conf_bus[221] ),
    .S(psn_net_21),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _05576_ (.A0(\cb_east.inst.cb_conf_bus[221] ),
    .A1(\cb_east.inst.cb_conf_bus[222] ),
    .S(psn_net_21),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _05577_ (.A0(\cb_east.inst.cb_conf_bus[222] ),
    .A1(\cb_east.inst.cb_conf_bus[223] ),
    .S(psn_net_21),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _05578_ (.A0(\cb_east.inst.cb_conf_bus[223] ),
    .A1(\cb_east.inst.cb_conf_bus[224] ),
    .S(psn_net_21),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _05579_ (.A0(\cb_east.inst.cb_conf_bus[224] ),
    .A1(\cb_east.inst.cb_conf_bus[225] ),
    .S(psn_net_21),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _05580_ (.A0(\cb_east.inst.cb_conf_bus[225] ),
    .A1(\cb_east.inst.cb_conf_bus[226] ),
    .S(psn_net_21),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _05581_ (.A0(\cb_east.inst.cb_conf_bus[226] ),
    .A1(\cb_east.inst.cb_conf_bus[227] ),
    .S(psn_net_1),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _05582_ (.A0(\cb_east.inst.cb_conf_bus[227] ),
    .A1(\cb_east.inst.cb_conf_bus[228] ),
    .S(psn_net_1),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _05583_ (.A0(\cb_east.inst.cb_conf_bus[228] ),
    .A1(\cb_east.inst.cb_conf_bus[229] ),
    .S(psn_net_1),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _05584_ (.A0(\cb_east.inst.cb_conf_bus[229] ),
    .A1(\cb_east.inst.cb_conf_bus[230] ),
    .S(psn_net_1),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _05585_ (.A0(\cb_east.inst.cb_conf_bus[230] ),
    .A1(\cb_east.inst.cb_conf_bus[231] ),
    .S(psn_net_1),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _05586_ (.A0(\cb_east.inst.cb_conf_bus[231] ),
    .A1(\cb_east.inst.cb_conf_bus[232] ),
    .S(psn_net_1),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _05587_ (.A0(\cb_east.inst.cb_conf_bus[232] ),
    .A1(\cb_east.inst.cb_conf_bus[233] ),
    .S(psn_net_1),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _05588_ (.A0(\cb_east.inst.cb_conf_bus[233] ),
    .A1(\cb_east.inst.cb_conf_bus[234] ),
    .S(psn_net_1),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _05589_ (.A0(\cb_east.inst.cb_conf_bus[234] ),
    .A1(\cb_east.inst.cb_conf_bus[235] ),
    .S(psn_net_1),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _05590_ (.A0(\cb_east.inst.cb_conf_bus[235] ),
    .A1(\cb_east.inst.cb_conf_bus[236] ),
    .S(psn_net_1),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _05591_ (.A0(\cb_east.inst.cb_conf_bus[236] ),
    .A1(\cb_east.inst.cb_conf_bus[237] ),
    .S(psn_net_1),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _05592_ (.A0(\cb_east.inst.cb_conf_bus[237] ),
    .A1(\cb_east.inst.cb_conf_bus[238] ),
    .S(psn_net_1),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _05593_ (.A0(\cb_east.inst.cb_conf_bus[238] ),
    .A1(\cb_east.inst.cb_conf_bus[239] ),
    .S(psn_net_1),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _05594_ (.A0(\cb_east.inst.cb_conf_bus[239] ),
    .A1(\cb_east.inst.cb_conf_bus[240] ),
    .S(psn_net_1),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _05595_ (.A0(\cb_east.inst.cb_conf_bus[240] ),
    .A1(\cb_east.inst.cb_conf_bus[241] ),
    .S(psn_net_1),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _05596_ (.A0(\cb_east.inst.cb_conf_bus[241] ),
    .A1(\cb_east.inst.cb_conf_bus[242] ),
    .S(psn_net_1),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _05597_ (.A0(\cb_east.inst.cb_conf_bus[242] ),
    .A1(\cb_east.inst.cb_conf_bus[243] ),
    .S(psn_net_1),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _05598_ (.A0(\cb_east.inst.cb_conf_bus[243] ),
    .A1(\cb_east.inst.cb_conf_bus[244] ),
    .S(psn_net_1),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _05599_ (.A0(\cb_east.inst.cb_conf_bus[244] ),
    .A1(\cb_east.inst.cb_conf_bus[245] ),
    .S(psn_net_1),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _05600_ (.A0(\cb_east.inst.cb_conf_bus[245] ),
    .A1(\cb_east.inst.cb_conf_bus[246] ),
    .S(psn_net_1),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _05601_ (.A0(\cb_east.inst.cb_conf_bus[246] ),
    .A1(\cb_east.inst.cb_conf_bus[247] ),
    .S(psn_net_1),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _05602_ (.A0(\cb_east.inst.cb_conf_bus[247] ),
    .A1(\cb_east.inst.cb_conf_bus[248] ),
    .S(psn_net_1),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _05603_ (.A0(\cb_east.inst.cb_conf_bus[248] ),
    .A1(\cb_east.inst.cb_conf_bus[249] ),
    .S(psn_net_1),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _05604_ (.A0(\cb_east.inst.cb_conf_bus[249] ),
    .A1(\cb_east.inst.cb_conf_bus[250] ),
    .S(psn_net_1),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _05605_ (.A0(\cb_east.inst.cb_conf_bus[250] ),
    .A1(\cb_east.inst.cb_conf_bus[251] ),
    .S(psn_net_1),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _05606_ (.A0(\cb_east.inst.cb_conf_bus[251] ),
    .A1(\cb_east.inst.cb_conf_bus[252] ),
    .S(psn_net_1),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _05607_ (.A0(\cb_east.inst.cb_conf_bus[252] ),
    .A1(\cb_east.inst.cb_conf_bus[253] ),
    .S(psn_net_1),
    .X(_02544_));
 sky130_fd_sc_hd__mux2_1 _05608_ (.A0(\cb_east.inst.cb_conf_bus[253] ),
    .A1(\cb_east.inst.cb_conf_bus[254] ),
    .S(psn_net_1),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_1 _05609_ (.A0(\cb_east.inst.cb_conf_bus[254] ),
    .A1(\cb_east.inst.cb_conf_bus[255] ),
    .S(psn_net_1),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _05610_ (.A0(\cb_east.inst.cb_conf_bus[255] ),
    .A1(\cb_east.inst.cb_conf_bus[256] ),
    .S(psn_net_1),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _05611_ (.A0(\cb_east.inst.cb_conf_bus[256] ),
    .A1(\cb_east.inst.cb_conf_bus[257] ),
    .S(psn_net_1),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _05612_ (.A0(\cb_east.inst.cb_conf_bus[257] ),
    .A1(\cb_east.inst.cb_conf_bus[258] ),
    .S(psn_net_1),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _05613_ (.A0(\cb_east.inst.cb_conf_bus[258] ),
    .A1(\cb_east.inst.cb_conf_bus[259] ),
    .S(psn_net_1),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _05614_ (.A0(\cb_east.inst.cb_conf_bus[259] ),
    .A1(\cb_east.inst.cb_conf_bus[260] ),
    .S(psn_net_1),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _05615_ (.A0(\cb_east.inst.cb_conf_bus[260] ),
    .A1(\cb_east.inst.cb_conf_bus[261] ),
    .S(psn_net_15),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _05616_ (.A0(\cb_east.inst.cb_conf_bus[261] ),
    .A1(\cb_east.inst.cb_conf_bus[262] ),
    .S(psn_net_15),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _05617_ (.A0(\cb_east.inst.cb_conf_bus[262] ),
    .A1(\cb_east.inst.cb_conf_bus[263] ),
    .S(psn_net_15),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _05618_ (.A0(\cb_east.inst.cb_conf_bus[263] ),
    .A1(\cb_east.inst.cb_conf_bus[264] ),
    .S(psn_net_15),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _05619_ (.A0(\cb_east.inst.cb_conf_bus[264] ),
    .A1(\cb_east.inst.cb_conf_bus[265] ),
    .S(psn_net_15),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _05620_ (.A0(\cb_east.inst.cb_conf_bus[265] ),
    .A1(\cb_east.inst.cb_conf_bus[266] ),
    .S(psn_net_15),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _05621_ (.A0(\cb_east.inst.cb_conf_bus[266] ),
    .A1(\cb_east.inst.cb_conf_bus[267] ),
    .S(psn_net_15),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_1 _05622_ (.A0(\cb_east.inst.cb_conf_bus[267] ),
    .A1(\cb_east.inst.cb_conf_bus[268] ),
    .S(psn_net_15),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _05623_ (.A0(\cb_east.inst.cb_conf_bus[268] ),
    .A1(\cb_east.inst.cb_conf_bus[269] ),
    .S(psn_net_15),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_1 _05624_ (.A0(\cb_east.inst.cb_conf_bus[269] ),
    .A1(\cb_east.inst.cb_conf_bus[270] ),
    .S(psn_net_15),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _05625_ (.A0(\cb_east.inst.cb_conf_bus[270] ),
    .A1(\cb_east.inst.cb_conf_bus[271] ),
    .S(psn_net_15),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _05626_ (.A0(\cb_east.inst.cb_conf_bus[271] ),
    .A1(\cb_east.inst.cb_conf_bus[272] ),
    .S(psn_net_15),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _05627_ (.A0(\cb_east.inst.cb_conf_bus[272] ),
    .A1(\cb_east.inst.cb_conf_bus[273] ),
    .S(psn_net_15),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _05628_ (.A0(\cb_east.inst.cb_conf_bus[273] ),
    .A1(\cb_east.inst.cb_conf_bus[274] ),
    .S(psn_net_15),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _05629_ (.A0(\cb_east.inst.cb_conf_bus[274] ),
    .A1(\cb_east.inst.cb_conf_bus[275] ),
    .S(psn_net_15),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _05630_ (.A0(\cb_east.inst.cb_conf_bus[275] ),
    .A1(\cb_east.inst.cb_conf_bus[276] ),
    .S(psn_net_15),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _05631_ (.A0(\cb_east.inst.cb_conf_bus[276] ),
    .A1(\cb_east.inst.cb_conf_bus[277] ),
    .S(psn_net_15),
    .X(_02592_));
 sky130_fd_sc_hd__mux2_1 _05632_ (.A0(\cb_east.inst.cb_conf_bus[277] ),
    .A1(\cb_east.inst.cb_conf_bus[278] ),
    .S(psn_net_15),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _05633_ (.A0(\cb_east.inst.cb_conf_bus[278] ),
    .A1(\cb_east.inst.cb_conf_bus[279] ),
    .S(psn_net_15),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _05634_ (.A0(\cb_east.inst.cb_conf_bus[279] ),
    .A1(\cb_east.inst.cb_conf_bus[280] ),
    .S(psn_net_15),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _05635_ (.A0(\cb_east.inst.cb_conf_bus[280] ),
    .A1(\cb_east.inst.cb_conf_bus[281] ),
    .S(psn_net_15),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _05636_ (.A0(\cb_east.inst.cb_conf_bus[281] ),
    .A1(\cb_east.inst.cb_conf_bus[282] ),
    .S(psn_net_15),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _05637_ (.A0(\cb_east.inst.cb_conf_bus[282] ),
    .A1(\cb_east.inst.cb_conf_bus[283] ),
    .S(psn_net_15),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _05638_ (.A0(\cb_east.inst.cb_conf_bus[283] ),
    .A1(\cb_east.inst.cb_conf_bus[284] ),
    .S(psn_net_15),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _05639_ (.A0(\cb_east.inst.cb_conf_bus[284] ),
    .A1(\cb_east.inst.cb_conf_bus[285] ),
    .S(psn_net_15),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _05640_ (.A0(\cb_east.inst.cb_conf_bus[285] ),
    .A1(\cb_east.inst.cb_conf_bus[286] ),
    .S(psn_net_15),
    .X(_02610_));
 sky130_fd_sc_hd__mux2_1 _05641_ (.A0(\cb_east.inst.cb_conf_bus[286] ),
    .A1(\cb_east.inst.cb_conf_bus[287] ),
    .S(psn_net_15),
    .X(_02612_));
 sky130_fd_sc_hd__mux2_1 _05642_ (.A0(\cb_east.inst.cb_conf_bus[287] ),
    .A1(\cb_east.inst.cb_conf_bus[288] ),
    .S(psn_net_15),
    .X(_02614_));
 sky130_fd_sc_hd__mux2_1 _05643_ (.A0(\cb_east.inst.cb_conf_bus[288] ),
    .A1(\cb_east.inst.cb_conf_bus[289] ),
    .S(psn_net_15),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _05644_ (.A0(\cb_east.inst.cb_conf_bus[289] ),
    .A1(\cb_east.inst.cb_conf_bus[290] ),
    .S(psn_net_15),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _05645_ (.A0(\cb_east.inst.cb_conf_bus[290] ),
    .A1(\cb_east.inst.cb_conf_bus[291] ),
    .S(psn_net_15),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _05646_ (.A0(\cb_east.inst.cb_conf_bus[291] ),
    .A1(\cb_east.inst.cb_conf_bus[292] ),
    .S(psn_net_15),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _05647_ (.A0(\cb_east.inst.cb_conf_bus[292] ),
    .A1(\cb_east.inst.cb_conf_bus[293] ),
    .S(psn_net_15),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _05648_ (.A0(\cb_east.inst.cb_conf_bus[293] ),
    .A1(\cb_east.inst.cb_conf_bus[294] ),
    .S(psn_net_15),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _05649_ (.A0(\cb_east.inst.cb_conf_bus[294] ),
    .A1(\cb_east.inst.cb_conf_bus[295] ),
    .S(psn_net_15),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _05650_ (.A0(\cb_east.inst.cb_conf_bus[295] ),
    .A1(\cb_east.inst.cb_conf_bus[296] ),
    .S(psn_net_15),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _05651_ (.A0(\cb_east.inst.cb_conf_bus[296] ),
    .A1(\cb_east.inst.cb_conf_bus[297] ),
    .S(psn_net_15),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _05652_ (.A0(\cb_east.inst.cb_conf_bus[297] ),
    .A1(\cb_east.inst.cb_conf_bus[298] ),
    .S(psn_net_15),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _05653_ (.A0(\cb_east.inst.cb_conf_bus[298] ),
    .A1(\cb_east.inst.cb_conf_bus[299] ),
    .S(psn_net_15),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _05654_ (.A0(\cb_east.inst.cb_conf_bus[299] ),
    .A1(\cb_east.inst.cb_conf_bus[300] ),
    .S(psn_net_15),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _05655_ (.A0(\cb_east.inst.cb_conf_bus[300] ),
    .A1(\cb_east.inst.cb_conf_bus[301] ),
    .S(psn_net_15),
    .X(_02640_));
 sky130_fd_sc_hd__mux2_1 _05656_ (.A0(\cb_east.inst.cb_conf_bus[301] ),
    .A1(\cb_east.inst.cb_conf_bus[302] ),
    .S(psn_net_15),
    .X(_02642_));
 sky130_fd_sc_hd__mux2_1 _05657_ (.A0(\cb_east.inst.cb_conf_bus[302] ),
    .A1(\cb_east.inst.cb_conf_bus[303] ),
    .S(psn_net_15),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _05658_ (.A0(\cb_east.inst.cb_conf_bus[303] ),
    .A1(\cb_east.inst.cb_conf_bus[304] ),
    .S(psn_net_15),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _05659_ (.A0(\cb_east.inst.cb_conf_bus[304] ),
    .A1(\cb_east.inst.cb_conf_bus[305] ),
    .S(psn_net_15),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _05660_ (.A0(\cb_east.inst.cb_conf_bus[305] ),
    .A1(\cb_east.inst.cb_conf_bus[306] ),
    .S(psn_net_15),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _05661_ (.A0(\cb_east.inst.cb_conf_bus[306] ),
    .A1(\cb_east.inst.cb_conf_bus[307] ),
    .S(psn_net_15),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _05662_ (.A0(\cb_east.inst.cb_conf_bus[307] ),
    .A1(\cb_east.inst.cb_conf_bus[308] ),
    .S(psn_net_15),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _05663_ (.A0(\cb_east.inst.cb_conf_bus[308] ),
    .A1(\cb_east.inst.cb_conf_bus[309] ),
    .S(psn_net_15),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _05664_ (.A0(\cb_east.inst.cb_conf_bus[309] ),
    .A1(\cb_east.inst.cb_conf_bus[310] ),
    .S(psn_net_15),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _05665_ (.A0(\cb_east.inst.cb_conf_bus[310] ),
    .A1(\cb_east.inst.cb_conf_bus[311] ),
    .S(psn_net_15),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _05666_ (.A0(\cb_east.inst.cb_conf_bus[311] ),
    .A1(\cb_east.inst.cb_conf_bus[312] ),
    .S(psn_net_15),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _05667_ (.A0(\cb_east.inst.cb_conf_bus[312] ),
    .A1(\cb_east.inst.cb_conf_bus[313] ),
    .S(psn_net_15),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _05668_ (.A0(\cb_east.inst.cb_conf_bus[313] ),
    .A1(\cb_east.inst.cb_conf_bus[314] ),
    .S(psn_net_15),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _05669_ (.A0(\cb_east.inst.cb_conf_bus[314] ),
    .A1(\cb_east.inst.cb_conf_bus[315] ),
    .S(psn_net_15),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _05670_ (.A0(\cb_east.inst.cb_conf_bus[315] ),
    .A1(\cb_east.inst.cb_conf_bus[316] ),
    .S(psn_net_15),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _05671_ (.A0(\cb_east.inst.cb_conf_bus[316] ),
    .A1(\cb_east.inst.cb_conf_bus[317] ),
    .S(psn_net_15),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _05672_ (.A0(\cb_east.inst.cb_conf_bus[317] ),
    .A1(\cb_east.inst.cb_conf_bus[318] ),
    .S(psn_net_15),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _05673_ (.A0(\cb_east.inst.cb_conf_bus[318] ),
    .A1(\cb_east.inst.cb_conf_bus[319] ),
    .S(psn_net_15),
    .X(_02676_));
 sky130_fd_sc_hd__mux2_1 _05674_ (.A0(\cb_east.inst.cb_conf_bus[319] ),
    .A1(\cb_east.inst.cb_conf_bus[320] ),
    .S(psn_net_15),
    .X(_02678_));
 sky130_fd_sc_hd__mux2_1 _05675_ (.A0(\cb_east.inst.cb_conf_bus[320] ),
    .A1(\cb_east.inst.cb_conf_bus[321] ),
    .S(psn_net_15),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _05676_ (.A0(\cb_east.inst.cb_conf_bus[321] ),
    .A1(\cb_east.inst.cb_conf_bus[322] ),
    .S(psn_net_15),
    .X(_02682_));
 sky130_fd_sc_hd__mux2_1 _05677_ (.A0(\cb_east.inst.cb_conf_bus[322] ),
    .A1(\cb_east.inst.cb_conf_bus[323] ),
    .S(psn_net_15),
    .X(_02684_));
 sky130_fd_sc_hd__mux2_1 _05678_ (.A0(\cb_east.inst.cb_conf_bus[323] ),
    .A1(\cb_east.inst.cb_conf_bus[324] ),
    .S(psn_net_15),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _05679_ (.A0(\cb_east.inst.cb_conf_bus[324] ),
    .A1(\cb_east.inst.cb_conf_bus[325] ),
    .S(psn_net_15),
    .X(_02688_));
 sky130_fd_sc_hd__mux2_1 _05680_ (.A0(\cb_east.inst.cb_conf_bus[325] ),
    .A1(\cb_east.inst.cb_conf_bus[326] ),
    .S(psn_net_15),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _05681_ (.A0(\cb_east.inst.cb_conf_bus[326] ),
    .A1(\cb_east.inst.cb_conf_bus[327] ),
    .S(psn_net_15),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _05682_ (.A0(\cb_east.inst.cb_conf_bus[327] ),
    .A1(\cb_east.inst.cb_conf_bus[328] ),
    .S(psn_net_15),
    .X(_02694_));
 sky130_fd_sc_hd__mux2_1 _05683_ (.A0(\cb_east.inst.cb_conf_bus[328] ),
    .A1(\cb_east.inst.cb_conf_bus[329] ),
    .S(psn_net_15),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _05684_ (.A0(\cb_east.inst.cb_conf_bus[329] ),
    .A1(\cb_east.inst.cb_conf_bus[330] ),
    .S(psn_net_15),
    .X(_02698_));
 sky130_fd_sc_hd__mux2_1 _05685_ (.A0(\cb_east.inst.cb_conf_bus[330] ),
    .A1(\cb_east.inst.cb_conf_bus[331] ),
    .S(psn_net_15),
    .X(_02700_));
 sky130_fd_sc_hd__mux2_1 _05686_ (.A0(\cb_east.inst.cb_conf_bus[331] ),
    .A1(\cb_east.inst.cb_conf_bus[332] ),
    .S(psn_net_15),
    .X(_02702_));
 sky130_fd_sc_hd__mux2_1 _05687_ (.A0(\cb_east.inst.cb_conf_bus[332] ),
    .A1(\cb_east.inst.cb_conf_bus[333] ),
    .S(psn_net_15),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _05688_ (.A0(\cb_east.inst.cb_conf_bus[333] ),
    .A1(\cb_east.inst.cb_conf_bus[334] ),
    .S(psn_net_15),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _05689_ (.A0(\cb_east.inst.cb_conf_bus[334] ),
    .A1(\cb_east.inst.cb_conf_bus[335] ),
    .S(psn_net_15),
    .X(_02708_));
 sky130_fd_sc_hd__mux2_1 _05690_ (.A0(\cb_east.inst.cb_conf_bus[335] ),
    .A1(\cb_east.inst.cb_conf_bus[336] ),
    .S(psn_net_15),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _05691_ (.A0(\cb_east.inst.cb_conf_bus[336] ),
    .A1(\cb_east.inst.cb_conf_bus[337] ),
    .S(psn_net_15),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _05692_ (.A0(\cb_east.inst.cb_conf_bus[337] ),
    .A1(\cb_east.inst.cb_conf_bus[338] ),
    .S(psn_net_15),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _05693_ (.A0(\cb_east.inst.cb_conf_bus[338] ),
    .A1(\cb_east.inst.cb_conf_bus[339] ),
    .S(psn_net_15),
    .X(_02716_));
 sky130_fd_sc_hd__mux2_1 _05694_ (.A0(\cb_east.inst.cb_conf_bus[339] ),
    .A1(\cb_east.inst.cb_conf_bus[340] ),
    .S(psn_net_15),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _05695_ (.A0(\cb_east.inst.cb_conf_bus[340] ),
    .A1(\cb_east.inst.cb_conf_bus[341] ),
    .S(psn_net_15),
    .X(_02720_));
 sky130_fd_sc_hd__mux2_1 _05696_ (.A0(\cb_east.inst.cb_conf_bus[341] ),
    .A1(\cb_east.inst.cb_conf_bus[342] ),
    .S(psn_net_15),
    .X(_02722_));
 sky130_fd_sc_hd__mux2_1 _05697_ (.A0(\cb_east.inst.cb_conf_bus[342] ),
    .A1(\cb_east.inst.cb_conf_bus[343] ),
    .S(psn_net_15),
    .X(_02724_));
 sky130_fd_sc_hd__mux2_1 _05698_ (.A0(\cb_east.inst.cb_conf_bus[343] ),
    .A1(\cb_east.inst.cb_conf_bus[344] ),
    .S(psn_net_15),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _05699_ (.A0(\cb_east.inst.cb_conf_bus[344] ),
    .A1(\cb_east.inst.cb_conf_bus[345] ),
    .S(psn_net_15),
    .X(_02728_));
 sky130_fd_sc_hd__mux2_1 _05700_ (.A0(\cb_east.inst.cb_conf_bus[345] ),
    .A1(\cb_east.inst.cb_conf_bus[346] ),
    .S(psn_net_15),
    .X(_02730_));
 sky130_fd_sc_hd__mux2_1 _05701_ (.A0(\cb_east.inst.cb_conf_bus[346] ),
    .A1(\cb_east.inst.cb_conf_bus[347] ),
    .S(psn_net_15),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_1 _05702_ (.A0(\cb_east.inst.cb_conf_bus[347] ),
    .A1(\cb_east.inst.cb_conf_bus[348] ),
    .S(psn_net_15),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _05703_ (.A0(\cb_east.inst.cb_conf_bus[348] ),
    .A1(\cb_east.inst.cb_conf_bus[349] ),
    .S(psn_net_15),
    .X(_02736_));
 sky130_fd_sc_hd__mux2_1 _05704_ (.A0(\cb_east.inst.cb_conf_bus[349] ),
    .A1(\cb_east.inst.cb_conf_bus[350] ),
    .S(psn_net_15),
    .X(_02738_));
 sky130_fd_sc_hd__mux2_1 _05705_ (.A0(\cb_east.inst.cb_conf_bus[350] ),
    .A1(\cb_east.inst.cb_conf_bus[351] ),
    .S(psn_net_15),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _05706_ (.A0(\cb_east.inst.cb_conf_bus[351] ),
    .A1(\cb_east.inst.cb_conf_bus[352] ),
    .S(psn_net_15),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _05707_ (.A0(\cb_east.inst.cb_conf_bus[352] ),
    .A1(\cb_east.inst.cb_conf_bus[353] ),
    .S(psn_net_15),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _05708_ (.A0(\cb_east.inst.cb_conf_bus[353] ),
    .A1(\cb_east.inst.cb_conf_bus[354] ),
    .S(psn_net_15),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _05709_ (.A0(\cb_east.inst.cb_conf_bus[354] ),
    .A1(\cb_east.inst.cb_conf_bus[355] ),
    .S(psn_net_15),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _05710_ (.A0(\cb_east.inst.cb_conf_bus[355] ),
    .A1(\cb_east.inst.cb_conf_bus[356] ),
    .S(psn_net_15),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _05711_ (.A0(\cb_east.inst.cb_conf_bus[356] ),
    .A1(\cb_east.inst.cb_conf_bus[357] ),
    .S(psn_net_15),
    .X(_02752_));
 sky130_fd_sc_hd__mux2_1 _05712_ (.A0(\cb_east.inst.cb_conf_bus[357] ),
    .A1(\cb_east.inst.cb_conf_bus[358] ),
    .S(psn_net_15),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _05713_ (.A0(\cb_east.inst.cb_conf_bus[358] ),
    .A1(\cb_east.inst.cb_conf_bus[359] ),
    .S(psn_net_15),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _05714_ (.A0(\cb_east.inst.cb_conf_bus[359] ),
    .A1(\cb_east.inst.cb_conf_bus[360] ),
    .S(psn_net_13),
    .X(_02758_));
 sky130_fd_sc_hd__mux2_1 _05715_ (.A0(\cb_east.inst.cb_conf_bus[360] ),
    .A1(\cb_east.inst.cb_conf_bus[361] ),
    .S(psn_net_13),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _05716_ (.A0(\cb_east.inst.cb_conf_bus[361] ),
    .A1(\cb_east.inst.cb_conf_bus[362] ),
    .S(psn_net_13),
    .X(_02762_));
 sky130_fd_sc_hd__mux2_1 _05717_ (.A0(\cb_east.inst.cb_conf_bus[362] ),
    .A1(\cb_east.inst.cb_conf_bus[363] ),
    .S(psn_net_13),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _05718_ (.A0(\cb_east.inst.cb_conf_bus[363] ),
    .A1(\cb_east.inst.cb_conf_bus[364] ),
    .S(psn_net_13),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _05719_ (.A0(\cb_east.inst.cb_conf_bus[364] ),
    .A1(\cb_east.inst.cb_conf_bus[365] ),
    .S(psn_net_13),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _05720_ (.A0(\cb_east.inst.cb_conf_bus[365] ),
    .A1(\cb_east.inst.cb_conf_bus[366] ),
    .S(psn_net_13),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _05721_ (.A0(\cb_east.inst.cb_conf_bus[366] ),
    .A1(\cb_east.inst.cb_conf_bus[367] ),
    .S(psn_net_15),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _05722_ (.A0(\cb_east.inst.cb_conf_bus[367] ),
    .A1(\cb_east.inst.cb_conf_bus[368] ),
    .S(psn_net_15),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _05723_ (.A0(\cb_east.inst.cb_conf_bus[368] ),
    .A1(\cb_east.inst.cb_conf_bus[369] ),
    .S(psn_net_15),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _05724_ (.A0(\cb_east.inst.cb_conf_bus[369] ),
    .A1(\cb_east.inst.cb_conf_bus[370] ),
    .S(psn_net_15),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _05725_ (.A0(\cb_east.inst.cb_conf_bus[370] ),
    .A1(\cb_east.inst.cb_conf_bus[371] ),
    .S(psn_net_15),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _05726_ (.A0(\cb_east.inst.cb_conf_bus[371] ),
    .A1(\cb_east.inst.cb_conf_bus[372] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _05727_ (.A0(\cb_east.inst.cb_conf_bus[372] ),
    .A1(\cb_east.inst.cb_conf_bus[373] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _05728_ (.A0(\cb_east.inst.cb_conf_bus[373] ),
    .A1(\cb_east.inst.cb_conf_bus[374] ),
    .S(psn_net_13),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _05729_ (.A0(\cb_east.inst.cb_conf_bus[374] ),
    .A1(\cb_east.inst.cb_conf_bus[375] ),
    .S(psn_net_14),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _05730_ (.A0(\cb_east.inst.cb_conf_bus[375] ),
    .A1(\cb_east.inst.cb_conf_bus[376] ),
    .S(psn_net_14),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _05731_ (.A0(\cb_east.inst.cb_conf_bus[376] ),
    .A1(\cb_east.inst.cb_conf_bus[377] ),
    .S(psn_net_14),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _05732_ (.A0(\cb_east.inst.cb_conf_bus[377] ),
    .A1(\cb_east.inst.cb_conf_bus[378] ),
    .S(psn_net_14),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _05733_ (.A0(\cb_east.inst.cb_conf_bus[378] ),
    .A1(\cb_east.inst.cb_conf_bus[379] ),
    .S(psn_net_14),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _05734_ (.A0(\cb_east.inst.cb_conf_bus[379] ),
    .A1(\cb_east.inst.cb_conf_bus[380] ),
    .S(psn_net_1),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _05735_ (.A0(\cb_east.inst.cb_conf_bus[380] ),
    .A1(\cb_east.inst.cb_conf_bus[381] ),
    .S(psn_net_1),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _05736_ (.A0(\cb_east.inst.cb_conf_bus[381] ),
    .A1(\cb_east.inst.cb_conf_bus[382] ),
    .S(psn_net_1),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _05737_ (.A0(\cb_east.inst.cb_conf_bus[382] ),
    .A1(\cb_east.inst.cb_conf_bus[383] ),
    .S(psn_net_1),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _05738_ (.A0(\cb_east.inst.cb_conf_bus[383] ),
    .A1(\cb_east.inst.cb_conf_bus[384] ),
    .S(psn_net_1),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _05739_ (.A0(\cb_east.inst.cb_conf_bus[384] ),
    .A1(\cb_east.inst.cb_conf_bus[385] ),
    .S(psn_net_1),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _05740_ (.A0(\cb_east.inst.cb_conf_bus[385] ),
    .A1(\cb_east.inst.cb_conf_bus[386] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _05741_ (.A0(\cb_east.inst.cb_conf_bus[386] ),
    .A1(\cb_east.inst.cb_conf_bus[387] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _05742_ (.A0(\cb_east.inst.cb_conf_bus[387] ),
    .A1(\cb_east.inst.cb_conf_bus[388] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _05743_ (.A0(\cb_east.inst.cb_conf_bus[388] ),
    .A1(\cb_east.inst.cb_conf_bus[389] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _05744_ (.A0(\cb_east.inst.cb_conf_bus[389] ),
    .A1(\cb_east.inst.cb_conf_bus[390] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _05745_ (.A0(\cb_east.inst.cb_conf_bus[390] ),
    .A1(\cb_east.inst.cb_conf_bus[391] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _05746_ (.A0(\cb_east.inst.cb_conf_bus[391] ),
    .A1(\cb_east.inst.cb_conf_bus[392] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _05747_ (.A0(\cb_east.inst.cb_conf_bus[392] ),
    .A1(\cb_east.inst.cb_conf_bus[393] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _05748_ (.A0(\cb_east.inst.cb_conf_bus[393] ),
    .A1(\cb_east.inst.cb_conf_bus[394] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _05749_ (.A0(\cb_east.inst.cb_conf_bus[394] ),
    .A1(\cb_east.inst.cb_conf_bus[395] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _05750_ (.A0(\cb_east.inst.cb_conf_bus[395] ),
    .A1(\cb_east.inst.cb_conf_bus[396] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _05751_ (.A0(\cb_east.inst.cb_conf_bus[396] ),
    .A1(\cb_east.inst.cb_conf_bus[397] ),
    .S(psn_net_24),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _05752_ (.A0(\cb_east.inst.cb_conf_bus[397] ),
    .A1(\cb_east.inst.cb_conf_bus[398] ),
    .S(psn_net_24),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _05753_ (.A0(\cb_east.inst.cb_conf_bus[398] ),
    .A1(\cb_east.inst.cb_conf_bus[399] ),
    .S(psn_net_24),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _05754_ (.A0(\cb_east.inst.cb_conf_bus[399] ),
    .A1(\cb_east.inst.cb_conf_bus[400] ),
    .S(psn_net_24),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _05755_ (.A0(\cb_east.inst.cb_conf_bus[400] ),
    .A1(\cb_east.inst.cb_conf_bus[401] ),
    .S(psn_net_24),
    .X(_02840_));
 sky130_fd_sc_hd__mux2_1 _05756_ (.A0(\cb_east.inst.cb_conf_bus[401] ),
    .A1(\cb_east.inst.cb_conf_bus[402] ),
    .S(psn_net_24),
    .X(_02842_));
 sky130_fd_sc_hd__mux2_1 _05757_ (.A0(\cb_east.inst.cb_conf_bus[402] ),
    .A1(\cb_east.inst.cb_conf_bus[403] ),
    .S(psn_net_24),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _05758_ (.A0(\cb_east.inst.cb_conf_bus[403] ),
    .A1(\cb_east.inst.cb_conf_bus[404] ),
    .S(psn_net_1),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _05759_ (.A0(\cb_east.inst.cb_conf_bus[404] ),
    .A1(\cb_east.inst.cb_conf_bus[405] ),
    .S(psn_net_1),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _05760_ (.A0(\cb_east.inst.cb_conf_bus[405] ),
    .A1(\cb_east.inst.cb_conf_bus[406] ),
    .S(psn_net_1),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _05761_ (.A0(\cb_east.inst.cb_conf_bus[406] ),
    .A1(\cb_east.inst.cb_conf_bus[407] ),
    .S(psn_net_1),
    .X(_02852_));
 sky130_fd_sc_hd__mux2_1 _05762_ (.A0(\cb_east.inst.cb_conf_bus[407] ),
    .A1(\cb_east.inst.cb_conf_bus[408] ),
    .S(psn_net_1),
    .X(_02854_));
 sky130_fd_sc_hd__mux2_1 _05763_ (.A0(\cb_east.inst.cb_conf_bus[408] ),
    .A1(\cb_east.inst.cb_conf_bus[409] ),
    .S(psn_net_1),
    .X(_02856_));
 sky130_fd_sc_hd__mux2_1 _05764_ (.A0(\cb_east.inst.cb_conf_bus[409] ),
    .A1(\cb_east.inst.cb_conf_bus[410] ),
    .S(psn_net_1),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _05765_ (.A0(\cb_east.inst.cb_conf_bus[410] ),
    .A1(\cb_east.inst.cb_conf_bus[411] ),
    .S(psn_net_1),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _05766_ (.A0(\cb_east.inst.cb_conf_bus[411] ),
    .A1(\cb_east.inst.cb_conf_bus[412] ),
    .S(psn_net_1),
    .X(_02862_));
 sky130_fd_sc_hd__mux2_1 _05767_ (.A0(\cb_east.inst.cb_conf_bus[412] ),
    .A1(\cb_east.inst.cb_conf_bus[413] ),
    .S(psn_net_1),
    .X(_02864_));
 sky130_fd_sc_hd__mux2_1 _05768_ (.A0(\cb_east.inst.cb_conf_bus[413] ),
    .A1(\cb_east.inst.cb_conf_bus[414] ),
    .S(psn_net_1),
    .X(_02866_));
 sky130_fd_sc_hd__mux2_1 _05769_ (.A0(\cb_east.inst.cb_conf_bus[414] ),
    .A1(\cb_east.inst.cb_conf_bus[415] ),
    .S(psn_net_1),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _05770_ (.A0(\cb_east.inst.cb_conf_bus[415] ),
    .A1(\cb_east.inst.cb_conf_bus[416] ),
    .S(psn_net_21),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _05771_ (.A0(\cb_east.inst.cb_conf_bus[416] ),
    .A1(\cb_east.inst.cb_conf_bus[417] ),
    .S(psn_net_21),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _05772_ (.A0(\cb_east.inst.cb_conf_bus[417] ),
    .A1(\cb_east.inst.cb_conf_bus[418] ),
    .S(psn_net_21),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _05773_ (.A0(\cb_east.inst.cb_conf_bus[418] ),
    .A1(\cb_east.inst.cb_conf_bus[419] ),
    .S(psn_net_21),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _05774_ (.A0(\cb_east.inst.cb_conf_bus[419] ),
    .A1(\cb_east.inst.configuroni.comb_shifter.config_data[420] ),
    .S(psn_net_14),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _05775_ (.A0(\cb_east.inst.configuroni.comb_shifter.config_data[420] ),
    .A1(\cb_east.inst.configuroni.comb_shifter.config_data[421] ),
    .S(psn_net_14),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _05776_ (.A0(\sb.configuroni.comb_shifter.config_data[48] ),
    .A1(\sb.configuroni.comb_shifter.config_data[49] ),
    .S(psn_net_11),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _05777_ (.A0(\sb.configuroni.comb_config[47] ),
    .A1(\sb.configuroni.comb_shifter.config_data[48] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _05778_ (.A0(\sb.configuroni.comb_config[46] ),
    .A1(\sb.configuroni.comb_config[47] ),
    .S(psn_net_15),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _05779_ (.A0(\sb.configuroni.comb_config[45] ),
    .A1(\sb.configuroni.comb_config[46] ),
    .S(psn_net_15),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _05780_ (.A0(\sb.configuroni.comb_config[44] ),
    .A1(\sb.configuroni.comb_config[45] ),
    .S(psn_net_15),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _05781_ (.A0(\sb.configuroni.comb_config[43] ),
    .A1(\sb.configuroni.comb_config[44] ),
    .S(psn_net_15),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _05782_ (.A0(\sb.configuroni.comb_config[42] ),
    .A1(\sb.configuroni.comb_config[43] ),
    .S(psn_net_15),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _05783_ (.A0(\sb.configuroni.comb_config[41] ),
    .A1(\sb.configuroni.comb_config[42] ),
    .S(psn_net_15),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _05784_ (.A0(\sb.configuroni.comb_config[40] ),
    .A1(\sb.configuroni.comb_config[41] ),
    .S(psn_net_15),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _05785_ (.A0(\sb.configuroni.comb_config[39] ),
    .A1(\sb.configuroni.comb_config[40] ),
    .S(psn_net_15),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _05786_ (.A0(\sb.configuroni.comb_config[38] ),
    .A1(\sb.configuroni.comb_config[39] ),
    .S(psn_net_15),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _05787_ (.A0(\sb.configuroni.comb_config[37] ),
    .A1(\sb.configuroni.comb_config[38] ),
    .S(psn_net_15),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _05788_ (.A0(\sb.configuroni.comb_config[36] ),
    .A1(\sb.configuroni.comb_config[37] ),
    .S(psn_net_15),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _05789_ (.A0(\sb.configuroni.comb_config[35] ),
    .A1(\sb.configuroni.comb_config[36] ),
    .S(psn_net_15),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _05790_ (.A0(\sb.configuroni.comb_config[34] ),
    .A1(\sb.configuroni.comb_config[35] ),
    .S(psn_net_15),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _05791_ (.A0(\sb.configuroni.comb_config[33] ),
    .A1(\sb.configuroni.comb_config[34] ),
    .S(psn_net_15),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _05792_ (.A0(\sb.configuroni.comb_config[32] ),
    .A1(\sb.configuroni.comb_config[33] ),
    .S(psn_net_15),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _05793_ (.A0(\sb.configuroni.comb_config[31] ),
    .A1(\sb.configuroni.comb_config[32] ),
    .S(psn_net_15),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _05794_ (.A0(\sb.configuroni.comb_config[30] ),
    .A1(\sb.configuroni.comb_config[31] ),
    .S(psn_net_15),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _05795_ (.A0(\sb.configuroni.comb_config[29] ),
    .A1(\sb.configuroni.comb_config[30] ),
    .S(psn_net_15),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _05796_ (.A0(\sb.configuroni.comb_config[28] ),
    .A1(\sb.configuroni.comb_config[29] ),
    .S(psn_net_15),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _05797_ (.A0(\sb.configuroni.comb_config[27] ),
    .A1(\sb.configuroni.comb_config[28] ),
    .S(psn_net_15),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _05798_ (.A0(\sb.configuroni.comb_config[26] ),
    .A1(\sb.configuroni.comb_config[27] ),
    .S(psn_net_15),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _05799_ (.A0(\sb.configuroni.comb_config[25] ),
    .A1(\sb.configuroni.comb_config[26] ),
    .S(psn_net_15),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _05800_ (.A0(\sb.configuroni.comb_config[24] ),
    .A1(\sb.configuroni.comb_config[25] ),
    .S(psn_net_15),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _05801_ (.A0(\sb.configuroni.comb_config[23] ),
    .A1(\sb.configuroni.comb_config[24] ),
    .S(psn_net_15),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _05802_ (.A0(\sb.configuroni.comb_config[22] ),
    .A1(\sb.configuroni.comb_config[23] ),
    .S(psn_net_16),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _05803_ (.A0(\sb.configuroni.comb_config[21] ),
    .A1(\sb.configuroni.comb_config[22] ),
    .S(psn_net_12),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _05804_ (.A0(\sb.configuroni.comb_config[20] ),
    .A1(\sb.configuroni.comb_config[21] ),
    .S(psn_net_12),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _05805_ (.A0(\sb.configuroni.comb_config[19] ),
    .A1(\sb.configuroni.comb_config[20] ),
    .S(psn_net_12),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _05806_ (.A0(\sb.configuroni.comb_config[18] ),
    .A1(\sb.configuroni.comb_config[19] ),
    .S(psn_net_11),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _05807_ (.A0(\sb.configuroni.comb_config[17] ),
    .A1(\sb.configuroni.comb_config[18] ),
    .S(psn_net_11),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _05808_ (.A0(\sb.configuroni.comb_config[16] ),
    .A1(\sb.configuroni.comb_config[17] ),
    .S(psn_net_11),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _05809_ (.A0(\sb.configuroni.comb_config[15] ),
    .A1(\sb.configuroni.comb_config[16] ),
    .S(psn_net_11),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _05810_ (.A0(\sb.configuroni.comb_config[14] ),
    .A1(\sb.configuroni.comb_config[15] ),
    .S(psn_net_11),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _05811_ (.A0(\sb.configuroni.comb_config[13] ),
    .A1(\sb.configuroni.comb_config[14] ),
    .S(psn_net_11),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _05812_ (.A0(\sb.configuroni.comb_config[12] ),
    .A1(\sb.configuroni.comb_config[13] ),
    .S(psn_net_11),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _05813_ (.A0(\sb.configuroni.comb_config[11] ),
    .A1(\sb.configuroni.comb_config[12] ),
    .S(psn_net_11),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _05814_ (.A0(\sb.configuroni.comb_config[10] ),
    .A1(\sb.configuroni.comb_config[11] ),
    .S(psn_net_11),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _05815_ (.A0(\sb.configuroni.comb_config[9] ),
    .A1(\sb.configuroni.comb_config[10] ),
    .S(psn_net_11),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _05816_ (.A0(\sb.configuroni.comb_config[8] ),
    .A1(\sb.configuroni.comb_config[9] ),
    .S(psn_net_11),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _05817_ (.A0(\sb.configuroni.comb_config[7] ),
    .A1(\sb.configuroni.comb_config[8] ),
    .S(psn_net_11),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _05818_ (.A0(\sb.configuroni.comb_config[6] ),
    .A1(\sb.configuroni.comb_config[7] ),
    .S(psn_net_11),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _05819_ (.A0(\sb.configuroni.comb_config[5] ),
    .A1(\sb.configuroni.comb_config[6] ),
    .S(psn_net_11),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _05820_ (.A0(\sb.configuroni.comb_config[4] ),
    .A1(\sb.configuroni.comb_config[5] ),
    .S(psn_net_11),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _05821_ (.A0(\sb.configuroni.comb_config[3] ),
    .A1(\sb.configuroni.comb_config[4] ),
    .S(psn_net_11),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _05822_ (.A0(\sb.configuroni.comb_config[2] ),
    .A1(\sb.configuroni.comb_config[3] ),
    .S(psn_net_11),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _05823_ (.A0(\sb.configuroni.comb_config[1] ),
    .A1(\sb.configuroni.comb_config[2] ),
    .S(psn_net_11),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _05824_ (.A0(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .A1(\sb.configuroni.comb_config[1] ),
    .S(psn_net_11),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _05825_ (.A0(\sb.configuroni.comb_shifter.config_data[49] ),
    .A1(\cb_north.inst.cb_conf_bus[0] ),
    .S(psn_net_11),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _05826_ (.A0(\slice.configuroni.mem_ctrl ),
    .A1(\slice.configuroni.comb_shifter.config_data[135] ),
    .S(set_out_hard),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _05827_ (.A0(\slice.configuroni.input_mux ),
    .A1(\slice.configuroni.comb_shifter.config_data[136] ),
    .S(set_out_hard),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _05828_ (.A0(\slice.configuroni.comb_shifter.config_data[135] ),
    .A1(\slice.configuroni.comb_shifter.config_data[136] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _05829_ (.A0(\slice.configuroni.comb_config[134] ),
    .A1(\slice.configuroni.comb_shifter.config_data[135] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _05830_ (.A0(\slice.configuroni.comb_config[133] ),
    .A1(\slice.configuroni.comb_config[134] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _05831_ (.A0(\slice.configuroni.comb_config[132] ),
    .A1(\slice.configuroni.comb_config[133] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _05832_ (.A0(\slice.configuroni.comb_config[131] ),
    .A1(\slice.configuroni.comb_config[132] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _05833_ (.A0(\slice.configuroni.comb_config[130] ),
    .A1(\slice.configuroni.comb_config[131] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _05834_ (.A0(\slice.configuroni.comb_config[129] ),
    .A1(\slice.configuroni.comb_config[130] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _05835_ (.A0(\slice.configuroni.comb_config[128] ),
    .A1(\slice.configuroni.comb_config[129] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _05836_ (.A0(\slice.configuroni.comb_config[127] ),
    .A1(\slice.configuroni.comb_config[128] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _05837_ (.A0(\slice.configuroni.comb_config[126] ),
    .A1(\slice.configuroni.comb_config[127] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _05838_ (.A0(\slice.configuroni.comb_config[125] ),
    .A1(\slice.configuroni.comb_config[126] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _05839_ (.A0(\slice.configuroni.comb_config[124] ),
    .A1(\slice.configuroni.comb_config[125] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _05840_ (.A0(\slice.configuroni.comb_config[123] ),
    .A1(\slice.configuroni.comb_config[124] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _05841_ (.A0(\slice.configuroni.comb_config[122] ),
    .A1(\slice.configuroni.comb_config[123] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _05842_ (.A0(\slice.configuroni.comb_config[121] ),
    .A1(\slice.configuroni.comb_config[122] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _05843_ (.A0(\slice.configuroni.comb_config[120] ),
    .A1(\slice.configuroni.comb_config[121] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _05844_ (.A0(\slice.configuroni.comb_config[119] ),
    .A1(\slice.configuroni.comb_config[120] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _05845_ (.A0(\slice.configuroni.comb_config[118] ),
    .A1(\slice.configuroni.comb_config[119] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _05846_ (.A0(\slice.configuroni.comb_config[117] ),
    .A1(\slice.configuroni.comb_config[118] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _05847_ (.A0(\slice.configuroni.comb_config[116] ),
    .A1(\slice.configuroni.comb_config[117] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_1 _05848_ (.A0(\slice.configuroni.comb_config[115] ),
    .A1(\slice.configuroni.comb_config[116] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _05849_ (.A0(\slice.configuroni.comb_config[114] ),
    .A1(\slice.configuroni.comb_config[115] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _05850_ (.A0(\slice.configuroni.comb_config[113] ),
    .A1(\slice.configuroni.comb_config[114] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03030_));
 sky130_fd_sc_hd__mux2_1 _05851_ (.A0(\slice.configuroni.comb_config[112] ),
    .A1(\slice.configuroni.comb_config[113] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03032_));
 sky130_fd_sc_hd__mux2_1 _05852_ (.A0(\slice.configuroni.comb_config[111] ),
    .A1(\slice.configuroni.comb_config[112] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _05853_ (.A0(\slice.configuroni.comb_config[110] ),
    .A1(\slice.configuroni.comb_config[111] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03036_));
 sky130_fd_sc_hd__mux2_1 _05854_ (.A0(\slice.configuroni.comb_config[109] ),
    .A1(\slice.configuroni.comb_config[110] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _05855_ (.A0(\slice.configuroni.comb_config[108] ),
    .A1(\slice.configuroni.comb_config[109] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _05856_ (.A0(\slice.configuroni.comb_config[107] ),
    .A1(\slice.configuroni.comb_config[108] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _05857_ (.A0(\slice.configuroni.comb_config[106] ),
    .A1(\slice.configuroni.comb_config[107] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _05858_ (.A0(\slice.configuroni.comb_config[105] ),
    .A1(\slice.configuroni.comb_config[106] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03046_));
 sky130_fd_sc_hd__mux2_1 _05859_ (.A0(\slice.configuroni.comb_config[104] ),
    .A1(\slice.configuroni.comb_config[105] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _05860_ (.A0(\slice.configuroni.comb_config[103] ),
    .A1(\slice.configuroni.comb_config[104] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03050_));
 sky130_fd_sc_hd__mux2_1 _05861_ (.A0(\slice.configuroni.comb_config[102] ),
    .A1(\slice.configuroni.comb_config[103] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03052_));
 sky130_fd_sc_hd__mux2_1 _05862_ (.A0(\slice.configuroni.comb_config[101] ),
    .A1(\slice.configuroni.comb_config[102] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03054_));
 sky130_fd_sc_hd__mux2_1 _05863_ (.A0(\slice.configuroni.comb_config[100] ),
    .A1(\slice.configuroni.comb_config[101] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03056_));
 sky130_fd_sc_hd__mux2_1 _05864_ (.A0(\slice.configuroni.comb_config[99] ),
    .A1(\slice.configuroni.comb_config[100] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03058_));
 sky130_fd_sc_hd__mux2_1 _05865_ (.A0(\slice.configuroni.comb_config[98] ),
    .A1(\slice.configuroni.comb_config[99] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _05866_ (.A0(\slice.configuroni.comb_config[97] ),
    .A1(\slice.configuroni.comb_config[98] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _05867_ (.A0(\slice.configuroni.comb_config[96] ),
    .A1(\slice.configuroni.comb_config[97] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _05868_ (.A0(\slice.configuroni.comb_config[95] ),
    .A1(\slice.configuroni.comb_config[96] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03066_));
 sky130_fd_sc_hd__mux2_1 _05869_ (.A0(\slice.configuroni.comb_config[94] ),
    .A1(\slice.configuroni.comb_config[95] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _05870_ (.A0(\slice.configuroni.comb_config[93] ),
    .A1(\slice.configuroni.comb_config[94] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _05871_ (.A0(\slice.configuroni.comb_config[92] ),
    .A1(\slice.configuroni.comb_config[93] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _05872_ (.A0(\slice.configuroni.comb_config[91] ),
    .A1(\slice.configuroni.comb_config[92] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _05873_ (.A0(\slice.configuroni.comb_config[90] ),
    .A1(\slice.configuroni.comb_config[91] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _05874_ (.A0(\slice.configuroni.comb_config[89] ),
    .A1(\slice.configuroni.comb_config[90] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _05875_ (.A0(\slice.configuroni.comb_config[88] ),
    .A1(\slice.configuroni.comb_config[89] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _05876_ (.A0(\slice.configuroni.comb_config[87] ),
    .A1(\slice.configuroni.comb_config[88] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _05877_ (.A0(\slice.configuroni.comb_config[86] ),
    .A1(\slice.configuroni.comb_config[87] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _05878_ (.A0(\slice.configuroni.comb_config[85] ),
    .A1(\slice.configuroni.comb_config[86] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _05879_ (.A0(\slice.configuroni.comb_config[84] ),
    .A1(\slice.configuroni.comb_config[85] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _05880_ (.A0(\slice.configuroni.comb_config[83] ),
    .A1(\slice.configuroni.comb_config[84] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _05881_ (.A0(\slice.configuroni.comb_config[82] ),
    .A1(\slice.configuroni.comb_config[83] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _05882_ (.A0(\slice.configuroni.comb_config[81] ),
    .A1(\slice.configuroni.comb_config[82] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _05883_ (.A0(\slice.configuroni.comb_config[80] ),
    .A1(\slice.configuroni.comb_config[81] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _05884_ (.A0(\slice.configuroni.comb_config[79] ),
    .A1(\slice.configuroni.comb_config[80] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _05885_ (.A0(\slice.configuroni.comb_config[78] ),
    .A1(\slice.configuroni.comb_config[79] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_1 _05886_ (.A0(\slice.configuroni.comb_config[77] ),
    .A1(\slice.configuroni.comb_config[78] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _05887_ (.A0(\slice.configuroni.comb_config[76] ),
    .A1(\slice.configuroni.comb_config[77] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _05888_ (.A0(\slice.configuroni.comb_config[75] ),
    .A1(\slice.configuroni.comb_config[76] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _05889_ (.A0(\slice.configuroni.comb_config[74] ),
    .A1(\slice.configuroni.comb_config[75] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03108_));
 sky130_fd_sc_hd__mux2_1 _05890_ (.A0(\slice.configuroni.comb_config[73] ),
    .A1(\slice.configuroni.comb_config[74] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03110_));
 sky130_fd_sc_hd__mux2_1 _05891_ (.A0(\slice.configuroni.comb_config[72] ),
    .A1(\slice.configuroni.comb_config[73] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03112_));
 sky130_fd_sc_hd__mux2_1 _05892_ (.A0(\slice.configuroni.comb_config[71] ),
    .A1(\slice.configuroni.comb_config[72] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _05893_ (.A0(\slice.configuroni.comb_config[70] ),
    .A1(\slice.configuroni.comb_config[71] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _05894_ (.A0(\slice.configuroni.comb_config[69] ),
    .A1(\slice.configuroni.comb_config[70] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03118_));
 sky130_fd_sc_hd__mux2_1 _05895_ (.A0(\slice.configuroni.comb_config[68] ),
    .A1(\slice.configuroni.comb_config[69] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03120_));
 sky130_fd_sc_hd__mux2_1 _05896_ (.A0(\slice.configuroni.comb_config[67] ),
    .A1(\slice.configuroni.comb_config[68] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _05897_ (.A0(\slice.configuroni.comb_config[66] ),
    .A1(\slice.configuroni.comb_config[67] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _05898_ (.A0(\slice.configuroni.comb_config[65] ),
    .A1(\slice.configuroni.comb_config[66] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _05899_ (.A0(\slice.configuroni.comb_config[64] ),
    .A1(\slice.configuroni.comb_config[65] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _05900_ (.A0(\slice.configuroni.comb_config[63] ),
    .A1(\slice.configuroni.comb_config[64] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _05901_ (.A0(\slice.configuroni.comb_config[62] ),
    .A1(\slice.configuroni.comb_config[63] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _05902_ (.A0(\slice.configuroni.comb_config[61] ),
    .A1(\slice.configuroni.comb_config[62] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_1 _05903_ (.A0(\slice.configuroni.comb_config[60] ),
    .A1(\slice.configuroni.comb_config[61] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _05904_ (.A0(\slice.configuroni.comb_config[59] ),
    .A1(\slice.configuroni.comb_config[60] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _05905_ (.A0(\slice.configuroni.comb_config[58] ),
    .A1(\slice.configuroni.comb_config[59] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_1 _05906_ (.A0(\slice.configuroni.comb_config[57] ),
    .A1(\slice.configuroni.comb_config[58] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03142_));
 sky130_fd_sc_hd__mux2_1 _05907_ (.A0(\slice.configuroni.comb_config[56] ),
    .A1(\slice.configuroni.comb_config[57] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _05908_ (.A0(\slice.configuroni.comb_config[55] ),
    .A1(\slice.configuroni.comb_config[56] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _05909_ (.A0(\slice.configuroni.comb_config[54] ),
    .A1(\slice.configuroni.comb_config[55] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _05910_ (.A0(\slice.configuroni.comb_config[53] ),
    .A1(\slice.configuroni.comb_config[54] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_1 _05911_ (.A0(\slice.configuroni.comb_config[52] ),
    .A1(\slice.configuroni.comb_config[53] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _05912_ (.A0(\slice.configuroni.comb_config[51] ),
    .A1(\slice.configuroni.comb_config[52] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03154_));
 sky130_fd_sc_hd__mux2_1 _05913_ (.A0(\slice.configuroni.comb_config[50] ),
    .A1(\slice.configuroni.comb_config[51] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03156_));
 sky130_fd_sc_hd__mux2_1 _05914_ (.A0(\slice.configuroni.comb_config[49] ),
    .A1(\slice.configuroni.comb_config[50] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03158_));
 sky130_fd_sc_hd__mux2_1 _05915_ (.A0(\slice.configuroni.comb_config[48] ),
    .A1(\slice.configuroni.comb_config[49] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03160_));
 sky130_fd_sc_hd__mux2_1 _05916_ (.A0(\slice.configuroni.comb_config[47] ),
    .A1(\slice.configuroni.comb_config[48] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03162_));
 sky130_fd_sc_hd__mux2_1 _05917_ (.A0(\slice.configuroni.comb_config[46] ),
    .A1(\slice.configuroni.comb_config[47] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03164_));
 sky130_fd_sc_hd__mux2_1 _05918_ (.A0(\slice.configuroni.comb_config[45] ),
    .A1(\slice.configuroni.comb_config[46] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03166_));
 sky130_fd_sc_hd__mux2_1 _05919_ (.A0(\slice.configuroni.comb_config[44] ),
    .A1(\slice.configuroni.comb_config[45] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03168_));
 sky130_fd_sc_hd__mux2_1 _05920_ (.A0(\slice.configuroni.comb_config[43] ),
    .A1(\slice.configuroni.comb_config[44] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03170_));
 sky130_fd_sc_hd__mux2_1 _05921_ (.A0(\slice.configuroni.comb_config[42] ),
    .A1(\slice.configuroni.comb_config[43] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03172_));
 sky130_fd_sc_hd__mux2_1 _05922_ (.A0(\slice.configuroni.comb_config[41] ),
    .A1(\slice.configuroni.comb_config[42] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _05923_ (.A0(\slice.configuroni.comb_config[40] ),
    .A1(\slice.configuroni.comb_config[41] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03176_));
 sky130_fd_sc_hd__mux2_1 _05924_ (.A0(\slice.configuroni.comb_config[39] ),
    .A1(\slice.configuroni.comb_config[40] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03178_));
 sky130_fd_sc_hd__mux2_1 _05925_ (.A0(\slice.configuroni.comb_config[38] ),
    .A1(\slice.configuroni.comb_config[39] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _05926_ (.A0(\slice.configuroni.comb_config[37] ),
    .A1(\slice.configuroni.comb_config[38] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _05927_ (.A0(\slice.configuroni.comb_config[36] ),
    .A1(\slice.configuroni.comb_config[37] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _05928_ (.A0(\slice.configuroni.comb_config[35] ),
    .A1(\slice.configuroni.comb_config[36] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03186_));
 sky130_fd_sc_hd__mux2_1 _05929_ (.A0(\slice.configuroni.comb_config[34] ),
    .A1(\slice.configuroni.comb_config[35] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _05930_ (.A0(\slice.configuroni.comb_config[33] ),
    .A1(\slice.configuroni.comb_config[34] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _05931_ (.A0(\slice.configuroni.comb_config[32] ),
    .A1(\slice.configuroni.comb_config[33] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03192_));
 sky130_fd_sc_hd__mux2_1 _05932_ (.A0(\slice.configuroni.comb_config[31] ),
    .A1(\slice.configuroni.comb_config[32] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _05933_ (.A0(\slice.configuroni.comb_config[30] ),
    .A1(\slice.configuroni.comb_config[31] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _05934_ (.A0(\slice.configuroni.comb_config[29] ),
    .A1(\slice.configuroni.comb_config[30] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _05935_ (.A0(\slice.configuroni.comb_config[28] ),
    .A1(\slice.configuroni.comb_config[29] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03200_));
 sky130_fd_sc_hd__mux2_1 _05936_ (.A0(\slice.configuroni.comb_config[27] ),
    .A1(\slice.configuroni.comb_config[28] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03202_));
 sky130_fd_sc_hd__mux2_1 _05937_ (.A0(\slice.configuroni.comb_config[26] ),
    .A1(\slice.configuroni.comb_config[27] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_1 _05938_ (.A0(\slice.configuroni.comb_config[25] ),
    .A1(\slice.configuroni.comb_config[26] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03206_));
 sky130_fd_sc_hd__mux2_1 _05939_ (.A0(\slice.configuroni.comb_config[24] ),
    .A1(\slice.configuroni.comb_config[25] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03208_));
 sky130_fd_sc_hd__mux2_1 _05940_ (.A0(\slice.configuroni.comb_config[23] ),
    .A1(\slice.configuroni.comb_config[24] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _05941_ (.A0(\slice.configuroni.comb_config[22] ),
    .A1(\slice.configuroni.comb_config[23] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _05942_ (.A0(\slice.configuroni.comb_config[21] ),
    .A1(\slice.configuroni.comb_config[22] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _05943_ (.A0(\slice.configuroni.comb_config[20] ),
    .A1(\slice.configuroni.comb_config[21] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _05944_ (.A0(\slice.configuroni.comb_config[19] ),
    .A1(\slice.configuroni.comb_config[20] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _05945_ (.A0(\slice.configuroni.comb_config[18] ),
    .A1(\slice.configuroni.comb_config[19] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _05946_ (.A0(\slice.configuroni.comb_config[17] ),
    .A1(\slice.configuroni.comb_config[18] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _05947_ (.A0(\slice.configuroni.comb_config[16] ),
    .A1(\slice.configuroni.comb_config[17] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _05948_ (.A0(\slice.configuroni.comb_config[15] ),
    .A1(\slice.configuroni.comb_config[16] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _05949_ (.A0(\slice.configuroni.comb_config[14] ),
    .A1(\slice.configuroni.comb_config[15] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_1 _05950_ (.A0(\slice.configuroni.comb_config[13] ),
    .A1(\slice.configuroni.comb_config[14] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _05951_ (.A0(\slice.configuroni.comb_config[12] ),
    .A1(\slice.configuroni.comb_config[13] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _05952_ (.A0(\slice.configuroni.comb_config[11] ),
    .A1(\slice.configuroni.comb_config[12] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _05953_ (.A0(\slice.configuroni.comb_config[10] ),
    .A1(\slice.configuroni.comb_config[11] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_1 _05954_ (.A0(\slice.configuroni.comb_config[9] ),
    .A1(\slice.configuroni.comb_config[10] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _05955_ (.A0(\slice.configuroni.comb_config[8] ),
    .A1(\slice.configuroni.comb_config[9] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _05956_ (.A0(\slice.configuroni.comb_config[7] ),
    .A1(\slice.configuroni.comb_config[8] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_1 _05957_ (.A0(\slice.configuroni.comb_config[6] ),
    .A1(\slice.configuroni.comb_config[7] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _05958_ (.A0(\slice.configuroni.comb_config[5] ),
    .A1(\slice.configuroni.comb_config[6] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _05959_ (.A0(\slice.configuroni.comb_config[4] ),
    .A1(\slice.configuroni.comb_config[5] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03248_));
 sky130_fd_sc_hd__mux2_1 _05960_ (.A0(\slice.configuroni.comb_config[3] ),
    .A1(\slice.configuroni.comb_config[4] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_1 _05961_ (.A0(\slice.configuroni.comb_config[2] ),
    .A1(\slice.configuroni.comb_config[3] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03252_));
 sky130_fd_sc_hd__mux2_1 _05962_ (.A0(\slice.configuroni.comb_config[1] ),
    .A1(\slice.configuroni.comb_config[2] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _05963_ (.A0(\slice.configuroni.comb_config[0] ),
    .A1(\slice.configuroni.comb_config[1] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03256_));
 sky130_fd_sc_hd__mux2_1 _05964_ (.A0(\slice.configuroni.comb_shifter.config_data[136] ),
    .A1(\slice.configuroni.comb_shifter.head_bit.shift_in ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_1 _05965_ (.A0(\slice.configuroni.mem_config[6] ),
    .A1(\slice.configuroni.mem_config[7] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03260_));
 sky130_fd_sc_hd__mux2_1 _05966_ (.A0(\slice.configuroni.mem_config[5] ),
    .A1(\slice.configuroni.mem_config[6] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03262_));
 sky130_fd_sc_hd__mux2_1 _05967_ (.A0(\slice.configuroni.mem_config[4] ),
    .A1(\slice.configuroni.mem_config[5] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03264_));
 sky130_fd_sc_hd__mux2_1 _05968_ (.A0(\slice.configuroni.mem_config[3] ),
    .A1(\slice.configuroni.mem_config[4] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03266_));
 sky130_fd_sc_hd__mux2_1 _05969_ (.A0(\slice.configuroni.mem_config[2] ),
    .A1(\slice.configuroni.mem_config[3] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03268_));
 sky130_fd_sc_hd__mux2_1 _05970_ (.A0(\slice.configuroni.mem_config[1] ),
    .A1(\slice.configuroni.mem_config[2] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03270_));
 sky130_fd_sc_hd__mux2_1 _05971_ (.A0(\cb_north.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .A1(\slice.configuroni.mem_config[1] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03272_));
 sky130_fd_sc_hd__mux2_1 _05972_ (.A0(\slice.configuroni.mem_config[7] ),
    .A1(\slice.configuroni.comb_config[0] ),
    .S(\slice.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03274_));
 sky130_fd_sc_hd__mux2_1 _05973_ (.A0(\cb_north.inst.configuroni.comb_shifter.config_data[421] ),
    .A1(\cb_north.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .S(psn_net_3),
    .X(_03276_));
 sky130_fd_sc_hd__mux2_1 _05974_ (.A0(\cb_north.inst.cb_conf_bus[0] ),
    .A1(\cb_north.inst.cb_conf_bus[1] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03278_));
 sky130_fd_sc_hd__mux2_1 _05975_ (.A0(\cb_north.inst.cb_conf_bus[1] ),
    .A1(\cb_north.inst.cb_conf_bus[2] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _05976_ (.A0(\cb_north.inst.cb_conf_bus[2] ),
    .A1(\cb_north.inst.cb_conf_bus[3] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _05977_ (.A0(\cb_north.inst.cb_conf_bus[3] ),
    .A1(\cb_north.inst.cb_conf_bus[4] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _05978_ (.A0(\cb_north.inst.cb_conf_bus[4] ),
    .A1(\cb_north.inst.cb_conf_bus[5] ),
    .S(psn_net_6),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _05979_ (.A0(\cb_north.inst.cb_conf_bus[5] ),
    .A1(\cb_north.inst.cb_conf_bus[6] ),
    .S(psn_net_6),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _05980_ (.A0(\cb_north.inst.cb_conf_bus[6] ),
    .A1(\cb_north.inst.cb_conf_bus[7] ),
    .S(psn_net_6),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _05981_ (.A0(\cb_north.inst.cb_conf_bus[7] ),
    .A1(\cb_north.inst.cb_conf_bus[8] ),
    .S(psn_net_6),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _05982_ (.A0(\cb_north.inst.cb_conf_bus[8] ),
    .A1(\cb_north.inst.cb_conf_bus[9] ),
    .S(psn_net_6),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _05983_ (.A0(\cb_north.inst.cb_conf_bus[9] ),
    .A1(\cb_north.inst.cb_conf_bus[10] ),
    .S(psn_net_5),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _05984_ (.A0(\cb_north.inst.cb_conf_bus[10] ),
    .A1(\cb_north.inst.cb_conf_bus[11] ),
    .S(psn_net_8),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _05985_ (.A0(\cb_north.inst.cb_conf_bus[11] ),
    .A1(\cb_north.inst.cb_conf_bus[12] ),
    .S(psn_net_3),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _05986_ (.A0(\cb_north.inst.cb_conf_bus[12] ),
    .A1(\cb_north.inst.cb_conf_bus[13] ),
    .S(psn_net_3),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _05987_ (.A0(\cb_north.inst.cb_conf_bus[13] ),
    .A1(\cb_north.inst.cb_conf_bus[14] ),
    .S(psn_net_3),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _05988_ (.A0(\cb_north.inst.cb_conf_bus[14] ),
    .A1(\cb_north.inst.cb_conf_bus[15] ),
    .S(psn_net_3),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _05989_ (.A0(\cb_north.inst.cb_conf_bus[15] ),
    .A1(\cb_north.inst.cb_conf_bus[16] ),
    .S(psn_net_3),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _05990_ (.A0(\cb_north.inst.cb_conf_bus[16] ),
    .A1(\cb_north.inst.cb_conf_bus[17] ),
    .S(psn_net_3),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _05991_ (.A0(\cb_north.inst.cb_conf_bus[17] ),
    .A1(\cb_north.inst.cb_conf_bus[18] ),
    .S(psn_net_3),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _05992_ (.A0(\cb_north.inst.cb_conf_bus[18] ),
    .A1(\cb_north.inst.cb_conf_bus[19] ),
    .S(psn_net_3),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _05993_ (.A0(\cb_north.inst.cb_conf_bus[19] ),
    .A1(\cb_north.inst.cb_conf_bus[20] ),
    .S(psn_net_3),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _05994_ (.A0(\cb_north.inst.cb_conf_bus[20] ),
    .A1(\cb_north.inst.cb_conf_bus[21] ),
    .S(psn_net_3),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _05995_ (.A0(\cb_north.inst.cb_conf_bus[21] ),
    .A1(\cb_north.inst.cb_conf_bus[22] ),
    .S(psn_net_3),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _05996_ (.A0(\cb_north.inst.cb_conf_bus[22] ),
    .A1(\cb_north.inst.cb_conf_bus[23] ),
    .S(psn_net_3),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _05997_ (.A0(\cb_north.inst.cb_conf_bus[23] ),
    .A1(\cb_north.inst.cb_conf_bus[24] ),
    .S(psn_net_3),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _05998_ (.A0(\cb_north.inst.cb_conf_bus[24] ),
    .A1(\cb_north.inst.cb_conf_bus[25] ),
    .S(psn_net_9),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _05999_ (.A0(\cb_north.inst.cb_conf_bus[25] ),
    .A1(\cb_north.inst.cb_conf_bus[26] ),
    .S(psn_net_8),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _06000_ (.A0(\cb_north.inst.cb_conf_bus[26] ),
    .A1(\cb_north.inst.cb_conf_bus[27] ),
    .S(psn_net_3),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _06001_ (.A0(\cb_north.inst.cb_conf_bus[27] ),
    .A1(\cb_north.inst.cb_conf_bus[28] ),
    .S(psn_net_3),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _06002_ (.A0(\cb_north.inst.cb_conf_bus[28] ),
    .A1(\cb_north.inst.cb_conf_bus[29] ),
    .S(psn_net_3),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _06003_ (.A0(\cb_north.inst.cb_conf_bus[29] ),
    .A1(\cb_north.inst.cb_conf_bus[30] ),
    .S(psn_net_3),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _06004_ (.A0(\cb_north.inst.cb_conf_bus[30] ),
    .A1(\cb_north.inst.cb_conf_bus[31] ),
    .S(psn_net_3),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _06005_ (.A0(\cb_north.inst.cb_conf_bus[31] ),
    .A1(\cb_north.inst.cb_conf_bus[32] ),
    .S(psn_net_3),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _06006_ (.A0(\cb_north.inst.cb_conf_bus[32] ),
    .A1(\cb_north.inst.cb_conf_bus[33] ),
    .S(psn_net_3),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _06007_ (.A0(\cb_north.inst.cb_conf_bus[33] ),
    .A1(\cb_north.inst.cb_conf_bus[34] ),
    .S(psn_net_3),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _06008_ (.A0(\cb_north.inst.cb_conf_bus[34] ),
    .A1(\cb_north.inst.cb_conf_bus[35] ),
    .S(psn_net_3),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _06009_ (.A0(\cb_north.inst.cb_conf_bus[35] ),
    .A1(\cb_north.inst.cb_conf_bus[36] ),
    .S(psn_net_3),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _06010_ (.A0(\cb_north.inst.cb_conf_bus[36] ),
    .A1(\cb_north.inst.cb_conf_bus[37] ),
    .S(psn_net_3),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _06011_ (.A0(\cb_north.inst.cb_conf_bus[37] ),
    .A1(\cb_north.inst.cb_conf_bus[38] ),
    .S(psn_net_3),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _06012_ (.A0(\cb_north.inst.cb_conf_bus[38] ),
    .A1(\cb_north.inst.cb_conf_bus[39] ),
    .S(psn_net_3),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _06013_ (.A0(\cb_north.inst.cb_conf_bus[39] ),
    .A1(\cb_north.inst.cb_conf_bus[40] ),
    .S(psn_net_3),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _06014_ (.A0(\cb_north.inst.cb_conf_bus[40] ),
    .A1(\cb_north.inst.cb_conf_bus[41] ),
    .S(psn_net_3),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _06015_ (.A0(\cb_north.inst.cb_conf_bus[41] ),
    .A1(\cb_north.inst.cb_conf_bus[42] ),
    .S(psn_net_8),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _06016_ (.A0(\cb_north.inst.cb_conf_bus[42] ),
    .A1(\cb_north.inst.cb_conf_bus[43] ),
    .S(psn_net_8),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _06017_ (.A0(\cb_north.inst.cb_conf_bus[43] ),
    .A1(\cb_north.inst.cb_conf_bus[44] ),
    .S(psn_net_8),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _06018_ (.A0(\cb_north.inst.cb_conf_bus[44] ),
    .A1(\cb_north.inst.cb_conf_bus[45] ),
    .S(psn_net_8),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _06019_ (.A0(\cb_north.inst.cb_conf_bus[45] ),
    .A1(\cb_north.inst.cb_conf_bus[46] ),
    .S(psn_net_8),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _06020_ (.A0(\cb_north.inst.cb_conf_bus[46] ),
    .A1(\cb_north.inst.cb_conf_bus[47] ),
    .S(psn_net_8),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _06021_ (.A0(\cb_north.inst.cb_conf_bus[47] ),
    .A1(\cb_north.inst.cb_conf_bus[48] ),
    .S(psn_net_8),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _06022_ (.A0(\cb_north.inst.cb_conf_bus[48] ),
    .A1(\cb_north.inst.cb_conf_bus[49] ),
    .S(psn_net_8),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _06023_ (.A0(\cb_north.inst.cb_conf_bus[49] ),
    .A1(\cb_north.inst.cb_conf_bus[50] ),
    .S(psn_net_8),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _06024_ (.A0(\cb_north.inst.cb_conf_bus[50] ),
    .A1(\cb_north.inst.cb_conf_bus[51] ),
    .S(psn_net_8),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_1 _06025_ (.A0(\cb_north.inst.cb_conf_bus[51] ),
    .A1(\cb_north.inst.cb_conf_bus[52] ),
    .S(psn_net_9),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _06026_ (.A0(\cb_north.inst.cb_conf_bus[52] ),
    .A1(\cb_north.inst.cb_conf_bus[53] ),
    .S(psn_net_9),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _06027_ (.A0(\cb_north.inst.cb_conf_bus[53] ),
    .A1(\cb_north.inst.cb_conf_bus[54] ),
    .S(psn_net_9),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_1 _06028_ (.A0(\cb_north.inst.cb_conf_bus[54] ),
    .A1(\cb_north.inst.cb_conf_bus[55] ),
    .S(psn_net_9),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _06029_ (.A0(\cb_north.inst.cb_conf_bus[55] ),
    .A1(\cb_north.inst.cb_conf_bus[56] ),
    .S(psn_net_9),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_1 _06030_ (.A0(\cb_north.inst.cb_conf_bus[56] ),
    .A1(\cb_north.inst.cb_conf_bus[57] ),
    .S(psn_net_9),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_1 _06031_ (.A0(\cb_north.inst.cb_conf_bus[57] ),
    .A1(\cb_north.inst.cb_conf_bus[58] ),
    .S(psn_net_9),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _06032_ (.A0(\cb_north.inst.cb_conf_bus[58] ),
    .A1(\cb_north.inst.cb_conf_bus[59] ),
    .S(psn_net_9),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_1 _06033_ (.A0(\cb_north.inst.cb_conf_bus[59] ),
    .A1(\cb_north.inst.cb_conf_bus[60] ),
    .S(psn_net_9),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_1 _06034_ (.A0(\cb_north.inst.cb_conf_bus[60] ),
    .A1(\cb_north.inst.cb_conf_bus[61] ),
    .S(psn_net_9),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _06035_ (.A0(\cb_north.inst.cb_conf_bus[61] ),
    .A1(\cb_north.inst.cb_conf_bus[62] ),
    .S(psn_net_9),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _06036_ (.A0(\cb_north.inst.cb_conf_bus[62] ),
    .A1(\cb_north.inst.cb_conf_bus[63] ),
    .S(psn_net_9),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _06037_ (.A0(\cb_north.inst.cb_conf_bus[63] ),
    .A1(\cb_north.inst.cb_conf_bus[64] ),
    .S(psn_net_9),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _06038_ (.A0(\cb_north.inst.cb_conf_bus[64] ),
    .A1(\cb_north.inst.cb_conf_bus[65] ),
    .S(psn_net_9),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _06039_ (.A0(\cb_north.inst.cb_conf_bus[65] ),
    .A1(\cb_north.inst.cb_conf_bus[66] ),
    .S(psn_net_9),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _06040_ (.A0(\cb_north.inst.cb_conf_bus[66] ),
    .A1(\cb_north.inst.cb_conf_bus[67] ),
    .S(psn_net_9),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_1 _06041_ (.A0(\cb_north.inst.cb_conf_bus[67] ),
    .A1(\cb_north.inst.cb_conf_bus[68] ),
    .S(psn_net_9),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_1 _06042_ (.A0(\cb_north.inst.cb_conf_bus[68] ),
    .A1(\cb_north.inst.cb_conf_bus[69] ),
    .S(psn_net_9),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _06043_ (.A0(\cb_north.inst.cb_conf_bus[69] ),
    .A1(\cb_north.inst.cb_conf_bus[70] ),
    .S(psn_net_9),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _06044_ (.A0(\cb_north.inst.cb_conf_bus[70] ),
    .A1(\cb_north.inst.cb_conf_bus[71] ),
    .S(psn_net_9),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _06045_ (.A0(\cb_north.inst.cb_conf_bus[71] ),
    .A1(\cb_north.inst.cb_conf_bus[72] ),
    .S(psn_net_9),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _06046_ (.A0(\cb_north.inst.cb_conf_bus[72] ),
    .A1(\cb_north.inst.cb_conf_bus[73] ),
    .S(psn_net_9),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _06047_ (.A0(\cb_north.inst.cb_conf_bus[73] ),
    .A1(\cb_north.inst.cb_conf_bus[74] ),
    .S(psn_net_9),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _06048_ (.A0(\cb_north.inst.cb_conf_bus[74] ),
    .A1(\cb_north.inst.cb_conf_bus[75] ),
    .S(psn_net_9),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _06049_ (.A0(\cb_north.inst.cb_conf_bus[75] ),
    .A1(\cb_north.inst.cb_conf_bus[76] ),
    .S(psn_net_9),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _06050_ (.A0(\cb_north.inst.cb_conf_bus[76] ),
    .A1(\cb_north.inst.cb_conf_bus[77] ),
    .S(psn_net_3),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _06051_ (.A0(\cb_north.inst.cb_conf_bus[77] ),
    .A1(\cb_north.inst.cb_conf_bus[78] ),
    .S(psn_net_3),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _06052_ (.A0(\cb_north.inst.cb_conf_bus[78] ),
    .A1(\cb_north.inst.cb_conf_bus[79] ),
    .S(psn_net_3),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_1 _06053_ (.A0(\cb_north.inst.cb_conf_bus[79] ),
    .A1(\cb_north.inst.cb_conf_bus[80] ),
    .S(psn_net_3),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_1 _06054_ (.A0(\cb_north.inst.cb_conf_bus[80] ),
    .A1(\cb_north.inst.cb_conf_bus[81] ),
    .S(psn_net_3),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _06055_ (.A0(\cb_north.inst.cb_conf_bus[81] ),
    .A1(\cb_north.inst.cb_conf_bus[82] ),
    .S(psn_net_3),
    .X(_03440_));
 sky130_fd_sc_hd__mux2_1 _06056_ (.A0(\cb_north.inst.cb_conf_bus[82] ),
    .A1(\cb_north.inst.cb_conf_bus[83] ),
    .S(psn_net_3),
    .X(_03442_));
 sky130_fd_sc_hd__mux2_1 _06057_ (.A0(\cb_north.inst.cb_conf_bus[83] ),
    .A1(\cb_north.inst.cb_conf_bus[84] ),
    .S(psn_net_3),
    .X(_03444_));
 sky130_fd_sc_hd__mux2_1 _06058_ (.A0(\cb_north.inst.cb_conf_bus[84] ),
    .A1(\cb_north.inst.cb_conf_bus[85] ),
    .S(psn_net_3),
    .X(_03446_));
 sky130_fd_sc_hd__mux2_1 _06059_ (.A0(\cb_north.inst.cb_conf_bus[85] ),
    .A1(\cb_north.inst.cb_conf_bus[86] ),
    .S(psn_net_3),
    .X(_03448_));
 sky130_fd_sc_hd__mux2_1 _06060_ (.A0(\cb_north.inst.cb_conf_bus[86] ),
    .A1(\cb_north.inst.cb_conf_bus[87] ),
    .S(psn_net_3),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_1 _06061_ (.A0(\cb_north.inst.cb_conf_bus[87] ),
    .A1(\cb_north.inst.cb_conf_bus[88] ),
    .S(psn_net_3),
    .X(_03452_));
 sky130_fd_sc_hd__mux2_1 _06062_ (.A0(\cb_north.inst.cb_conf_bus[88] ),
    .A1(\cb_north.inst.cb_conf_bus[89] ),
    .S(psn_net_3),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_1 _06063_ (.A0(\cb_north.inst.cb_conf_bus[89] ),
    .A1(\cb_north.inst.cb_conf_bus[90] ),
    .S(psn_net_3),
    .X(_03456_));
 sky130_fd_sc_hd__mux2_1 _06064_ (.A0(\cb_north.inst.cb_conf_bus[90] ),
    .A1(\cb_north.inst.cb_conf_bus[91] ),
    .S(psn_net_3),
    .X(_03458_));
 sky130_fd_sc_hd__mux2_1 _06065_ (.A0(\cb_north.inst.cb_conf_bus[91] ),
    .A1(\cb_north.inst.cb_conf_bus[92] ),
    .S(psn_net_3),
    .X(_03460_));
 sky130_fd_sc_hd__mux2_1 _06066_ (.A0(\cb_north.inst.cb_conf_bus[92] ),
    .A1(\cb_north.inst.cb_conf_bus[93] ),
    .S(psn_net_9),
    .X(_03462_));
 sky130_fd_sc_hd__mux2_1 _06067_ (.A0(\cb_north.inst.cb_conf_bus[93] ),
    .A1(\cb_north.inst.cb_conf_bus[94] ),
    .S(psn_net_9),
    .X(_03464_));
 sky130_fd_sc_hd__mux2_1 _06068_ (.A0(\cb_north.inst.cb_conf_bus[94] ),
    .A1(\cb_north.inst.cb_conf_bus[95] ),
    .S(psn_net_9),
    .X(_03466_));
 sky130_fd_sc_hd__mux2_1 _06069_ (.A0(\cb_north.inst.cb_conf_bus[95] ),
    .A1(\cb_north.inst.cb_conf_bus[96] ),
    .S(psn_net_9),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _06070_ (.A0(\cb_north.inst.cb_conf_bus[96] ),
    .A1(\cb_north.inst.cb_conf_bus[97] ),
    .S(psn_net_9),
    .X(_03470_));
 sky130_fd_sc_hd__mux2_1 _06071_ (.A0(\cb_north.inst.cb_conf_bus[97] ),
    .A1(\cb_north.inst.cb_conf_bus[98] ),
    .S(psn_net_9),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _06072_ (.A0(\cb_north.inst.cb_conf_bus[98] ),
    .A1(\cb_north.inst.cb_conf_bus[99] ),
    .S(psn_net_9),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _06073_ (.A0(\cb_north.inst.cb_conf_bus[99] ),
    .A1(\cb_north.inst.cb_conf_bus[100] ),
    .S(psn_net_9),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_1 _06074_ (.A0(\cb_north.inst.cb_conf_bus[100] ),
    .A1(\cb_north.inst.cb_conf_bus[101] ),
    .S(psn_net_9),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _06075_ (.A0(\cb_north.inst.cb_conf_bus[101] ),
    .A1(\cb_north.inst.cb_conf_bus[102] ),
    .S(psn_net_9),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _06076_ (.A0(\cb_north.inst.cb_conf_bus[102] ),
    .A1(\cb_north.inst.cb_conf_bus[103] ),
    .S(psn_net_9),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_1 _06077_ (.A0(\cb_north.inst.cb_conf_bus[103] ),
    .A1(\cb_north.inst.cb_conf_bus[104] ),
    .S(psn_net_9),
    .X(_03484_));
 sky130_fd_sc_hd__mux2_1 _06078_ (.A0(\cb_north.inst.cb_conf_bus[104] ),
    .A1(\cb_north.inst.cb_conf_bus[105] ),
    .S(psn_net_9),
    .X(_03486_));
 sky130_fd_sc_hd__mux2_1 _06079_ (.A0(\cb_north.inst.cb_conf_bus[105] ),
    .A1(\cb_north.inst.cb_conf_bus[106] ),
    .S(psn_net_9),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_1 _06080_ (.A0(\cb_north.inst.cb_conf_bus[106] ),
    .A1(\cb_north.inst.cb_conf_bus[107] ),
    .S(psn_net_9),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _06081_ (.A0(\cb_north.inst.cb_conf_bus[107] ),
    .A1(\cb_north.inst.cb_conf_bus[108] ),
    .S(psn_net_9),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_1 _06082_ (.A0(\cb_north.inst.cb_conf_bus[108] ),
    .A1(\cb_north.inst.cb_conf_bus[109] ),
    .S(psn_net_9),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_1 _06083_ (.A0(\cb_north.inst.cb_conf_bus[109] ),
    .A1(\cb_north.inst.cb_conf_bus[110] ),
    .S(psn_net_9),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_1 _06084_ (.A0(\cb_north.inst.cb_conf_bus[110] ),
    .A1(\cb_north.inst.cb_conf_bus[111] ),
    .S(psn_net_9),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _06085_ (.A0(\cb_north.inst.cb_conf_bus[111] ),
    .A1(\cb_north.inst.cb_conf_bus[112] ),
    .S(psn_net_9),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_1 _06086_ (.A0(\cb_north.inst.cb_conf_bus[112] ),
    .A1(\cb_north.inst.cb_conf_bus[113] ),
    .S(psn_net_9),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_1 _06087_ (.A0(\cb_north.inst.cb_conf_bus[113] ),
    .A1(\cb_north.inst.cb_conf_bus[114] ),
    .S(psn_net_8),
    .X(_03504_));
 sky130_fd_sc_hd__mux2_1 _06088_ (.A0(\cb_north.inst.cb_conf_bus[114] ),
    .A1(\cb_north.inst.cb_conf_bus[115] ),
    .S(psn_net_8),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_1 _06089_ (.A0(\cb_north.inst.cb_conf_bus[115] ),
    .A1(\cb_north.inst.cb_conf_bus[116] ),
    .S(psn_net_8),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _06090_ (.A0(\cb_north.inst.cb_conf_bus[116] ),
    .A1(\cb_north.inst.cb_conf_bus[117] ),
    .S(psn_net_8),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _06091_ (.A0(\cb_north.inst.cb_conf_bus[117] ),
    .A1(\cb_north.inst.cb_conf_bus[118] ),
    .S(psn_net_8),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _06092_ (.A0(\cb_north.inst.cb_conf_bus[118] ),
    .A1(\cb_north.inst.cb_conf_bus[119] ),
    .S(psn_net_8),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _06093_ (.A0(\cb_north.inst.cb_conf_bus[119] ),
    .A1(\cb_north.inst.cb_conf_bus[120] ),
    .S(psn_net_8),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _06094_ (.A0(\cb_north.inst.cb_conf_bus[120] ),
    .A1(\cb_north.inst.cb_conf_bus[121] ),
    .S(psn_net_8),
    .X(_03518_));
 sky130_fd_sc_hd__mux2_1 _06095_ (.A0(\cb_north.inst.cb_conf_bus[121] ),
    .A1(\cb_north.inst.cb_conf_bus[122] ),
    .S(psn_net_8),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _06096_ (.A0(\cb_north.inst.cb_conf_bus[122] ),
    .A1(\cb_north.inst.cb_conf_bus[123] ),
    .S(psn_net_8),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_1 _06097_ (.A0(\cb_north.inst.cb_conf_bus[123] ),
    .A1(\cb_north.inst.cb_conf_bus[124] ),
    .S(psn_net_8),
    .X(_03524_));
 sky130_fd_sc_hd__mux2_1 _06098_ (.A0(\cb_north.inst.cb_conf_bus[124] ),
    .A1(\cb_north.inst.cb_conf_bus[125] ),
    .S(psn_net_8),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _06099_ (.A0(\cb_north.inst.cb_conf_bus[125] ),
    .A1(\cb_north.inst.cb_conf_bus[126] ),
    .S(psn_net_8),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _06100_ (.A0(\cb_north.inst.cb_conf_bus[126] ),
    .A1(\cb_north.inst.cb_conf_bus[127] ),
    .S(psn_net_8),
    .X(_03530_));
 sky130_fd_sc_hd__mux2_1 _06101_ (.A0(\cb_north.inst.cb_conf_bus[127] ),
    .A1(\cb_north.inst.cb_conf_bus[128] ),
    .S(psn_net_8),
    .X(_03532_));
 sky130_fd_sc_hd__mux2_1 _06102_ (.A0(\cb_north.inst.cb_conf_bus[128] ),
    .A1(\cb_north.inst.cb_conf_bus[129] ),
    .S(psn_net_8),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _06103_ (.A0(\cb_north.inst.cb_conf_bus[129] ),
    .A1(\cb_north.inst.cb_conf_bus[130] ),
    .S(psn_net_8),
    .X(_03536_));
 sky130_fd_sc_hd__mux2_1 _06104_ (.A0(\cb_north.inst.cb_conf_bus[130] ),
    .A1(\cb_north.inst.cb_conf_bus[131] ),
    .S(psn_net_8),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _06105_ (.A0(\cb_north.inst.cb_conf_bus[131] ),
    .A1(\cb_north.inst.cb_conf_bus[132] ),
    .S(psn_net_8),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _06106_ (.A0(\cb_north.inst.cb_conf_bus[132] ),
    .A1(\cb_north.inst.cb_conf_bus[133] ),
    .S(psn_net_8),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _06107_ (.A0(\cb_north.inst.cb_conf_bus[133] ),
    .A1(\cb_north.inst.cb_conf_bus[134] ),
    .S(psn_net_8),
    .X(_03544_));
 sky130_fd_sc_hd__mux2_1 _06108_ (.A0(\cb_north.inst.cb_conf_bus[134] ),
    .A1(\cb_north.inst.cb_conf_bus[135] ),
    .S(psn_net_8),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _06109_ (.A0(\cb_north.inst.cb_conf_bus[135] ),
    .A1(\cb_north.inst.cb_conf_bus[136] ),
    .S(psn_net_8),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_1 _06110_ (.A0(\cb_north.inst.cb_conf_bus[136] ),
    .A1(\cb_north.inst.cb_conf_bus[137] ),
    .S(psn_net_8),
    .X(_03550_));
 sky130_fd_sc_hd__mux2_1 _06111_ (.A0(\cb_north.inst.cb_conf_bus[137] ),
    .A1(\cb_north.inst.cb_conf_bus[138] ),
    .S(psn_net_8),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _06112_ (.A0(\cb_north.inst.cb_conf_bus[138] ),
    .A1(\cb_north.inst.cb_conf_bus[139] ),
    .S(psn_net_8),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_1 _06113_ (.A0(\cb_north.inst.cb_conf_bus[139] ),
    .A1(\cb_north.inst.cb_conf_bus[140] ),
    .S(psn_net_8),
    .X(_03556_));
 sky130_fd_sc_hd__mux2_1 _06114_ (.A0(\cb_north.inst.cb_conf_bus[140] ),
    .A1(\cb_north.inst.cb_conf_bus[141] ),
    .S(psn_net_4),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _06115_ (.A0(\cb_north.inst.cb_conf_bus[141] ),
    .A1(\cb_north.inst.cb_conf_bus[142] ),
    .S(psn_net_4),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _06116_ (.A0(\cb_north.inst.cb_conf_bus[142] ),
    .A1(\cb_north.inst.cb_conf_bus[143] ),
    .S(psn_net_4),
    .X(_03562_));
 sky130_fd_sc_hd__mux2_1 _06117_ (.A0(\cb_north.inst.cb_conf_bus[143] ),
    .A1(\cb_north.inst.cb_conf_bus[144] ),
    .S(psn_net_4),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _06118_ (.A0(\cb_north.inst.cb_conf_bus[144] ),
    .A1(\cb_north.inst.cb_conf_bus[145] ),
    .S(psn_net_4),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_1 _06119_ (.A0(\cb_north.inst.cb_conf_bus[145] ),
    .A1(\cb_north.inst.cb_conf_bus[146] ),
    .S(psn_net_4),
    .X(_03568_));
 sky130_fd_sc_hd__mux2_1 _06120_ (.A0(\cb_north.inst.cb_conf_bus[146] ),
    .A1(\cb_north.inst.cb_conf_bus[147] ),
    .S(psn_net_3),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_1 _06121_ (.A0(\cb_north.inst.cb_conf_bus[147] ),
    .A1(\cb_north.inst.cb_conf_bus[148] ),
    .S(psn_net_3),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _06122_ (.A0(\cb_north.inst.cb_conf_bus[148] ),
    .A1(\cb_north.inst.cb_conf_bus[149] ),
    .S(psn_net_3),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _06123_ (.A0(\cb_north.inst.cb_conf_bus[149] ),
    .A1(\cb_north.inst.cb_conf_bus[150] ),
    .S(psn_net_3),
    .X(_03576_));
 sky130_fd_sc_hd__mux2_1 _06124_ (.A0(\cb_north.inst.cb_conf_bus[150] ),
    .A1(\cb_north.inst.cb_conf_bus[151] ),
    .S(psn_net_3),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _06125_ (.A0(\cb_north.inst.cb_conf_bus[151] ),
    .A1(\cb_north.inst.cb_conf_bus[152] ),
    .S(psn_net_3),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _06126_ (.A0(\cb_north.inst.cb_conf_bus[152] ),
    .A1(\cb_north.inst.cb_conf_bus[153] ),
    .S(psn_net_3),
    .X(_03582_));
 sky130_fd_sc_hd__mux2_1 _06127_ (.A0(\cb_north.inst.cb_conf_bus[153] ),
    .A1(\cb_north.inst.cb_conf_bus[154] ),
    .S(psn_net_3),
    .X(_03584_));
 sky130_fd_sc_hd__mux2_1 _06128_ (.A0(\cb_north.inst.cb_conf_bus[154] ),
    .A1(\cb_north.inst.cb_conf_bus[155] ),
    .S(psn_net_3),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _06129_ (.A0(\cb_north.inst.cb_conf_bus[155] ),
    .A1(\cb_north.inst.cb_conf_bus[156] ),
    .S(psn_net_3),
    .X(_03588_));
 sky130_fd_sc_hd__mux2_1 _06130_ (.A0(\cb_north.inst.cb_conf_bus[156] ),
    .A1(\cb_north.inst.cb_conf_bus[157] ),
    .S(psn_net_3),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_1 _06131_ (.A0(\cb_north.inst.cb_conf_bus[157] ),
    .A1(\cb_north.inst.cb_conf_bus[158] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _06132_ (.A0(\cb_north.inst.cb_conf_bus[158] ),
    .A1(\cb_north.inst.cb_conf_bus[159] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03594_));
 sky130_fd_sc_hd__mux2_1 _06133_ (.A0(\cb_north.inst.cb_conf_bus[159] ),
    .A1(\cb_north.inst.cb_conf_bus[160] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _06134_ (.A0(\cb_north.inst.cb_conf_bus[160] ),
    .A1(\cb_north.inst.cb_conf_bus[161] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_1 _06135_ (.A0(\cb_north.inst.cb_conf_bus[161] ),
    .A1(\cb_north.inst.cb_conf_bus[162] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03600_));
 sky130_fd_sc_hd__mux2_1 _06136_ (.A0(\cb_north.inst.cb_conf_bus[162] ),
    .A1(\cb_north.inst.cb_conf_bus[163] ),
    .S(psn_net_5),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _06137_ (.A0(\cb_north.inst.cb_conf_bus[163] ),
    .A1(\cb_north.inst.cb_conf_bus[164] ),
    .S(psn_net_5),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _06138_ (.A0(\cb_north.inst.cb_conf_bus[164] ),
    .A1(\cb_north.inst.cb_conf_bus[165] ),
    .S(psn_net_5),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _06139_ (.A0(\cb_north.inst.cb_conf_bus[165] ),
    .A1(\cb_north.inst.cb_conf_bus[166] ),
    .S(psn_net_8),
    .X(_03608_));
 sky130_fd_sc_hd__mux2_1 _06140_ (.A0(\cb_north.inst.cb_conf_bus[166] ),
    .A1(\cb_north.inst.cb_conf_bus[167] ),
    .S(psn_net_8),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _06141_ (.A0(\cb_north.inst.cb_conf_bus[167] ),
    .A1(\cb_north.inst.cb_conf_bus[168] ),
    .S(psn_net_8),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _06142_ (.A0(\cb_north.inst.cb_conf_bus[168] ),
    .A1(\cb_north.inst.cb_conf_bus[169] ),
    .S(psn_net_8),
    .X(_03614_));
 sky130_fd_sc_hd__mux2_1 _06143_ (.A0(\cb_north.inst.cb_conf_bus[169] ),
    .A1(\cb_north.inst.cb_conf_bus[170] ),
    .S(psn_net_5),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _06144_ (.A0(\cb_north.inst.cb_conf_bus[170] ),
    .A1(\cb_north.inst.cb_conf_bus[171] ),
    .S(psn_net_5),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _06145_ (.A0(\cb_north.inst.cb_conf_bus[171] ),
    .A1(\cb_north.inst.cb_conf_bus[172] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03620_));
 sky130_fd_sc_hd__mux2_1 _06146_ (.A0(\cb_north.inst.cb_conf_bus[172] ),
    .A1(\cb_north.inst.cb_conf_bus[173] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _06147_ (.A0(\cb_north.inst.cb_conf_bus[173] ),
    .A1(\cb_north.inst.cb_conf_bus[174] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _06148_ (.A0(\cb_north.inst.cb_conf_bus[174] ),
    .A1(\cb_north.inst.cb_conf_bus[175] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03626_));
 sky130_fd_sc_hd__mux2_1 _06149_ (.A0(\cb_north.inst.cb_conf_bus[175] ),
    .A1(\cb_north.inst.cb_conf_bus[176] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _06150_ (.A0(\cb_north.inst.cb_conf_bus[176] ),
    .A1(\cb_north.inst.cb_conf_bus[177] ),
    .S(psn_net_18),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_1 _06151_ (.A0(\cb_north.inst.cb_conf_bus[177] ),
    .A1(\cb_north.inst.cb_conf_bus[178] ),
    .S(psn_net_18),
    .X(_03632_));
 sky130_fd_sc_hd__mux2_1 _06152_ (.A0(\cb_north.inst.cb_conf_bus[178] ),
    .A1(\cb_north.inst.cb_conf_bus[179] ),
    .S(psn_net_18),
    .X(_03634_));
 sky130_fd_sc_hd__mux2_1 _06153_ (.A0(\cb_north.inst.cb_conf_bus[179] ),
    .A1(\cb_north.inst.cb_conf_bus[180] ),
    .S(psn_net_11),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _06154_ (.A0(\cb_north.inst.cb_conf_bus[180] ),
    .A1(\cb_north.inst.cb_conf_bus[181] ),
    .S(psn_net_11),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _06155_ (.A0(\cb_north.inst.cb_conf_bus[181] ),
    .A1(\cb_north.inst.cb_conf_bus[182] ),
    .S(psn_net_11),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _06156_ (.A0(\cb_north.inst.cb_conf_bus[182] ),
    .A1(\cb_north.inst.cb_conf_bus[183] ),
    .S(psn_net_11),
    .X(_03642_));
 sky130_fd_sc_hd__mux2_1 _06157_ (.A0(\cb_north.inst.cb_conf_bus[183] ),
    .A1(\cb_north.inst.cb_conf_bus[184] ),
    .S(psn_net_11),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _06158_ (.A0(\cb_north.inst.cb_conf_bus[184] ),
    .A1(\cb_north.inst.cb_conf_bus[185] ),
    .S(psn_net_11),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _06159_ (.A0(\cb_north.inst.cb_conf_bus[185] ),
    .A1(\cb_north.inst.cb_conf_bus[186] ),
    .S(psn_net_11),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _06160_ (.A0(\cb_north.inst.cb_conf_bus[186] ),
    .A1(\cb_north.inst.cb_conf_bus[187] ),
    .S(psn_net_11),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _06161_ (.A0(\cb_north.inst.cb_conf_bus[187] ),
    .A1(\cb_north.inst.cb_conf_bus[188] ),
    .S(psn_net_11),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _06162_ (.A0(\cb_north.inst.cb_conf_bus[188] ),
    .A1(\cb_north.inst.cb_conf_bus[189] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _06163_ (.A0(\cb_north.inst.cb_conf_bus[189] ),
    .A1(\cb_north.inst.cb_conf_bus[190] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _06164_ (.A0(\cb_north.inst.cb_conf_bus[190] ),
    .A1(\cb_north.inst.cb_conf_bus[191] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _06165_ (.A0(\cb_north.inst.cb_conf_bus[191] ),
    .A1(\cb_north.inst.cb_conf_bus[192] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03660_));
 sky130_fd_sc_hd__mux2_1 _06166_ (.A0(\cb_north.inst.cb_conf_bus[192] ),
    .A1(\cb_north.inst.cb_conf_bus[193] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03662_));
 sky130_fd_sc_hd__mux2_1 _06167_ (.A0(\cb_north.inst.cb_conf_bus[193] ),
    .A1(\cb_north.inst.cb_conf_bus[194] ),
    .S(psn_net_7),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _06168_ (.A0(\cb_north.inst.cb_conf_bus[194] ),
    .A1(\cb_north.inst.cb_conf_bus[195] ),
    .S(psn_net_7),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _06169_ (.A0(\cb_north.inst.cb_conf_bus[195] ),
    .A1(\cb_north.inst.cb_conf_bus[196] ),
    .S(psn_net_7),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _06170_ (.A0(\cb_north.inst.cb_conf_bus[196] ),
    .A1(\cb_north.inst.cb_conf_bus[197] ),
    .S(psn_net_7),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_1 _06171_ (.A0(\cb_north.inst.cb_conf_bus[197] ),
    .A1(\cb_north.inst.cb_conf_bus[198] ),
    .S(psn_net_8),
    .X(_03672_));
 sky130_fd_sc_hd__mux2_1 _06172_ (.A0(\cb_north.inst.cb_conf_bus[198] ),
    .A1(\cb_north.inst.cb_conf_bus[199] ),
    .S(psn_net_8),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _06173_ (.A0(\cb_north.inst.cb_conf_bus[199] ),
    .A1(\cb_north.inst.cb_conf_bus[200] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _06174_ (.A0(\cb_north.inst.cb_conf_bus[200] ),
    .A1(\cb_north.inst.cb_conf_bus[201] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03678_));
 sky130_fd_sc_hd__mux2_1 _06175_ (.A0(\cb_north.inst.cb_conf_bus[201] ),
    .A1(\cb_north.inst.cb_conf_bus[202] ),
    .S(psn_net_10),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _06176_ (.A0(\cb_north.inst.cb_conf_bus[202] ),
    .A1(\cb_north.inst.cb_conf_bus[203] ),
    .S(psn_net_10),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _06177_ (.A0(\cb_north.inst.cb_conf_bus[203] ),
    .A1(\cb_north.inst.cb_conf_bus[204] ),
    .S(psn_net_10),
    .X(_03684_));
 sky130_fd_sc_hd__mux2_1 _06178_ (.A0(\cb_north.inst.cb_conf_bus[204] ),
    .A1(\cb_north.inst.cb_conf_bus[205] ),
    .S(psn_net_10),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _06179_ (.A0(\cb_north.inst.cb_conf_bus[205] ),
    .A1(\cb_north.inst.cb_conf_bus[206] ),
    .S(psn_net_10),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _06180_ (.A0(\cb_north.inst.cb_conf_bus[206] ),
    .A1(\cb_north.inst.cb_conf_bus[207] ),
    .S(psn_net_10),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _06181_ (.A0(\cb_north.inst.cb_conf_bus[207] ),
    .A1(\cb_north.inst.cb_conf_bus[208] ),
    .S(psn_net_10),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _06182_ (.A0(\cb_north.inst.cb_conf_bus[208] ),
    .A1(\cb_north.inst.cb_conf_bus[209] ),
    .S(psn_net_10),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _06183_ (.A0(\cb_north.inst.cb_conf_bus[209] ),
    .A1(\cb_north.inst.cb_conf_bus[210] ),
    .S(psn_net_10),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _06184_ (.A0(\cb_north.inst.cb_conf_bus[210] ),
    .A1(\cb_north.inst.cb_conf_bus[211] ),
    .S(psn_net_10),
    .X(_03698_));
 sky130_fd_sc_hd__mux2_1 _06185_ (.A0(\cb_north.inst.cb_conf_bus[211] ),
    .A1(\cb_north.inst.cb_conf_bus[212] ),
    .S(psn_net_10),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _06186_ (.A0(\cb_north.inst.cb_conf_bus[212] ),
    .A1(\cb_north.inst.cb_conf_bus[213] ),
    .S(psn_net_10),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _06187_ (.A0(\cb_north.inst.cb_conf_bus[213] ),
    .A1(\cb_north.inst.cb_conf_bus[214] ),
    .S(psn_net_10),
    .X(_03704_));
 sky130_fd_sc_hd__mux2_1 _06188_ (.A0(\cb_north.inst.cb_conf_bus[214] ),
    .A1(\cb_north.inst.cb_conf_bus[215] ),
    .S(psn_net_10),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _06189_ (.A0(\cb_north.inst.cb_conf_bus[215] ),
    .A1(\cb_north.inst.cb_conf_bus[216] ),
    .S(psn_net_10),
    .X(_03708_));
 sky130_fd_sc_hd__mux2_1 _06190_ (.A0(\cb_north.inst.cb_conf_bus[216] ),
    .A1(\cb_north.inst.cb_conf_bus[217] ),
    .S(psn_net_10),
    .X(_03710_));
 sky130_fd_sc_hd__mux2_1 _06191_ (.A0(\cb_north.inst.cb_conf_bus[217] ),
    .A1(\cb_north.inst.cb_conf_bus[218] ),
    .S(psn_net_10),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_1 _06192_ (.A0(\cb_north.inst.cb_conf_bus[218] ),
    .A1(\cb_north.inst.cb_conf_bus[219] ),
    .S(psn_net_10),
    .X(_03714_));
 sky130_fd_sc_hd__mux2_1 _06193_ (.A0(\cb_north.inst.cb_conf_bus[219] ),
    .A1(\cb_north.inst.cb_conf_bus[220] ),
    .S(psn_net_10),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_1 _06194_ (.A0(\cb_north.inst.cb_conf_bus[220] ),
    .A1(\cb_north.inst.cb_conf_bus[221] ),
    .S(psn_net_10),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_1 _06195_ (.A0(\cb_north.inst.cb_conf_bus[221] ),
    .A1(\cb_north.inst.cb_conf_bus[222] ),
    .S(psn_net_10),
    .X(_03720_));
 sky130_fd_sc_hd__mux2_1 _06196_ (.A0(\cb_north.inst.cb_conf_bus[222] ),
    .A1(\cb_north.inst.cb_conf_bus[223] ),
    .S(psn_net_10),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _06197_ (.A0(\cb_north.inst.cb_conf_bus[223] ),
    .A1(\cb_north.inst.cb_conf_bus[224] ),
    .S(psn_net_10),
    .X(_03724_));
 sky130_fd_sc_hd__mux2_1 _06198_ (.A0(\cb_north.inst.cb_conf_bus[224] ),
    .A1(\cb_north.inst.cb_conf_bus[225] ),
    .S(psn_net_10),
    .X(_03726_));
 sky130_fd_sc_hd__mux2_1 _06199_ (.A0(\cb_north.inst.cb_conf_bus[225] ),
    .A1(\cb_north.inst.cb_conf_bus[226] ),
    .S(psn_net_10),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _06200_ (.A0(\cb_north.inst.cb_conf_bus[226] ),
    .A1(\cb_north.inst.cb_conf_bus[227] ),
    .S(psn_net_10),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _06201_ (.A0(\cb_north.inst.cb_conf_bus[227] ),
    .A1(\cb_north.inst.cb_conf_bus[228] ),
    .S(psn_net_10),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _06202_ (.A0(\cb_north.inst.cb_conf_bus[228] ),
    .A1(\cb_north.inst.cb_conf_bus[229] ),
    .S(psn_net_10),
    .X(_03734_));
 sky130_fd_sc_hd__mux2_1 _06203_ (.A0(\cb_north.inst.cb_conf_bus[229] ),
    .A1(\cb_north.inst.cb_conf_bus[230] ),
    .S(psn_net_10),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _06204_ (.A0(\cb_north.inst.cb_conf_bus[230] ),
    .A1(\cb_north.inst.cb_conf_bus[231] ),
    .S(psn_net_10),
    .X(_03738_));
 sky130_fd_sc_hd__mux2_1 _06205_ (.A0(\cb_north.inst.cb_conf_bus[231] ),
    .A1(\cb_north.inst.cb_conf_bus[232] ),
    .S(psn_net_10),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _06206_ (.A0(\cb_north.inst.cb_conf_bus[232] ),
    .A1(\cb_north.inst.cb_conf_bus[233] ),
    .S(psn_net_10),
    .X(_03742_));
 sky130_fd_sc_hd__mux2_1 _06207_ (.A0(\cb_north.inst.cb_conf_bus[233] ),
    .A1(\cb_north.inst.cb_conf_bus[234] ),
    .S(psn_net_10),
    .X(_03744_));
 sky130_fd_sc_hd__mux2_1 _06208_ (.A0(\cb_north.inst.cb_conf_bus[234] ),
    .A1(\cb_north.inst.cb_conf_bus[235] ),
    .S(psn_net_10),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _06209_ (.A0(\cb_north.inst.cb_conf_bus[235] ),
    .A1(\cb_north.inst.cb_conf_bus[236] ),
    .S(psn_net_10),
    .X(_03748_));
 sky130_fd_sc_hd__mux2_1 _06210_ (.A0(\cb_north.inst.cb_conf_bus[236] ),
    .A1(\cb_north.inst.cb_conf_bus[237] ),
    .S(psn_net_10),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_1 _06211_ (.A0(\cb_north.inst.cb_conf_bus[237] ),
    .A1(\cb_north.inst.cb_conf_bus[238] ),
    .S(psn_net_10),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_1 _06212_ (.A0(\cb_north.inst.cb_conf_bus[238] ),
    .A1(\cb_north.inst.cb_conf_bus[239] ),
    .S(psn_net_10),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _06213_ (.A0(\cb_north.inst.cb_conf_bus[239] ),
    .A1(\cb_north.inst.cb_conf_bus[240] ),
    .S(psn_net_10),
    .X(_03756_));
 sky130_fd_sc_hd__mux2_1 _06214_ (.A0(\cb_north.inst.cb_conf_bus[240] ),
    .A1(\cb_north.inst.cb_conf_bus[241] ),
    .S(psn_net_10),
    .X(_03758_));
 sky130_fd_sc_hd__mux2_1 _06215_ (.A0(\cb_north.inst.cb_conf_bus[241] ),
    .A1(\cb_north.inst.cb_conf_bus[242] ),
    .S(psn_net_10),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _06216_ (.A0(\cb_north.inst.cb_conf_bus[242] ),
    .A1(\cb_north.inst.cb_conf_bus[243] ),
    .S(psn_net_10),
    .X(_03762_));
 sky130_fd_sc_hd__mux2_1 _06217_ (.A0(\cb_north.inst.cb_conf_bus[243] ),
    .A1(\cb_north.inst.cb_conf_bus[244] ),
    .S(psn_net_10),
    .X(_03764_));
 sky130_fd_sc_hd__mux2_1 _06218_ (.A0(\cb_north.inst.cb_conf_bus[244] ),
    .A1(\cb_north.inst.cb_conf_bus[245] ),
    .S(psn_net_10),
    .X(_03766_));
 sky130_fd_sc_hd__mux2_1 _06219_ (.A0(\cb_north.inst.cb_conf_bus[245] ),
    .A1(\cb_north.inst.cb_conf_bus[246] ),
    .S(psn_net_10),
    .X(_03768_));
 sky130_fd_sc_hd__mux2_1 _06220_ (.A0(\cb_north.inst.cb_conf_bus[246] ),
    .A1(\cb_north.inst.cb_conf_bus[247] ),
    .S(psn_net_10),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_1 _06221_ (.A0(\cb_north.inst.cb_conf_bus[247] ),
    .A1(\cb_north.inst.cb_conf_bus[248] ),
    .S(psn_net_10),
    .X(_03772_));
 sky130_fd_sc_hd__mux2_1 _06222_ (.A0(\cb_north.inst.cb_conf_bus[248] ),
    .A1(\cb_north.inst.cb_conf_bus[249] ),
    .S(psn_net_10),
    .X(_03774_));
 sky130_fd_sc_hd__mux2_1 _06223_ (.A0(\cb_north.inst.cb_conf_bus[249] ),
    .A1(\cb_north.inst.cb_conf_bus[250] ),
    .S(psn_net_10),
    .X(_03776_));
 sky130_fd_sc_hd__mux2_1 _06224_ (.A0(\cb_north.inst.cb_conf_bus[250] ),
    .A1(\cb_north.inst.cb_conf_bus[251] ),
    .S(psn_net_10),
    .X(_03778_));
 sky130_fd_sc_hd__mux2_1 _06225_ (.A0(\cb_north.inst.cb_conf_bus[251] ),
    .A1(\cb_north.inst.cb_conf_bus[252] ),
    .S(psn_net_10),
    .X(_03780_));
 sky130_fd_sc_hd__mux2_1 _06226_ (.A0(\cb_north.inst.cb_conf_bus[252] ),
    .A1(\cb_north.inst.cb_conf_bus[253] ),
    .S(psn_net_10),
    .X(_03782_));
 sky130_fd_sc_hd__mux2_1 _06227_ (.A0(\cb_north.inst.cb_conf_bus[253] ),
    .A1(\cb_north.inst.cb_conf_bus[254] ),
    .S(psn_net_10),
    .X(_03784_));
 sky130_fd_sc_hd__mux2_1 _06228_ (.A0(\cb_north.inst.cb_conf_bus[254] ),
    .A1(\cb_north.inst.cb_conf_bus[255] ),
    .S(psn_net_10),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_1 _06229_ (.A0(\cb_north.inst.cb_conf_bus[255] ),
    .A1(\cb_north.inst.cb_conf_bus[256] ),
    .S(psn_net_10),
    .X(_03788_));
 sky130_fd_sc_hd__mux2_1 _06230_ (.A0(\cb_north.inst.cb_conf_bus[256] ),
    .A1(\cb_north.inst.cb_conf_bus[257] ),
    .S(psn_net_10),
    .X(_03790_));
 sky130_fd_sc_hd__mux2_1 _06231_ (.A0(\cb_north.inst.cb_conf_bus[257] ),
    .A1(\cb_north.inst.cb_conf_bus[258] ),
    .S(psn_net_10),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_1 _06232_ (.A0(\cb_north.inst.cb_conf_bus[258] ),
    .A1(\cb_north.inst.cb_conf_bus[259] ),
    .S(psn_net_10),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_1 _06233_ (.A0(\cb_north.inst.cb_conf_bus[259] ),
    .A1(\cb_north.inst.cb_conf_bus[260] ),
    .S(psn_net_10),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_1 _06234_ (.A0(\cb_north.inst.cb_conf_bus[260] ),
    .A1(\cb_north.inst.cb_conf_bus[261] ),
    .S(psn_net_10),
    .X(_03798_));
 sky130_fd_sc_hd__mux2_1 _06235_ (.A0(\cb_north.inst.cb_conf_bus[261] ),
    .A1(\cb_north.inst.cb_conf_bus[262] ),
    .S(psn_net_10),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_1 _06236_ (.A0(\cb_north.inst.cb_conf_bus[262] ),
    .A1(\cb_north.inst.cb_conf_bus[263] ),
    .S(psn_net_10),
    .X(_03802_));
 sky130_fd_sc_hd__mux2_1 _06237_ (.A0(\cb_north.inst.cb_conf_bus[263] ),
    .A1(\cb_north.inst.cb_conf_bus[264] ),
    .S(psn_net_10),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _06238_ (.A0(\cb_north.inst.cb_conf_bus[264] ),
    .A1(\cb_north.inst.cb_conf_bus[265] ),
    .S(psn_net_10),
    .X(_03806_));
 sky130_fd_sc_hd__mux2_1 _06239_ (.A0(\cb_north.inst.cb_conf_bus[265] ),
    .A1(\cb_north.inst.cb_conf_bus[266] ),
    .S(psn_net_10),
    .X(_03808_));
 sky130_fd_sc_hd__mux2_1 _06240_ (.A0(\cb_north.inst.cb_conf_bus[266] ),
    .A1(\cb_north.inst.cb_conf_bus[267] ),
    .S(psn_net_10),
    .X(_03810_));
 sky130_fd_sc_hd__mux2_1 _06241_ (.A0(\cb_north.inst.cb_conf_bus[267] ),
    .A1(\cb_north.inst.cb_conf_bus[268] ),
    .S(psn_net_10),
    .X(_03812_));
 sky130_fd_sc_hd__mux2_1 _06242_ (.A0(\cb_north.inst.cb_conf_bus[268] ),
    .A1(\cb_north.inst.cb_conf_bus[269] ),
    .S(psn_net_10),
    .X(_03814_));
 sky130_fd_sc_hd__mux2_1 _06243_ (.A0(\cb_north.inst.cb_conf_bus[269] ),
    .A1(\cb_north.inst.cb_conf_bus[270] ),
    .S(psn_net_10),
    .X(_03816_));
 sky130_fd_sc_hd__mux2_1 _06244_ (.A0(\cb_north.inst.cb_conf_bus[270] ),
    .A1(\cb_north.inst.cb_conf_bus[271] ),
    .S(psn_net_10),
    .X(_03818_));
 sky130_fd_sc_hd__mux2_1 _06245_ (.A0(\cb_north.inst.cb_conf_bus[271] ),
    .A1(\cb_north.inst.cb_conf_bus[272] ),
    .S(psn_net_10),
    .X(_03820_));
 sky130_fd_sc_hd__mux2_1 _06246_ (.A0(\cb_north.inst.cb_conf_bus[272] ),
    .A1(\cb_north.inst.cb_conf_bus[273] ),
    .S(psn_net_10),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_1 _06247_ (.A0(\cb_north.inst.cb_conf_bus[273] ),
    .A1(\cb_north.inst.cb_conf_bus[274] ),
    .S(psn_net_10),
    .X(_03824_));
 sky130_fd_sc_hd__mux2_1 _06248_ (.A0(\cb_north.inst.cb_conf_bus[274] ),
    .A1(\cb_north.inst.cb_conf_bus[275] ),
    .S(psn_net_10),
    .X(_03826_));
 sky130_fd_sc_hd__mux2_1 _06249_ (.A0(\cb_north.inst.cb_conf_bus[275] ),
    .A1(\cb_north.inst.cb_conf_bus[276] ),
    .S(psn_net_10),
    .X(_03828_));
 sky130_fd_sc_hd__mux2_1 _06250_ (.A0(\cb_north.inst.cb_conf_bus[276] ),
    .A1(\cb_north.inst.cb_conf_bus[277] ),
    .S(psn_net_10),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _06251_ (.A0(\cb_north.inst.cb_conf_bus[277] ),
    .A1(\cb_north.inst.cb_conf_bus[278] ),
    .S(psn_net_10),
    .X(_03832_));
 sky130_fd_sc_hd__mux2_1 _06252_ (.A0(\cb_north.inst.cb_conf_bus[278] ),
    .A1(\cb_north.inst.cb_conf_bus[279] ),
    .S(psn_net_10),
    .X(_03834_));
 sky130_fd_sc_hd__mux2_1 _06253_ (.A0(\cb_north.inst.cb_conf_bus[279] ),
    .A1(\cb_north.inst.cb_conf_bus[280] ),
    .S(psn_net_10),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _06254_ (.A0(\cb_north.inst.cb_conf_bus[280] ),
    .A1(\cb_north.inst.cb_conf_bus[281] ),
    .S(psn_net_10),
    .X(_03838_));
 sky130_fd_sc_hd__mux2_1 _06255_ (.A0(\cb_north.inst.cb_conf_bus[281] ),
    .A1(\cb_north.inst.cb_conf_bus[282] ),
    .S(psn_net_10),
    .X(_03840_));
 sky130_fd_sc_hd__mux2_1 _06256_ (.A0(\cb_north.inst.cb_conf_bus[282] ),
    .A1(\cb_north.inst.cb_conf_bus[283] ),
    .S(psn_net_10),
    .X(_03842_));
 sky130_fd_sc_hd__mux2_1 _06257_ (.A0(\cb_north.inst.cb_conf_bus[283] ),
    .A1(\cb_north.inst.cb_conf_bus[284] ),
    .S(psn_net_10),
    .X(_03844_));
 sky130_fd_sc_hd__mux2_1 _06258_ (.A0(\cb_north.inst.cb_conf_bus[284] ),
    .A1(\cb_north.inst.cb_conf_bus[285] ),
    .S(psn_net_10),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_1 _06259_ (.A0(\cb_north.inst.cb_conf_bus[285] ),
    .A1(\cb_north.inst.cb_conf_bus[286] ),
    .S(psn_net_10),
    .X(_03848_));
 sky130_fd_sc_hd__mux2_1 _06260_ (.A0(\cb_north.inst.cb_conf_bus[286] ),
    .A1(\cb_north.inst.cb_conf_bus[287] ),
    .S(psn_net_10),
    .X(_03850_));
 sky130_fd_sc_hd__mux2_1 _06261_ (.A0(\cb_north.inst.cb_conf_bus[287] ),
    .A1(\cb_north.inst.cb_conf_bus[288] ),
    .S(psn_net_10),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_1 _06262_ (.A0(\cb_north.inst.cb_conf_bus[288] ),
    .A1(\cb_north.inst.cb_conf_bus[289] ),
    .S(psn_net_10),
    .X(_03854_));
 sky130_fd_sc_hd__mux2_1 _06263_ (.A0(\cb_north.inst.cb_conf_bus[289] ),
    .A1(\cb_north.inst.cb_conf_bus[290] ),
    .S(psn_net_10),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _06264_ (.A0(\cb_north.inst.cb_conf_bus[290] ),
    .A1(\cb_north.inst.cb_conf_bus[291] ),
    .S(psn_net_10),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_1 _06265_ (.A0(\cb_north.inst.cb_conf_bus[291] ),
    .A1(\cb_north.inst.cb_conf_bus[292] ),
    .S(psn_net_10),
    .X(_03860_));
 sky130_fd_sc_hd__mux2_1 _06266_ (.A0(\cb_north.inst.cb_conf_bus[292] ),
    .A1(\cb_north.inst.cb_conf_bus[293] ),
    .S(psn_net_10),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_1 _06267_ (.A0(\cb_north.inst.cb_conf_bus[293] ),
    .A1(\cb_north.inst.cb_conf_bus[294] ),
    .S(psn_net_16),
    .X(_03864_));
 sky130_fd_sc_hd__mux2_1 _06268_ (.A0(\cb_north.inst.cb_conf_bus[294] ),
    .A1(\cb_north.inst.cb_conf_bus[295] ),
    .S(psn_net_16),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_1 _06269_ (.A0(\cb_north.inst.cb_conf_bus[295] ),
    .A1(\cb_north.inst.cb_conf_bus[296] ),
    .S(psn_net_16),
    .X(_03868_));
 sky130_fd_sc_hd__mux2_1 _06270_ (.A0(\cb_north.inst.cb_conf_bus[296] ),
    .A1(\cb_north.inst.cb_conf_bus[297] ),
    .S(psn_net_16),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _06271_ (.A0(\cb_north.inst.cb_conf_bus[297] ),
    .A1(\cb_north.inst.cb_conf_bus[298] ),
    .S(psn_net_16),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _06272_ (.A0(\cb_north.inst.cb_conf_bus[298] ),
    .A1(\cb_north.inst.cb_conf_bus[299] ),
    .S(psn_net_16),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _06273_ (.A0(\cb_north.inst.cb_conf_bus[299] ),
    .A1(\cb_north.inst.cb_conf_bus[300] ),
    .S(psn_net_16),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _06274_ (.A0(\cb_north.inst.cb_conf_bus[300] ),
    .A1(\cb_north.inst.cb_conf_bus[301] ),
    .S(psn_net_16),
    .X(_03878_));
 sky130_fd_sc_hd__mux2_1 _06275_ (.A0(\cb_north.inst.cb_conf_bus[301] ),
    .A1(\cb_north.inst.cb_conf_bus[302] ),
    .S(psn_net_16),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _06276_ (.A0(\cb_north.inst.cb_conf_bus[302] ),
    .A1(\cb_north.inst.cb_conf_bus[303] ),
    .S(psn_net_16),
    .X(_03882_));
 sky130_fd_sc_hd__mux2_1 _06277_ (.A0(\cb_north.inst.cb_conf_bus[303] ),
    .A1(\cb_north.inst.cb_conf_bus[304] ),
    .S(psn_net_16),
    .X(_03884_));
 sky130_fd_sc_hd__mux2_1 _06278_ (.A0(\cb_north.inst.cb_conf_bus[304] ),
    .A1(\cb_north.inst.cb_conf_bus[305] ),
    .S(psn_net_16),
    .X(_03886_));
 sky130_fd_sc_hd__mux2_1 _06279_ (.A0(\cb_north.inst.cb_conf_bus[305] ),
    .A1(\cb_north.inst.cb_conf_bus[306] ),
    .S(psn_net_16),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _06280_ (.A0(\cb_north.inst.cb_conf_bus[306] ),
    .A1(\cb_north.inst.cb_conf_bus[307] ),
    .S(psn_net_16),
    .X(_03890_));
 sky130_fd_sc_hd__mux2_1 _06281_ (.A0(\cb_north.inst.cb_conf_bus[307] ),
    .A1(\cb_north.inst.cb_conf_bus[308] ),
    .S(psn_net_16),
    .X(_03892_));
 sky130_fd_sc_hd__mux2_1 _06282_ (.A0(\cb_north.inst.cb_conf_bus[308] ),
    .A1(\cb_north.inst.cb_conf_bus[309] ),
    .S(psn_net_16),
    .X(_03894_));
 sky130_fd_sc_hd__mux2_1 _06283_ (.A0(\cb_north.inst.cb_conf_bus[309] ),
    .A1(\cb_north.inst.cb_conf_bus[310] ),
    .S(psn_net_16),
    .X(_03896_));
 sky130_fd_sc_hd__mux2_1 _06284_ (.A0(\cb_north.inst.cb_conf_bus[310] ),
    .A1(\cb_north.inst.cb_conf_bus[311] ),
    .S(psn_net_16),
    .X(_03898_));
 sky130_fd_sc_hd__mux2_1 _06285_ (.A0(\cb_north.inst.cb_conf_bus[311] ),
    .A1(\cb_north.inst.cb_conf_bus[312] ),
    .S(psn_net_16),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _06286_ (.A0(\cb_north.inst.cb_conf_bus[312] ),
    .A1(\cb_north.inst.cb_conf_bus[313] ),
    .S(psn_net_16),
    .X(_03902_));
 sky130_fd_sc_hd__mux2_1 _06287_ (.A0(\cb_north.inst.cb_conf_bus[313] ),
    .A1(\cb_north.inst.cb_conf_bus[314] ),
    .S(psn_net_16),
    .X(_03904_));
 sky130_fd_sc_hd__mux2_1 _06288_ (.A0(\cb_north.inst.cb_conf_bus[314] ),
    .A1(\cb_north.inst.cb_conf_bus[315] ),
    .S(psn_net_16),
    .X(_03906_));
 sky130_fd_sc_hd__mux2_1 _06289_ (.A0(\cb_north.inst.cb_conf_bus[315] ),
    .A1(\cb_north.inst.cb_conf_bus[316] ),
    .S(psn_net_16),
    .X(_03908_));
 sky130_fd_sc_hd__mux2_1 _06290_ (.A0(\cb_north.inst.cb_conf_bus[316] ),
    .A1(\cb_north.inst.cb_conf_bus[317] ),
    .S(psn_net_16),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _06291_ (.A0(\cb_north.inst.cb_conf_bus[317] ),
    .A1(\cb_north.inst.cb_conf_bus[318] ),
    .S(psn_net_16),
    .X(_03912_));
 sky130_fd_sc_hd__mux2_1 _06292_ (.A0(\cb_north.inst.cb_conf_bus[318] ),
    .A1(\cb_north.inst.cb_conf_bus[319] ),
    .S(psn_net_16),
    .X(_03914_));
 sky130_fd_sc_hd__mux2_1 _06293_ (.A0(\cb_north.inst.cb_conf_bus[319] ),
    .A1(\cb_north.inst.cb_conf_bus[320] ),
    .S(psn_net_16),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_1 _06294_ (.A0(\cb_north.inst.cb_conf_bus[320] ),
    .A1(\cb_north.inst.cb_conf_bus[321] ),
    .S(psn_net_16),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _06295_ (.A0(\cb_north.inst.cb_conf_bus[321] ),
    .A1(\cb_north.inst.cb_conf_bus[322] ),
    .S(psn_net_16),
    .X(_03920_));
 sky130_fd_sc_hd__mux2_1 _06296_ (.A0(\cb_north.inst.cb_conf_bus[322] ),
    .A1(\cb_north.inst.cb_conf_bus[323] ),
    .S(psn_net_16),
    .X(_03922_));
 sky130_fd_sc_hd__mux2_1 _06297_ (.A0(\cb_north.inst.cb_conf_bus[323] ),
    .A1(\cb_north.inst.cb_conf_bus[324] ),
    .S(psn_net_16),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_1 _06298_ (.A0(\cb_north.inst.cb_conf_bus[324] ),
    .A1(\cb_north.inst.cb_conf_bus[325] ),
    .S(psn_net_16),
    .X(_03926_));
 sky130_fd_sc_hd__mux2_1 _06299_ (.A0(\cb_north.inst.cb_conf_bus[325] ),
    .A1(\cb_north.inst.cb_conf_bus[326] ),
    .S(psn_net_16),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_1 _06300_ (.A0(\cb_north.inst.cb_conf_bus[326] ),
    .A1(\cb_north.inst.cb_conf_bus[327] ),
    .S(psn_net_16),
    .X(_03930_));
 sky130_fd_sc_hd__mux2_1 _06301_ (.A0(\cb_north.inst.cb_conf_bus[327] ),
    .A1(\cb_north.inst.cb_conf_bus[328] ),
    .S(psn_net_16),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _06302_ (.A0(\cb_north.inst.cb_conf_bus[328] ),
    .A1(\cb_north.inst.cb_conf_bus[329] ),
    .S(psn_net_16),
    .X(_03934_));
 sky130_fd_sc_hd__mux2_1 _06303_ (.A0(\cb_north.inst.cb_conf_bus[329] ),
    .A1(\cb_north.inst.cb_conf_bus[330] ),
    .S(psn_net_16),
    .X(_03936_));
 sky130_fd_sc_hd__mux2_1 _06304_ (.A0(\cb_north.inst.cb_conf_bus[330] ),
    .A1(\cb_north.inst.cb_conf_bus[331] ),
    .S(psn_net_16),
    .X(_03938_));
 sky130_fd_sc_hd__mux2_1 _06305_ (.A0(\cb_north.inst.cb_conf_bus[331] ),
    .A1(\cb_north.inst.cb_conf_bus[332] ),
    .S(psn_net_16),
    .X(_03940_));
 sky130_fd_sc_hd__mux2_1 _06306_ (.A0(\cb_north.inst.cb_conf_bus[332] ),
    .A1(\cb_north.inst.cb_conf_bus[333] ),
    .S(psn_net_16),
    .X(_03942_));
 sky130_fd_sc_hd__mux2_1 _06307_ (.A0(\cb_north.inst.cb_conf_bus[333] ),
    .A1(\cb_north.inst.cb_conf_bus[334] ),
    .S(psn_net_16),
    .X(_03944_));
 sky130_fd_sc_hd__mux2_1 _06308_ (.A0(\cb_north.inst.cb_conf_bus[334] ),
    .A1(\cb_north.inst.cb_conf_bus[335] ),
    .S(psn_net_16),
    .X(_03946_));
 sky130_fd_sc_hd__mux2_1 _06309_ (.A0(\cb_north.inst.cb_conf_bus[335] ),
    .A1(\cb_north.inst.cb_conf_bus[336] ),
    .S(psn_net_16),
    .X(_03948_));
 sky130_fd_sc_hd__mux2_1 _06310_ (.A0(\cb_north.inst.cb_conf_bus[336] ),
    .A1(\cb_north.inst.cb_conf_bus[337] ),
    .S(psn_net_16),
    .X(_03950_));
 sky130_fd_sc_hd__mux2_1 _06311_ (.A0(\cb_north.inst.cb_conf_bus[337] ),
    .A1(\cb_north.inst.cb_conf_bus[338] ),
    .S(psn_net_16),
    .X(_03952_));
 sky130_fd_sc_hd__mux2_1 _06312_ (.A0(\cb_north.inst.cb_conf_bus[338] ),
    .A1(\cb_north.inst.cb_conf_bus[339] ),
    .S(psn_net_16),
    .X(_03954_));
 sky130_fd_sc_hd__mux2_1 _06313_ (.A0(\cb_north.inst.cb_conf_bus[339] ),
    .A1(\cb_north.inst.cb_conf_bus[340] ),
    .S(psn_net_16),
    .X(_03956_));
 sky130_fd_sc_hd__mux2_1 _06314_ (.A0(\cb_north.inst.cb_conf_bus[340] ),
    .A1(\cb_north.inst.cb_conf_bus[341] ),
    .S(psn_net_16),
    .X(_03958_));
 sky130_fd_sc_hd__mux2_1 _06315_ (.A0(\cb_north.inst.cb_conf_bus[341] ),
    .A1(\cb_north.inst.cb_conf_bus[342] ),
    .S(psn_net_17),
    .X(_03960_));
 sky130_fd_sc_hd__mux2_1 _06316_ (.A0(\cb_north.inst.cb_conf_bus[342] ),
    .A1(\cb_north.inst.cb_conf_bus[343] ),
    .S(psn_net_17),
    .X(_03962_));
 sky130_fd_sc_hd__mux2_1 _06317_ (.A0(\cb_north.inst.cb_conf_bus[343] ),
    .A1(\cb_north.inst.cb_conf_bus[344] ),
    .S(psn_net_17),
    .X(_03964_));
 sky130_fd_sc_hd__mux2_1 _06318_ (.A0(\cb_north.inst.cb_conf_bus[344] ),
    .A1(\cb_north.inst.cb_conf_bus[345] ),
    .S(psn_net_16),
    .X(_03966_));
 sky130_fd_sc_hd__mux2_1 _06319_ (.A0(\cb_north.inst.cb_conf_bus[345] ),
    .A1(\cb_north.inst.cb_conf_bus[346] ),
    .S(psn_net_16),
    .X(_03968_));
 sky130_fd_sc_hd__mux2_1 _06320_ (.A0(\cb_north.inst.cb_conf_bus[346] ),
    .A1(\cb_north.inst.cb_conf_bus[347] ),
    .S(psn_net_16),
    .X(_03970_));
 sky130_fd_sc_hd__mux2_1 _06321_ (.A0(\cb_north.inst.cb_conf_bus[347] ),
    .A1(\cb_north.inst.cb_conf_bus[348] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03972_));
 sky130_fd_sc_hd__mux2_1 _06322_ (.A0(\cb_north.inst.cb_conf_bus[348] ),
    .A1(\cb_north.inst.cb_conf_bus[349] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03974_));
 sky130_fd_sc_hd__mux2_1 _06323_ (.A0(\cb_north.inst.cb_conf_bus[349] ),
    .A1(\cb_north.inst.cb_conf_bus[350] ),
    .S(psn_net_15),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _06324_ (.A0(\cb_north.inst.cb_conf_bus[350] ),
    .A1(\cb_north.inst.cb_conf_bus[351] ),
    .S(psn_net_15),
    .X(_03978_));
 sky130_fd_sc_hd__mux2_1 _06325_ (.A0(\cb_north.inst.cb_conf_bus[351] ),
    .A1(\cb_north.inst.cb_conf_bus[352] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03980_));
 sky130_fd_sc_hd__mux2_1 _06326_ (.A0(\cb_north.inst.cb_conf_bus[352] ),
    .A1(\cb_north.inst.cb_conf_bus[353] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03982_));
 sky130_fd_sc_hd__mux2_1 _06327_ (.A0(\cb_north.inst.cb_conf_bus[353] ),
    .A1(\cb_north.inst.cb_conf_bus[354] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03984_));
 sky130_fd_sc_hd__mux2_1 _06328_ (.A0(\cb_north.inst.cb_conf_bus[354] ),
    .A1(\cb_north.inst.cb_conf_bus[355] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03986_));
 sky130_fd_sc_hd__mux2_1 _06329_ (.A0(\cb_north.inst.cb_conf_bus[355] ),
    .A1(\cb_north.inst.cb_conf_bus[356] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_1 _06330_ (.A0(\cb_north.inst.cb_conf_bus[356] ),
    .A1(\cb_north.inst.cb_conf_bus[357] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03990_));
 sky130_fd_sc_hd__mux2_1 _06331_ (.A0(\cb_north.inst.cb_conf_bus[357] ),
    .A1(\cb_north.inst.cb_conf_bus[358] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03992_));
 sky130_fd_sc_hd__mux2_1 _06332_ (.A0(\cb_north.inst.cb_conf_bus[358] ),
    .A1(\cb_north.inst.cb_conf_bus[359] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _06333_ (.A0(\cb_north.inst.cb_conf_bus[359] ),
    .A1(\cb_north.inst.cb_conf_bus[360] ),
    .S(psn_net_17),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_1 _06334_ (.A0(\cb_north.inst.cb_conf_bus[360] ),
    .A1(\cb_north.inst.cb_conf_bus[361] ),
    .S(psn_net_17),
    .X(_03998_));
 sky130_fd_sc_hd__mux2_1 _06335_ (.A0(\cb_north.inst.cb_conf_bus[361] ),
    .A1(\cb_north.inst.cb_conf_bus[362] ),
    .S(psn_net_17),
    .X(_04000_));
 sky130_fd_sc_hd__mux2_1 _06336_ (.A0(\cb_north.inst.cb_conf_bus[362] ),
    .A1(\cb_north.inst.cb_conf_bus[363] ),
    .S(psn_net_17),
    .X(_04002_));
 sky130_fd_sc_hd__mux2_1 _06337_ (.A0(\cb_north.inst.cb_conf_bus[363] ),
    .A1(\cb_north.inst.cb_conf_bus[364] ),
    .S(psn_net_17),
    .X(_04004_));
 sky130_fd_sc_hd__mux2_1 _06338_ (.A0(\cb_north.inst.cb_conf_bus[364] ),
    .A1(\cb_north.inst.cb_conf_bus[365] ),
    .S(psn_net_17),
    .X(_04006_));
 sky130_fd_sc_hd__mux2_1 _06339_ (.A0(\cb_north.inst.cb_conf_bus[365] ),
    .A1(\cb_north.inst.cb_conf_bus[366] ),
    .S(psn_net_17),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _06340_ (.A0(\cb_north.inst.cb_conf_bus[366] ),
    .A1(\cb_north.inst.cb_conf_bus[367] ),
    .S(psn_net_17),
    .X(_04010_));
 sky130_fd_sc_hd__mux2_1 _06341_ (.A0(\cb_north.inst.cb_conf_bus[367] ),
    .A1(\cb_north.inst.cb_conf_bus[368] ),
    .S(psn_net_17),
    .X(_04012_));
 sky130_fd_sc_hd__mux2_1 _06342_ (.A0(\cb_north.inst.cb_conf_bus[368] ),
    .A1(\cb_north.inst.cb_conf_bus[369] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_04014_));
 sky130_fd_sc_hd__mux2_1 _06343_ (.A0(\cb_north.inst.cb_conf_bus[369] ),
    .A1(\cb_north.inst.cb_conf_bus[370] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_04016_));
 sky130_fd_sc_hd__mux2_1 _06344_ (.A0(\cb_north.inst.cb_conf_bus[370] ),
    .A1(\cb_north.inst.cb_conf_bus[371] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_04018_));
 sky130_fd_sc_hd__mux2_1 _06345_ (.A0(\cb_north.inst.cb_conf_bus[371] ),
    .A1(\cb_north.inst.cb_conf_bus[372] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_04020_));
 sky130_fd_sc_hd__mux2_1 _06346_ (.A0(\cb_north.inst.cb_conf_bus[372] ),
    .A1(\cb_north.inst.cb_conf_bus[373] ),
    .S(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(_04022_));
 sky130_fd_sc_hd__mux2_1 _06347_ (.A0(\cb_north.inst.cb_conf_bus[373] ),
    .A1(\cb_north.inst.cb_conf_bus[374] ),
    .S(psn_net_10),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_1 _06348_ (.A0(\cb_north.inst.cb_conf_bus[374] ),
    .A1(\cb_north.inst.cb_conf_bus[375] ),
    .S(psn_net_10),
    .X(_04026_));
 sky130_fd_sc_hd__mux2_1 _06349_ (.A0(\cb_north.inst.cb_conf_bus[375] ),
    .A1(\cb_north.inst.cb_conf_bus[376] ),
    .S(psn_net_10),
    .X(_04028_));
 sky130_fd_sc_hd__mux2_1 _06350_ (.A0(\cb_north.inst.cb_conf_bus[376] ),
    .A1(\cb_north.inst.cb_conf_bus[377] ),
    .S(psn_net_10),
    .X(_04030_));
 sky130_fd_sc_hd__mux2_1 _06351_ (.A0(\cb_north.inst.cb_conf_bus[377] ),
    .A1(\cb_north.inst.cb_conf_bus[378] ),
    .S(psn_net_10),
    .X(_04032_));
 sky130_fd_sc_hd__mux2_1 _06352_ (.A0(\cb_north.inst.cb_conf_bus[378] ),
    .A1(\cb_north.inst.cb_conf_bus[379] ),
    .S(psn_net_10),
    .X(_04034_));
 sky130_fd_sc_hd__mux2_1 _06353_ (.A0(\cb_north.inst.cb_conf_bus[379] ),
    .A1(\cb_north.inst.cb_conf_bus[380] ),
    .S(psn_net_10),
    .X(_04036_));
 sky130_fd_sc_hd__mux2_1 _06354_ (.A0(\cb_north.inst.cb_conf_bus[380] ),
    .A1(\cb_north.inst.cb_conf_bus[381] ),
    .S(psn_net_10),
    .X(_04038_));
 sky130_fd_sc_hd__mux2_1 _06355_ (.A0(\cb_north.inst.cb_conf_bus[381] ),
    .A1(\cb_north.inst.cb_conf_bus[382] ),
    .S(psn_net_10),
    .X(_04040_));
 sky130_fd_sc_hd__mux2_1 _06356_ (.A0(\cb_north.inst.cb_conf_bus[382] ),
    .A1(\cb_north.inst.cb_conf_bus[383] ),
    .S(psn_net_10),
    .X(_04042_));
 sky130_fd_sc_hd__mux2_1 _06357_ (.A0(\cb_north.inst.cb_conf_bus[383] ),
    .A1(\cb_north.inst.cb_conf_bus[384] ),
    .S(psn_net_10),
    .X(_04044_));
 sky130_fd_sc_hd__mux2_1 _06358_ (.A0(\cb_north.inst.cb_conf_bus[384] ),
    .A1(\cb_north.inst.cb_conf_bus[385] ),
    .S(psn_net_10),
    .X(_04046_));
 sky130_fd_sc_hd__mux2_1 _06359_ (.A0(\cb_north.inst.cb_conf_bus[385] ),
    .A1(\cb_north.inst.cb_conf_bus[386] ),
    .S(psn_net_9),
    .X(_04048_));
 sky130_fd_sc_hd__mux2_1 _06360_ (.A0(\cb_north.inst.cb_conf_bus[386] ),
    .A1(\cb_north.inst.cb_conf_bus[387] ),
    .S(psn_net_9),
    .X(_04050_));
 sky130_fd_sc_hd__mux2_1 _06361_ (.A0(\cb_north.inst.cb_conf_bus[387] ),
    .A1(\cb_north.inst.cb_conf_bus[388] ),
    .S(psn_net_9),
    .X(_04052_));
 sky130_fd_sc_hd__mux2_1 _06362_ (.A0(\cb_north.inst.cb_conf_bus[388] ),
    .A1(\cb_north.inst.cb_conf_bus[389] ),
    .S(psn_net_9),
    .X(_04054_));
 sky130_fd_sc_hd__mux2_1 _06363_ (.A0(\cb_north.inst.cb_conf_bus[389] ),
    .A1(\cb_north.inst.cb_conf_bus[390] ),
    .S(psn_net_9),
    .X(_04056_));
 sky130_fd_sc_hd__mux2_1 _06364_ (.A0(\cb_north.inst.cb_conf_bus[390] ),
    .A1(\cb_north.inst.cb_conf_bus[391] ),
    .S(psn_net_9),
    .X(_04058_));
 sky130_fd_sc_hd__mux2_1 _06365_ (.A0(\cb_north.inst.cb_conf_bus[391] ),
    .A1(\cb_north.inst.cb_conf_bus[392] ),
    .S(psn_net_9),
    .X(_04060_));
 sky130_fd_sc_hd__mux2_1 _06366_ (.A0(\cb_north.inst.cb_conf_bus[392] ),
    .A1(\cb_north.inst.cb_conf_bus[393] ),
    .S(psn_net_9),
    .X(_04062_));
 sky130_fd_sc_hd__mux2_1 _06367_ (.A0(\cb_north.inst.cb_conf_bus[393] ),
    .A1(\cb_north.inst.cb_conf_bus[394] ),
    .S(psn_net_9),
    .X(_04064_));
 sky130_fd_sc_hd__mux2_1 _06368_ (.A0(\cb_north.inst.cb_conf_bus[394] ),
    .A1(\cb_north.inst.cb_conf_bus[395] ),
    .S(psn_net_9),
    .X(_04066_));
 sky130_fd_sc_hd__mux2_1 _06369_ (.A0(\cb_north.inst.cb_conf_bus[395] ),
    .A1(\cb_north.inst.cb_conf_bus[396] ),
    .S(psn_net_9),
    .X(_04068_));
 sky130_fd_sc_hd__mux2_1 _06370_ (.A0(\cb_north.inst.cb_conf_bus[396] ),
    .A1(\cb_north.inst.cb_conf_bus[397] ),
    .S(psn_net_9),
    .X(_04070_));
 sky130_fd_sc_hd__mux2_1 _06371_ (.A0(\cb_north.inst.cb_conf_bus[397] ),
    .A1(\cb_north.inst.cb_conf_bus[398] ),
    .S(psn_net_9),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_1 _06372_ (.A0(\cb_north.inst.cb_conf_bus[398] ),
    .A1(\cb_north.inst.cb_conf_bus[399] ),
    .S(psn_net_9),
    .X(_04074_));
 sky130_fd_sc_hd__mux2_1 _06373_ (.A0(\cb_north.inst.cb_conf_bus[399] ),
    .A1(\cb_north.inst.cb_conf_bus[400] ),
    .S(psn_net_9),
    .X(_04076_));
 sky130_fd_sc_hd__mux2_1 _06374_ (.A0(\cb_north.inst.cb_conf_bus[400] ),
    .A1(\cb_north.inst.cb_conf_bus[401] ),
    .S(psn_net_9),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _06375_ (.A0(\cb_north.inst.cb_conf_bus[401] ),
    .A1(\cb_north.inst.cb_conf_bus[402] ),
    .S(psn_net_9),
    .X(_04080_));
 sky130_fd_sc_hd__mux2_1 _06376_ (.A0(\cb_north.inst.cb_conf_bus[402] ),
    .A1(\cb_north.inst.cb_conf_bus[403] ),
    .S(psn_net_9),
    .X(_04082_));
 sky130_fd_sc_hd__mux2_1 _06377_ (.A0(\cb_north.inst.cb_conf_bus[403] ),
    .A1(\cb_north.inst.cb_conf_bus[404] ),
    .S(psn_net_9),
    .X(_04084_));
 sky130_fd_sc_hd__mux2_1 _06378_ (.A0(\cb_north.inst.cb_conf_bus[404] ),
    .A1(\cb_north.inst.cb_conf_bus[405] ),
    .S(psn_net_9),
    .X(_04086_));
 sky130_fd_sc_hd__mux2_1 _06379_ (.A0(\cb_north.inst.cb_conf_bus[405] ),
    .A1(\cb_north.inst.cb_conf_bus[406] ),
    .S(psn_net_9),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_1 _06380_ (.A0(\cb_north.inst.cb_conf_bus[406] ),
    .A1(\cb_north.inst.cb_conf_bus[407] ),
    .S(psn_net_9),
    .X(_04090_));
 sky130_fd_sc_hd__mux2_1 _06381_ (.A0(\cb_north.inst.cb_conf_bus[407] ),
    .A1(\cb_north.inst.cb_conf_bus[408] ),
    .S(psn_net_9),
    .X(_04092_));
 sky130_fd_sc_hd__mux2_1 _06382_ (.A0(\cb_north.inst.cb_conf_bus[408] ),
    .A1(\cb_north.inst.cb_conf_bus[409] ),
    .S(psn_net_9),
    .X(_04094_));
 sky130_fd_sc_hd__mux2_1 _06383_ (.A0(\cb_north.inst.cb_conf_bus[409] ),
    .A1(\cb_north.inst.cb_conf_bus[410] ),
    .S(psn_net_9),
    .X(_04096_));
 sky130_fd_sc_hd__mux2_1 _06384_ (.A0(\cb_north.inst.cb_conf_bus[410] ),
    .A1(\cb_north.inst.cb_conf_bus[411] ),
    .S(psn_net_9),
    .X(_04098_));
 sky130_fd_sc_hd__mux2_1 _06385_ (.A0(\cb_north.inst.cb_conf_bus[411] ),
    .A1(\cb_north.inst.cb_conf_bus[412] ),
    .S(psn_net_9),
    .X(_04100_));
 sky130_fd_sc_hd__mux2_1 _06386_ (.A0(\cb_north.inst.cb_conf_bus[412] ),
    .A1(\cb_north.inst.cb_conf_bus[413] ),
    .S(psn_net_9),
    .X(_04102_));
 sky130_fd_sc_hd__mux2_1 _06387_ (.A0(\cb_north.inst.cb_conf_bus[413] ),
    .A1(\cb_north.inst.cb_conf_bus[414] ),
    .S(psn_net_9),
    .X(_04104_));
 sky130_fd_sc_hd__mux2_1 _06388_ (.A0(\cb_north.inst.cb_conf_bus[414] ),
    .A1(\cb_north.inst.cb_conf_bus[415] ),
    .S(psn_net_9),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _06389_ (.A0(\cb_north.inst.cb_conf_bus[415] ),
    .A1(\cb_north.inst.cb_conf_bus[416] ),
    .S(psn_net_8),
    .X(_04108_));
 sky130_fd_sc_hd__mux2_1 _06390_ (.A0(\cb_north.inst.cb_conf_bus[416] ),
    .A1(\cb_north.inst.cb_conf_bus[417] ),
    .S(psn_net_8),
    .X(_04110_));
 sky130_fd_sc_hd__mux2_1 _06391_ (.A0(\cb_north.inst.cb_conf_bus[417] ),
    .A1(\cb_north.inst.cb_conf_bus[418] ),
    .S(psn_net_8),
    .X(_04112_));
 sky130_fd_sc_hd__mux2_1 _06392_ (.A0(\cb_north.inst.cb_conf_bus[418] ),
    .A1(\cb_north.inst.cb_conf_bus[419] ),
    .S(psn_net_8),
    .X(_04114_));
 sky130_fd_sc_hd__mux2_1 _06393_ (.A0(\cb_north.inst.cb_conf_bus[419] ),
    .A1(\cb_north.inst.configuroni.comb_shifter.config_data[420] ),
    .S(psn_net_8),
    .X(_04116_));
 sky130_fd_sc_hd__mux2_1 _06394_ (.A0(\cb_north.inst.configuroni.comb_shifter.config_data[420] ),
    .A1(\cb_north.inst.configuroni.comb_shifter.config_data[421] ),
    .S(psn_net_8),
    .X(_04118_));
 sky130_fd_sc_hd__mux2_1 _06395_ (.A0(_02038_),
    .A1(_01541_),
    .S(rst),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _06396_ (.A0(_02040_),
    .A1(_01540_),
    .S(rst),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _06397_ (.A0(_02042_),
    .A1(_01539_),
    .S(rst),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _06398_ (.A0(_02044_),
    .A1(_01538_),
    .S(rst),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _06399_ (.A0(_02046_),
    .A1(_01537_),
    .S(rst),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _06400_ (.A0(_02048_),
    .A1(_01536_),
    .S(rst),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _06401_ (.A0(_02050_),
    .A1(_01535_),
    .S(rst),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _06402_ (.A0(_02052_),
    .A1(_01534_),
    .S(rst),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _06403_ (.A0(_02054_),
    .A1(_01533_),
    .S(rst),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _06404_ (.A0(_02056_),
    .A1(_01532_),
    .S(rst),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _06405_ (.A0(_02058_),
    .A1(_01531_),
    .S(rst),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _06406_ (.A0(_02060_),
    .A1(_01530_),
    .S(rst),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _06407_ (.A0(_02062_),
    .A1(_01529_),
    .S(rst),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _06408_ (.A0(_02064_),
    .A1(_01528_),
    .S(rst),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _06409_ (.A0(_02066_),
    .A1(_01527_),
    .S(rst),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _06410_ (.A0(_02068_),
    .A1(_01526_),
    .S(rst),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _06411_ (.A0(_02070_),
    .A1(_01525_),
    .S(rst),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _06412_ (.A0(_02072_),
    .A1(_01524_),
    .S(rst),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _06413_ (.A0(_02074_),
    .A1(_01523_),
    .S(rst),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _06414_ (.A0(_02076_),
    .A1(_01522_),
    .S(rst),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _06415_ (.A0(_02078_),
    .A1(_01521_),
    .S(rst),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _06416_ (.A0(_02080_),
    .A1(_01520_),
    .S(rst),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _06417_ (.A0(_02082_),
    .A1(_01519_),
    .S(rst),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _06418_ (.A0(_02084_),
    .A1(_01518_),
    .S(rst),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _06419_ (.A0(_02086_),
    .A1(_01517_),
    .S(rst),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _06420_ (.A0(_02088_),
    .A1(_01516_),
    .S(rst),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _06421_ (.A0(_02090_),
    .A1(_01515_),
    .S(rst),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _06422_ (.A0(_02092_),
    .A1(_01514_),
    .S(rst),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _06423_ (.A0(_02094_),
    .A1(_01513_),
    .S(rst),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _06424_ (.A0(_02096_),
    .A1(_01512_),
    .S(rst),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _06425_ (.A0(_02098_),
    .A1(_01511_),
    .S(rst),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _06426_ (.A0(_02100_),
    .A1(_01510_),
    .S(rst),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _06427_ (.A0(_02102_),
    .A1(_01509_),
    .S(rst),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _06428_ (.A0(_02104_),
    .A1(_01508_),
    .S(rst),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _06429_ (.A0(_02106_),
    .A1(_01507_),
    .S(rst),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _06430_ (.A0(_02108_),
    .A1(_01506_),
    .S(rst),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _06431_ (.A0(_02110_),
    .A1(_01505_),
    .S(rst),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _06432_ (.A0(_02112_),
    .A1(_01504_),
    .S(rst),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _06433_ (.A0(_02114_),
    .A1(_01503_),
    .S(rst),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _06434_ (.A0(_02116_),
    .A1(_01502_),
    .S(rst),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _06435_ (.A0(_02118_),
    .A1(_01501_),
    .S(rst),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _06436_ (.A0(_02120_),
    .A1(_01500_),
    .S(rst),
    .X(_02121_));
 sky130_fd_sc_hd__mux2_1 _06437_ (.A0(_02122_),
    .A1(_01499_),
    .S(rst),
    .X(_02123_));
 sky130_fd_sc_hd__mux2_1 _06438_ (.A0(_02124_),
    .A1(_01498_),
    .S(rst),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _06439_ (.A0(_02126_),
    .A1(_01497_),
    .S(rst),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _06440_ (.A0(_02128_),
    .A1(_01496_),
    .S(rst),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _06441_ (.A0(_02130_),
    .A1(_01495_),
    .S(rst),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _06442_ (.A0(_02132_),
    .A1(_01494_),
    .S(rst),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _06443_ (.A0(_02134_),
    .A1(_01493_),
    .S(rst),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _06444_ (.A0(_02136_),
    .A1(_01492_),
    .S(rst),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _06445_ (.A0(_02138_),
    .A1(_01491_),
    .S(rst),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _06446_ (.A0(_02140_),
    .A1(_01490_),
    .S(rst),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _06447_ (.A0(_02142_),
    .A1(_01489_),
    .S(rst),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _06448_ (.A0(_02144_),
    .A1(_01488_),
    .S(rst),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _06449_ (.A0(_02146_),
    .A1(_01487_),
    .S(rst),
    .X(_02147_));
 sky130_fd_sc_hd__mux2_1 _06450_ (.A0(_02148_),
    .A1(_01486_),
    .S(rst),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _06451_ (.A0(_02150_),
    .A1(_01485_),
    .S(rst),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _06452_ (.A0(_02152_),
    .A1(_01484_),
    .S(rst),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _06453_ (.A0(_02154_),
    .A1(_01483_),
    .S(rst),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _06454_ (.A0(_02156_),
    .A1(_01482_),
    .S(rst),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _06455_ (.A0(_02158_),
    .A1(_01481_),
    .S(rst),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _06456_ (.A0(_02160_),
    .A1(_01480_),
    .S(rst),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_1 _06457_ (.A0(_02162_),
    .A1(_01479_),
    .S(rst),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _06458_ (.A0(_02164_),
    .A1(_01478_),
    .S(rst),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _06459_ (.A0(_02166_),
    .A1(_01477_),
    .S(rst),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _06460_ (.A0(_02168_),
    .A1(_01476_),
    .S(rst),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _06461_ (.A0(_02170_),
    .A1(_01475_),
    .S(rst),
    .X(_02171_));
 sky130_fd_sc_hd__mux2_1 _06462_ (.A0(_02172_),
    .A1(_01474_),
    .S(rst),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _06463_ (.A0(_02174_),
    .A1(_01473_),
    .S(rst),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _06464_ (.A0(_02176_),
    .A1(_01472_),
    .S(rst),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_1 _06465_ (.A0(_02178_),
    .A1(_01471_),
    .S(rst),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _06466_ (.A0(_02180_),
    .A1(_01470_),
    .S(rst),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _06467_ (.A0(_02182_),
    .A1(_01469_),
    .S(rst),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _06468_ (.A0(_02184_),
    .A1(_01468_),
    .S(rst),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _06469_ (.A0(_02186_),
    .A1(_01467_),
    .S(rst),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _06470_ (.A0(_02188_),
    .A1(_01466_),
    .S(rst),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _06471_ (.A0(_02190_),
    .A1(_01465_),
    .S(rst),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _06472_ (.A0(_02192_),
    .A1(_01464_),
    .S(rst),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _06473_ (.A0(_02194_),
    .A1(_01463_),
    .S(rst),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _06474_ (.A0(_02196_),
    .A1(_01462_),
    .S(rst),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _06475_ (.A0(_02198_),
    .A1(_01461_),
    .S(rst),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _06476_ (.A0(_02200_),
    .A1(_01460_),
    .S(rst),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _06477_ (.A0(_02202_),
    .A1(_01459_),
    .S(rst),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _06478_ (.A0(_02204_),
    .A1(_01458_),
    .S(rst),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _06479_ (.A0(_02206_),
    .A1(_01457_),
    .S(rst),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _06480_ (.A0(_02208_),
    .A1(_01456_),
    .S(rst),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _06481_ (.A0(_02210_),
    .A1(_01455_),
    .S(rst),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _06482_ (.A0(_02212_),
    .A1(_01454_),
    .S(rst),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _06483_ (.A0(_02214_),
    .A1(_01453_),
    .S(rst),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _06484_ (.A0(_02216_),
    .A1(_01452_),
    .S(rst),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _06485_ (.A0(_02218_),
    .A1(_01451_),
    .S(rst),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _06486_ (.A0(_02220_),
    .A1(_01450_),
    .S(rst),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _06487_ (.A0(_02222_),
    .A1(_01449_),
    .S(rst),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _06488_ (.A0(_02224_),
    .A1(_01448_),
    .S(rst),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(_02226_),
    .A1(_01447_),
    .S(rst),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _06490_ (.A0(_02228_),
    .A1(_01446_),
    .S(rst),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _06491_ (.A0(_02230_),
    .A1(_01445_),
    .S(rst),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _06492_ (.A0(_02232_),
    .A1(_01444_),
    .S(rst),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _06493_ (.A0(_02234_),
    .A1(_01443_),
    .S(rst),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _06494_ (.A0(_02236_),
    .A1(_01442_),
    .S(rst),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _06495_ (.A0(_02238_),
    .A1(_01441_),
    .S(rst),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _06496_ (.A0(_02240_),
    .A1(_01440_),
    .S(rst),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _06497_ (.A0(_02242_),
    .A1(_01439_),
    .S(rst),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _06498_ (.A0(_02244_),
    .A1(_01438_),
    .S(rst),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _06499_ (.A0(_02246_),
    .A1(_01437_),
    .S(rst),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _06500_ (.A0(_02248_),
    .A1(_01436_),
    .S(rst),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _06501_ (.A0(_02250_),
    .A1(_01435_),
    .S(rst),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _06502_ (.A0(_02252_),
    .A1(_01434_),
    .S(rst),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _06503_ (.A0(_02254_),
    .A1(_01433_),
    .S(rst),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _06504_ (.A0(_02256_),
    .A1(_01432_),
    .S(rst),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _06505_ (.A0(_02258_),
    .A1(_01431_),
    .S(rst),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _06506_ (.A0(_02260_),
    .A1(_01430_),
    .S(rst),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _06507_ (.A0(_02262_),
    .A1(_01429_),
    .S(rst),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _06508_ (.A0(_02264_),
    .A1(_01428_),
    .S(rst),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _06509_ (.A0(_02266_),
    .A1(_01427_),
    .S(rst),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _06510_ (.A0(_02268_),
    .A1(_01426_),
    .S(rst),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _06511_ (.A0(_02270_),
    .A1(_01425_),
    .S(rst),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _06512_ (.A0(_02272_),
    .A1(_01424_),
    .S(rst),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _06513_ (.A0(_02274_),
    .A1(_01423_),
    .S(rst),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _06514_ (.A0(_02276_),
    .A1(_01422_),
    .S(rst),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _06515_ (.A0(_02278_),
    .A1(_01421_),
    .S(rst),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _06516_ (.A0(_02280_),
    .A1(_01420_),
    .S(rst),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _06517_ (.A0(_02282_),
    .A1(_01419_),
    .S(rst),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _06518_ (.A0(_02284_),
    .A1(_01418_),
    .S(rst),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _06519_ (.A0(_02286_),
    .A1(_01417_),
    .S(rst),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _06520_ (.A0(_02288_),
    .A1(_01416_),
    .S(rst),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _06521_ (.A0(_02290_),
    .A1(_01415_),
    .S(rst),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _06522_ (.A0(_02292_),
    .A1(_01414_),
    .S(rst),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _06523_ (.A0(_02294_),
    .A1(_01413_),
    .S(rst),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _06524_ (.A0(_02296_),
    .A1(_01412_),
    .S(rst),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _06525_ (.A0(_02298_),
    .A1(_01411_),
    .S(rst),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _06526_ (.A0(_02300_),
    .A1(_01410_),
    .S(rst),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _06527_ (.A0(_02302_),
    .A1(_01409_),
    .S(rst),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _06528_ (.A0(_02304_),
    .A1(_01408_),
    .S(rst),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _06529_ (.A0(_02306_),
    .A1(_01407_),
    .S(rst),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _06530_ (.A0(_02308_),
    .A1(_01406_),
    .S(rst),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _06531_ (.A0(_02310_),
    .A1(_01405_),
    .S(rst),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _06532_ (.A0(_02312_),
    .A1(_01404_),
    .S(rst),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _06533_ (.A0(_02314_),
    .A1(_01403_),
    .S(rst),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _06534_ (.A0(_02316_),
    .A1(_01402_),
    .S(rst),
    .X(_02317_));
 sky130_fd_sc_hd__mux2_1 _06535_ (.A0(_02318_),
    .A1(_01401_),
    .S(rst),
    .X(_02319_));
 sky130_fd_sc_hd__mux2_1 _06536_ (.A0(_02320_),
    .A1(_01400_),
    .S(rst),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _06537_ (.A0(_02322_),
    .A1(_01399_),
    .S(rst),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _06538_ (.A0(_02324_),
    .A1(_01398_),
    .S(rst),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _06539_ (.A0(_02326_),
    .A1(_01397_),
    .S(rst),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _06540_ (.A0(_02328_),
    .A1(_01396_),
    .S(rst),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _06541_ (.A0(_02330_),
    .A1(_01395_),
    .S(rst),
    .X(_02331_));
 sky130_fd_sc_hd__mux2_1 _06542_ (.A0(_02332_),
    .A1(_01394_),
    .S(rst),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _06543_ (.A0(_02334_),
    .A1(_01393_),
    .S(rst),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _06544_ (.A0(_02336_),
    .A1(_01392_),
    .S(rst),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _06545_ (.A0(_02338_),
    .A1(_01391_),
    .S(rst),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _06546_ (.A0(_02340_),
    .A1(_01390_),
    .S(rst),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _06547_ (.A0(_02342_),
    .A1(_01389_),
    .S(rst),
    .X(_02343_));
 sky130_fd_sc_hd__mux2_1 _06548_ (.A0(_02344_),
    .A1(_01388_),
    .S(rst),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _06549_ (.A0(_02346_),
    .A1(_01387_),
    .S(rst),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _06550_ (.A0(_02348_),
    .A1(_01386_),
    .S(rst),
    .X(_02349_));
 sky130_fd_sc_hd__mux2_1 _06551_ (.A0(_02350_),
    .A1(_01385_),
    .S(rst),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _06552_ (.A0(_02352_),
    .A1(_01384_),
    .S(rst),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _06553_ (.A0(_02354_),
    .A1(_01383_),
    .S(rst),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _06554_ (.A0(_02356_),
    .A1(_01382_),
    .S(rst),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _06555_ (.A0(_02358_),
    .A1(_01381_),
    .S(rst),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _06556_ (.A0(_02360_),
    .A1(_01380_),
    .S(rst),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _06557_ (.A0(_02362_),
    .A1(_01379_),
    .S(rst),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _06558_ (.A0(_02364_),
    .A1(_01378_),
    .S(rst),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _06559_ (.A0(_02366_),
    .A1(_01377_),
    .S(rst),
    .X(_02367_));
 sky130_fd_sc_hd__mux2_1 _06560_ (.A0(_02368_),
    .A1(_01376_),
    .S(rst),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _06561_ (.A0(_02370_),
    .A1(_01375_),
    .S(rst),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _06562_ (.A0(_02372_),
    .A1(_01374_),
    .S(rst),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _06563_ (.A0(_02374_),
    .A1(_01373_),
    .S(rst),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _06564_ (.A0(_02376_),
    .A1(_01372_),
    .S(rst),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _06565_ (.A0(_02378_),
    .A1(_01371_),
    .S(rst),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _06566_ (.A0(_02380_),
    .A1(_01370_),
    .S(rst),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _06567_ (.A0(_02382_),
    .A1(_01369_),
    .S(rst),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _06568_ (.A0(_02384_),
    .A1(_01368_),
    .S(rst),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _06569_ (.A0(_02386_),
    .A1(_01367_),
    .S(rst),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _06570_ (.A0(_02388_),
    .A1(_01366_),
    .S(rst),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _06571_ (.A0(_02390_),
    .A1(_01365_),
    .S(rst),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _06572_ (.A0(_02392_),
    .A1(_01364_),
    .S(rst),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _06573_ (.A0(_02394_),
    .A1(_01363_),
    .S(rst),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _06574_ (.A0(_02396_),
    .A1(_01362_),
    .S(rst),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _06575_ (.A0(_02398_),
    .A1(_01361_),
    .S(rst),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _06576_ (.A0(_02400_),
    .A1(_01360_),
    .S(rst),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _06577_ (.A0(_02402_),
    .A1(_01359_),
    .S(rst),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _06578_ (.A0(_02404_),
    .A1(_01358_),
    .S(rst),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _06579_ (.A0(_02406_),
    .A1(_01357_),
    .S(rst),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _06580_ (.A0(_02408_),
    .A1(_01356_),
    .S(rst),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _06581_ (.A0(_02410_),
    .A1(_01355_),
    .S(rst),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _06582_ (.A0(_02412_),
    .A1(_01354_),
    .S(rst),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _06583_ (.A0(_02414_),
    .A1(_01353_),
    .S(rst),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _06584_ (.A0(_02416_),
    .A1(_01352_),
    .S(rst),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _06585_ (.A0(_02418_),
    .A1(_01351_),
    .S(rst),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _06586_ (.A0(_02420_),
    .A1(_01350_),
    .S(rst),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _06587_ (.A0(_02422_),
    .A1(_01349_),
    .S(rst),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _06588_ (.A0(_02424_),
    .A1(_01348_),
    .S(rst),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _06589_ (.A0(_02426_),
    .A1(_01347_),
    .S(rst),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _06590_ (.A0(_02428_),
    .A1(_01346_),
    .S(rst),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _06591_ (.A0(_02430_),
    .A1(_01345_),
    .S(rst),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _06592_ (.A0(_02432_),
    .A1(_01344_),
    .S(rst),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _06593_ (.A0(_02434_),
    .A1(_01343_),
    .S(rst),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _06594_ (.A0(_02436_),
    .A1(_01342_),
    .S(rst),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _06595_ (.A0(_02438_),
    .A1(_01341_),
    .S(rst),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _06596_ (.A0(_02440_),
    .A1(_01340_),
    .S(rst),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _06597_ (.A0(_02442_),
    .A1(_01339_),
    .S(rst),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _06598_ (.A0(_02444_),
    .A1(_01338_),
    .S(rst),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _06599_ (.A0(_02446_),
    .A1(_01337_),
    .S(rst),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _06600_ (.A0(_02448_),
    .A1(_01336_),
    .S(rst),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _06601_ (.A0(_02450_),
    .A1(_01335_),
    .S(rst),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _06602_ (.A0(_02452_),
    .A1(_01334_),
    .S(rst),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _06603_ (.A0(_02454_),
    .A1(_01333_),
    .S(rst),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _06604_ (.A0(_02456_),
    .A1(_01332_),
    .S(rst),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _06605_ (.A0(_02458_),
    .A1(_01331_),
    .S(rst),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _06606_ (.A0(_02460_),
    .A1(_01330_),
    .S(rst),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _06607_ (.A0(_02462_),
    .A1(_01329_),
    .S(rst),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _06608_ (.A0(_02464_),
    .A1(_01328_),
    .S(rst),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _06609_ (.A0(_02466_),
    .A1(_01327_),
    .S(rst),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _06610_ (.A0(_02468_),
    .A1(_01326_),
    .S(rst),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _06611_ (.A0(_02470_),
    .A1(_01325_),
    .S(rst),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _06612_ (.A0(_02472_),
    .A1(_01324_),
    .S(rst),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _06613_ (.A0(_02474_),
    .A1(_01323_),
    .S(rst),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _06614_ (.A0(_02476_),
    .A1(_01322_),
    .S(rst),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _06615_ (.A0(_02478_),
    .A1(_01321_),
    .S(rst),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _06616_ (.A0(_02480_),
    .A1(_01320_),
    .S(rst),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _06617_ (.A0(_02482_),
    .A1(_01319_),
    .S(rst),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _06618_ (.A0(_02484_),
    .A1(_01318_),
    .S(rst),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _06619_ (.A0(_02486_),
    .A1(_01317_),
    .S(rst),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _06620_ (.A0(_02488_),
    .A1(_01316_),
    .S(rst),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _06621_ (.A0(_02490_),
    .A1(_01315_),
    .S(rst),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _06622_ (.A0(_02492_),
    .A1(_01314_),
    .S(rst),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _06623_ (.A0(_02494_),
    .A1(_01313_),
    .S(rst),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _06624_ (.A0(_02496_),
    .A1(_01312_),
    .S(rst),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _06625_ (.A0(_02498_),
    .A1(_01311_),
    .S(rst),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _06626_ (.A0(_02500_),
    .A1(_01310_),
    .S(rst),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _06627_ (.A0(_02502_),
    .A1(_01309_),
    .S(rst),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _06628_ (.A0(_02504_),
    .A1(_01308_),
    .S(rst),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _06629_ (.A0(_02506_),
    .A1(_01307_),
    .S(rst),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _06630_ (.A0(_02508_),
    .A1(_01306_),
    .S(rst),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _06631_ (.A0(_02510_),
    .A1(_01305_),
    .S(rst),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _06632_ (.A0(_02512_),
    .A1(_01304_),
    .S(rst),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _06633_ (.A0(_02514_),
    .A1(_01303_),
    .S(rst),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _06634_ (.A0(_02516_),
    .A1(_01302_),
    .S(rst),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _06635_ (.A0(_02518_),
    .A1(_01301_),
    .S(rst),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _06636_ (.A0(_02520_),
    .A1(_01300_),
    .S(rst),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _06637_ (.A0(_02522_),
    .A1(_01299_),
    .S(rst),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _06638_ (.A0(_02524_),
    .A1(_01298_),
    .S(rst),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _06639_ (.A0(_02526_),
    .A1(_01297_),
    .S(rst),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _06640_ (.A0(_02528_),
    .A1(_01296_),
    .S(rst),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _06641_ (.A0(_02530_),
    .A1(_01295_),
    .S(rst),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _06642_ (.A0(_02532_),
    .A1(_01294_),
    .S(rst),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _06643_ (.A0(_02534_),
    .A1(_01293_),
    .S(rst),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _06644_ (.A0(_02536_),
    .A1(_01292_),
    .S(rst),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _06645_ (.A0(_02538_),
    .A1(_01291_),
    .S(rst),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _06646_ (.A0(_02540_),
    .A1(_01290_),
    .S(rst),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _06647_ (.A0(_02542_),
    .A1(_01289_),
    .S(rst),
    .X(_02543_));
 sky130_fd_sc_hd__mux2_1 _06648_ (.A0(_02544_),
    .A1(_01288_),
    .S(rst),
    .X(_02545_));
 sky130_fd_sc_hd__mux2_1 _06649_ (.A0(_02546_),
    .A1(_01287_),
    .S(rst),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _06650_ (.A0(_02548_),
    .A1(_01286_),
    .S(rst),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _06651_ (.A0(_02550_),
    .A1(_01285_),
    .S(rst),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _06652_ (.A0(_02552_),
    .A1(_01284_),
    .S(rst),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _06653_ (.A0(_02554_),
    .A1(_01283_),
    .S(rst),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _06654_ (.A0(_02556_),
    .A1(_01282_),
    .S(rst),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _06655_ (.A0(_02558_),
    .A1(_01281_),
    .S(rst),
    .X(_02559_));
 sky130_fd_sc_hd__mux2_1 _06656_ (.A0(_02560_),
    .A1(_01280_),
    .S(rst),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _06657_ (.A0(_02562_),
    .A1(_01279_),
    .S(rst),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _06658_ (.A0(_02564_),
    .A1(_01278_),
    .S(rst),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _06659_ (.A0(_02566_),
    .A1(_01277_),
    .S(rst),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _06660_ (.A0(_02568_),
    .A1(_01276_),
    .S(rst),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _06661_ (.A0(_02570_),
    .A1(_01275_),
    .S(rst),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _06662_ (.A0(_02572_),
    .A1(_01274_),
    .S(rst),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _06663_ (.A0(_02574_),
    .A1(_01273_),
    .S(rst),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _06664_ (.A0(_02576_),
    .A1(_01272_),
    .S(rst),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _06665_ (.A0(_02578_),
    .A1(_01271_),
    .S(rst),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _06666_ (.A0(_02580_),
    .A1(_01270_),
    .S(rst),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _06667_ (.A0(_02582_),
    .A1(_01269_),
    .S(rst),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _06668_ (.A0(_02584_),
    .A1(_01268_),
    .S(rst),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _06669_ (.A0(_02586_),
    .A1(_01267_),
    .S(rst),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _06670_ (.A0(_02588_),
    .A1(_01266_),
    .S(rst),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _06671_ (.A0(_02590_),
    .A1(_01265_),
    .S(rst),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _06672_ (.A0(_02592_),
    .A1(_01264_),
    .S(rst),
    .X(_02593_));
 sky130_fd_sc_hd__mux2_1 _06673_ (.A0(_02594_),
    .A1(_01263_),
    .S(rst),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _06674_ (.A0(_02596_),
    .A1(_01262_),
    .S(rst),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _06675_ (.A0(_02598_),
    .A1(_01261_),
    .S(rst),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _06676_ (.A0(_02600_),
    .A1(_01260_),
    .S(rst),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _06677_ (.A0(_02602_),
    .A1(_01259_),
    .S(rst),
    .X(_02603_));
 sky130_fd_sc_hd__mux2_1 _06678_ (.A0(_02604_),
    .A1(_01258_),
    .S(rst),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _06679_ (.A0(_02606_),
    .A1(_01257_),
    .S(rst),
    .X(_02607_));
 sky130_fd_sc_hd__mux2_1 _06680_ (.A0(_02608_),
    .A1(_01256_),
    .S(rst),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _06681_ (.A0(_02610_),
    .A1(_01255_),
    .S(rst),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _06682_ (.A0(_02612_),
    .A1(_01254_),
    .S(rst),
    .X(_02613_));
 sky130_fd_sc_hd__mux2_1 _06683_ (.A0(_02614_),
    .A1(_01253_),
    .S(rst),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _06684_ (.A0(_02616_),
    .A1(_01252_),
    .S(rst),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _06685_ (.A0(_02618_),
    .A1(_01251_),
    .S(rst),
    .X(_02619_));
 sky130_fd_sc_hd__mux2_1 _06686_ (.A0(_02620_),
    .A1(_01250_),
    .S(rst),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _06687_ (.A0(_02622_),
    .A1(_01249_),
    .S(rst),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _06688_ (.A0(_02624_),
    .A1(_01248_),
    .S(rst),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _06689_ (.A0(_02626_),
    .A1(_01247_),
    .S(rst),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _06690_ (.A0(_02628_),
    .A1(_01246_),
    .S(rst),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _06691_ (.A0(_02630_),
    .A1(_01245_),
    .S(rst),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _06692_ (.A0(_02632_),
    .A1(_01244_),
    .S(rst),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _06693_ (.A0(_02634_),
    .A1(_01243_),
    .S(rst),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _06694_ (.A0(_02636_),
    .A1(_01242_),
    .S(rst),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _06695_ (.A0(_02638_),
    .A1(_01241_),
    .S(rst),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _06696_ (.A0(_02640_),
    .A1(_01240_),
    .S(rst),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _06697_ (.A0(_02642_),
    .A1(_01239_),
    .S(rst),
    .X(_02643_));
 sky130_fd_sc_hd__mux2_1 _06698_ (.A0(_02644_),
    .A1(_01238_),
    .S(rst),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _06699_ (.A0(_02646_),
    .A1(_01237_),
    .S(rst),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _06700_ (.A0(_02648_),
    .A1(_01236_),
    .S(rst),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _06701_ (.A0(_02650_),
    .A1(_01235_),
    .S(rst),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _06702_ (.A0(_02652_),
    .A1(_01234_),
    .S(rst),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _06703_ (.A0(_02654_),
    .A1(_01233_),
    .S(rst),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _06704_ (.A0(_02656_),
    .A1(_01232_),
    .S(rst),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _06705_ (.A0(_02658_),
    .A1(_01231_),
    .S(rst),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _06706_ (.A0(_02660_),
    .A1(_01230_),
    .S(rst),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _06707_ (.A0(_02662_),
    .A1(_01229_),
    .S(rst),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _06708_ (.A0(_02664_),
    .A1(_01228_),
    .S(rst),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _06709_ (.A0(_02666_),
    .A1(_01227_),
    .S(rst),
    .X(_02667_));
 sky130_fd_sc_hd__mux2_1 _06710_ (.A0(_02668_),
    .A1(_01226_),
    .S(rst),
    .X(_02669_));
 sky130_fd_sc_hd__mux2_1 _06711_ (.A0(_02670_),
    .A1(_01225_),
    .S(rst),
    .X(_02671_));
 sky130_fd_sc_hd__mux2_1 _06712_ (.A0(_02672_),
    .A1(_01224_),
    .S(rst),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _06713_ (.A0(_02674_),
    .A1(_01223_),
    .S(rst),
    .X(_02675_));
 sky130_fd_sc_hd__mux2_1 _06714_ (.A0(_02676_),
    .A1(_01222_),
    .S(rst),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _06715_ (.A0(_02678_),
    .A1(_01221_),
    .S(rst),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _06716_ (.A0(_02680_),
    .A1(_01220_),
    .S(rst),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _06717_ (.A0(_02682_),
    .A1(_01219_),
    .S(rst),
    .X(_02683_));
 sky130_fd_sc_hd__mux2_1 _06718_ (.A0(_02684_),
    .A1(_01218_),
    .S(rst),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _06719_ (.A0(_02686_),
    .A1(_01217_),
    .S(rst),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _06720_ (.A0(_02688_),
    .A1(_01216_),
    .S(rst),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_1 _06721_ (.A0(_02690_),
    .A1(_01215_),
    .S(rst),
    .X(_02691_));
 sky130_fd_sc_hd__mux2_1 _06722_ (.A0(_02692_),
    .A1(_01214_),
    .S(rst),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _06723_ (.A0(_02694_),
    .A1(_01213_),
    .S(rst),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _06724_ (.A0(_02696_),
    .A1(_01212_),
    .S(rst),
    .X(_02697_));
 sky130_fd_sc_hd__mux2_1 _06725_ (.A0(_02698_),
    .A1(_01211_),
    .S(rst),
    .X(_02699_));
 sky130_fd_sc_hd__mux2_1 _06726_ (.A0(_02700_),
    .A1(_01210_),
    .S(rst),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _06727_ (.A0(_02702_),
    .A1(_01209_),
    .S(rst),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _06728_ (.A0(_02704_),
    .A1(_01208_),
    .S(rst),
    .X(_02705_));
 sky130_fd_sc_hd__mux2_1 _06729_ (.A0(_02706_),
    .A1(_01207_),
    .S(rst),
    .X(_02707_));
 sky130_fd_sc_hd__mux2_1 _06730_ (.A0(_02708_),
    .A1(_01206_),
    .S(rst),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _06731_ (.A0(_02710_),
    .A1(_01205_),
    .S(rst),
    .X(_02711_));
 sky130_fd_sc_hd__mux2_1 _06732_ (.A0(_02712_),
    .A1(_01204_),
    .S(rst),
    .X(_02713_));
 sky130_fd_sc_hd__mux2_1 _06733_ (.A0(_02714_),
    .A1(_01203_),
    .S(rst),
    .X(_02715_));
 sky130_fd_sc_hd__mux2_1 _06734_ (.A0(_02716_),
    .A1(_01202_),
    .S(rst),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_1 _06735_ (.A0(_02718_),
    .A1(_01201_),
    .S(rst),
    .X(_02719_));
 sky130_fd_sc_hd__mux2_1 _06736_ (.A0(_02720_),
    .A1(_01200_),
    .S(rst),
    .X(_02721_));
 sky130_fd_sc_hd__mux2_1 _06737_ (.A0(_02722_),
    .A1(_01199_),
    .S(rst),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _06738_ (.A0(_02724_),
    .A1(_01198_),
    .S(rst),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_1 _06739_ (.A0(_02726_),
    .A1(_01197_),
    .S(rst),
    .X(_02727_));
 sky130_fd_sc_hd__mux2_1 _06740_ (.A0(_02728_),
    .A1(_01196_),
    .S(rst),
    .X(_02729_));
 sky130_fd_sc_hd__mux2_1 _06741_ (.A0(_02730_),
    .A1(_01195_),
    .S(rst),
    .X(_02731_));
 sky130_fd_sc_hd__mux2_1 _06742_ (.A0(_02732_),
    .A1(_01194_),
    .S(rst),
    .X(_02733_));
 sky130_fd_sc_hd__mux2_1 _06743_ (.A0(_02734_),
    .A1(_01193_),
    .S(rst),
    .X(_02735_));
 sky130_fd_sc_hd__mux2_1 _06744_ (.A0(_02736_),
    .A1(_01192_),
    .S(rst),
    .X(_02737_));
 sky130_fd_sc_hd__mux2_1 _06745_ (.A0(_02738_),
    .A1(_01191_),
    .S(rst),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _06746_ (.A0(_02740_),
    .A1(_01190_),
    .S(rst),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _06747_ (.A0(_02742_),
    .A1(_01189_),
    .S(rst),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _06748_ (.A0(_02744_),
    .A1(_01188_),
    .S(rst),
    .X(_02745_));
 sky130_fd_sc_hd__mux2_1 _06749_ (.A0(_02746_),
    .A1(_01187_),
    .S(rst),
    .X(_02747_));
 sky130_fd_sc_hd__mux2_1 _06750_ (.A0(_02748_),
    .A1(_01186_),
    .S(rst),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _06751_ (.A0(_02750_),
    .A1(_01185_),
    .S(rst),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _06752_ (.A0(_02752_),
    .A1(_01184_),
    .S(rst),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _06753_ (.A0(_02754_),
    .A1(_01183_),
    .S(rst),
    .X(_02755_));
 sky130_fd_sc_hd__mux2_1 _06754_ (.A0(_02756_),
    .A1(_01182_),
    .S(rst),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _06755_ (.A0(_02758_),
    .A1(_01181_),
    .S(rst),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _06756_ (.A0(_02760_),
    .A1(_01180_),
    .S(rst),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _06757_ (.A0(_02762_),
    .A1(_01179_),
    .S(rst),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _06758_ (.A0(_02764_),
    .A1(_01178_),
    .S(rst),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _06759_ (.A0(_02766_),
    .A1(_01177_),
    .S(rst),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _06760_ (.A0(_02768_),
    .A1(_01176_),
    .S(rst),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _06761_ (.A0(_02770_),
    .A1(_01175_),
    .S(rst),
    .X(_02771_));
 sky130_fd_sc_hd__mux2_1 _06762_ (.A0(_02772_),
    .A1(_01174_),
    .S(rst),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _06763_ (.A0(_02774_),
    .A1(_01173_),
    .S(rst),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _06764_ (.A0(_02776_),
    .A1(_01172_),
    .S(rst),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _06765_ (.A0(_02778_),
    .A1(_01171_),
    .S(rst),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _06766_ (.A0(_02780_),
    .A1(_01170_),
    .S(rst),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _06767_ (.A0(_02782_),
    .A1(_01169_),
    .S(rst),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _06768_ (.A0(_02784_),
    .A1(_01168_),
    .S(rst),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _06769_ (.A0(_02786_),
    .A1(_01167_),
    .S(rst),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _06770_ (.A0(_02788_),
    .A1(_01166_),
    .S(rst),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _06771_ (.A0(_02790_),
    .A1(_01165_),
    .S(rst),
    .X(_02791_));
 sky130_fd_sc_hd__mux2_1 _06772_ (.A0(_02792_),
    .A1(_01164_),
    .S(rst),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _06773_ (.A0(_02794_),
    .A1(_01163_),
    .S(rst),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _06774_ (.A0(_02796_),
    .A1(_01162_),
    .S(rst),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _06775_ (.A0(_02798_),
    .A1(_01161_),
    .S(rst),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _06776_ (.A0(_02800_),
    .A1(_01160_),
    .S(rst),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _06777_ (.A0(_02802_),
    .A1(_01159_),
    .S(rst),
    .X(_02803_));
 sky130_fd_sc_hd__mux2_1 _06778_ (.A0(_02804_),
    .A1(_01158_),
    .S(rst),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _06779_ (.A0(_02806_),
    .A1(_01157_),
    .S(rst),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _06780_ (.A0(_02808_),
    .A1(_01156_),
    .S(rst),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _06781_ (.A0(_02810_),
    .A1(_01155_),
    .S(rst),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _06782_ (.A0(_02812_),
    .A1(_01154_),
    .S(rst),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _06783_ (.A0(_02814_),
    .A1(_01153_),
    .S(rst),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _06784_ (.A0(_02816_),
    .A1(_01152_),
    .S(rst),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _06785_ (.A0(_02818_),
    .A1(_01151_),
    .S(rst),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _06786_ (.A0(_02820_),
    .A1(_01150_),
    .S(rst),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _06787_ (.A0(_02822_),
    .A1(_01149_),
    .S(rst),
    .X(_02823_));
 sky130_fd_sc_hd__mux2_1 _06788_ (.A0(_02824_),
    .A1(_01148_),
    .S(rst),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _06789_ (.A0(_02826_),
    .A1(_01147_),
    .S(rst),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _06790_ (.A0(_02828_),
    .A1(_01146_),
    .S(rst),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_1 _06791_ (.A0(_02830_),
    .A1(_01145_),
    .S(rst),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _06792_ (.A0(_02832_),
    .A1(_01144_),
    .S(rst),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _06793_ (.A0(_02834_),
    .A1(_01143_),
    .S(rst),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _06794_ (.A0(_02836_),
    .A1(_01142_),
    .S(rst),
    .X(_02837_));
 sky130_fd_sc_hd__mux2_1 _06795_ (.A0(_02838_),
    .A1(_01141_),
    .S(rst),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _06796_ (.A0(_02840_),
    .A1(_01140_),
    .S(rst),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _06797_ (.A0(_02842_),
    .A1(_01139_),
    .S(rst),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _06798_ (.A0(_02844_),
    .A1(_01138_),
    .S(rst),
    .X(_02845_));
 sky130_fd_sc_hd__mux2_1 _06799_ (.A0(_02846_),
    .A1(_01137_),
    .S(rst),
    .X(_02847_));
 sky130_fd_sc_hd__mux2_1 _06800_ (.A0(_02848_),
    .A1(_01136_),
    .S(rst),
    .X(_02849_));
 sky130_fd_sc_hd__mux2_1 _06801_ (.A0(_02850_),
    .A1(_01135_),
    .S(rst),
    .X(_02851_));
 sky130_fd_sc_hd__mux2_1 _06802_ (.A0(_02852_),
    .A1(_01134_),
    .S(rst),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _06803_ (.A0(_02854_),
    .A1(_01133_),
    .S(rst),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_1 _06804_ (.A0(_02856_),
    .A1(_01132_),
    .S(rst),
    .X(_02857_));
 sky130_fd_sc_hd__mux2_1 _06805_ (.A0(_02858_),
    .A1(_01131_),
    .S(rst),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _06806_ (.A0(_02860_),
    .A1(_01130_),
    .S(rst),
    .X(_02861_));
 sky130_fd_sc_hd__mux2_1 _06807_ (.A0(_02862_),
    .A1(_01129_),
    .S(rst),
    .X(_02863_));
 sky130_fd_sc_hd__mux2_1 _06808_ (.A0(_02864_),
    .A1(_01128_),
    .S(rst),
    .X(_02865_));
 sky130_fd_sc_hd__mux2_1 _06809_ (.A0(_02866_),
    .A1(_01127_),
    .S(rst),
    .X(_02867_));
 sky130_fd_sc_hd__mux2_1 _06810_ (.A0(_02868_),
    .A1(_01126_),
    .S(rst),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _06811_ (.A0(_02870_),
    .A1(_01125_),
    .S(rst),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _06812_ (.A0(_02872_),
    .A1(_01124_),
    .S(rst),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _06813_ (.A0(_02874_),
    .A1(_01123_),
    .S(rst),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _06814_ (.A0(_02876_),
    .A1(_01122_),
    .S(rst),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _06815_ (.A0(_02878_),
    .A1(_01121_),
    .S(rst),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _06816_ (.A0(_02880_),
    .A1(_01120_),
    .S(rst),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _06817_ (.A0(_02882_),
    .A1(_01119_),
    .S(rst),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _06818_ (.A0(_02884_),
    .A1(_01118_),
    .S(rst),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(_02886_),
    .A1(_01117_),
    .S(rst),
    .X(_02887_));
 sky130_fd_sc_hd__mux2_1 _06820_ (.A0(_02888_),
    .A1(_01116_),
    .S(rst),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _06821_ (.A0(_02890_),
    .A1(_01115_),
    .S(rst),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _06822_ (.A0(_02892_),
    .A1(_01114_),
    .S(rst),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_1 _06823_ (.A0(_02894_),
    .A1(_01113_),
    .S(rst),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _06824_ (.A0(_02896_),
    .A1(_01112_),
    .S(rst),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _06825_ (.A0(_02898_),
    .A1(_01111_),
    .S(rst),
    .X(_02899_));
 sky130_fd_sc_hd__mux2_1 _06826_ (.A0(_02900_),
    .A1(_01110_),
    .S(rst),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _06827_ (.A0(_02902_),
    .A1(_01109_),
    .S(rst),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _06828_ (.A0(_02904_),
    .A1(_01108_),
    .S(rst),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _06829_ (.A0(_02906_),
    .A1(_01107_),
    .S(rst),
    .X(_02907_));
 sky130_fd_sc_hd__mux2_1 _06830_ (.A0(_02908_),
    .A1(_01106_),
    .S(rst),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _06831_ (.A0(_02910_),
    .A1(_01105_),
    .S(rst),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _06832_ (.A0(_02912_),
    .A1(_01104_),
    .S(rst),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _06833_ (.A0(_02914_),
    .A1(_01103_),
    .S(rst),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _06834_ (.A0(_02916_),
    .A1(_01102_),
    .S(rst),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _06835_ (.A0(_02918_),
    .A1(_01101_),
    .S(rst),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _06836_ (.A0(_02920_),
    .A1(_01100_),
    .S(rst),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _06837_ (.A0(_02922_),
    .A1(_01099_),
    .S(rst),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _06838_ (.A0(_02924_),
    .A1(_01098_),
    .S(rst),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _06839_ (.A0(_02926_),
    .A1(_01097_),
    .S(rst),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _06840_ (.A0(_02928_),
    .A1(_01096_),
    .S(rst),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _06841_ (.A0(_02930_),
    .A1(_01095_),
    .S(rst),
    .X(_02931_));
 sky130_fd_sc_hd__mux2_1 _06842_ (.A0(_02932_),
    .A1(_01094_),
    .S(rst),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _06843_ (.A0(_02934_),
    .A1(_01093_),
    .S(rst),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _06844_ (.A0(_02936_),
    .A1(_01092_),
    .S(rst),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _06845_ (.A0(_02938_),
    .A1(_01091_),
    .S(rst),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _06846_ (.A0(_02940_),
    .A1(_01090_),
    .S(rst),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _06847_ (.A0(_02942_),
    .A1(_01089_),
    .S(rst),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _06848_ (.A0(_02944_),
    .A1(_01088_),
    .S(rst),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(_02946_),
    .A1(_01087_),
    .S(rst),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _06850_ (.A0(_02948_),
    .A1(_01086_),
    .S(rst),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _06851_ (.A0(_02950_),
    .A1(_01085_),
    .S(rst),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _06852_ (.A0(_02952_),
    .A1(_01084_),
    .S(rst),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _06853_ (.A0(_02954_),
    .A1(_01083_),
    .S(rst),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _06854_ (.A0(_02956_),
    .A1(_01082_),
    .S(rst),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _06855_ (.A0(_02958_),
    .A1(_01081_),
    .S(rst),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _06856_ (.A0(_02960_),
    .A1(_01080_),
    .S(rst),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _06857_ (.A0(_02962_),
    .A1(_01079_),
    .S(rst),
    .X(_02963_));
 sky130_fd_sc_hd__mux2_1 _06858_ (.A0(_02964_),
    .A1(_01078_),
    .S(rst),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _06859_ (.A0(_02966_),
    .A1(_01077_),
    .S(rst),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _06860_ (.A0(_02968_),
    .A1(_01076_),
    .S(rst),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _06861_ (.A0(_02970_),
    .A1(_01075_),
    .S(rst),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _06862_ (.A0(_02972_),
    .A1(_01074_),
    .S(rst),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _06863_ (.A0(_02974_),
    .A1(_01073_),
    .S(rst),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _06864_ (.A0(_02976_),
    .A1(_01072_),
    .S(rst),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_1 _06865_ (.A0(_02978_),
    .A1(_01071_),
    .S(rst),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _06866_ (.A0(_02980_),
    .A1(_01070_),
    .S(rst),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _06867_ (.A0(_02982_),
    .A1(_01069_),
    .S(rst),
    .X(_02983_));
 sky130_fd_sc_hd__mux2_1 _06868_ (.A0(_02984_),
    .A1(_01068_),
    .S(rst),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _06869_ (.A0(_02986_),
    .A1(_01067_),
    .S(rst),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _06870_ (.A0(_02988_),
    .A1(_01066_),
    .S(rst),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_1 _06871_ (.A0(_02990_),
    .A1(_01065_),
    .S(rst),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _06872_ (.A0(_02992_),
    .A1(_01064_),
    .S(rst),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _06873_ (.A0(_02994_),
    .A1(_01063_),
    .S(rst),
    .X(_02995_));
 sky130_fd_sc_hd__mux2_1 _06874_ (.A0(_02996_),
    .A1(_01062_),
    .S(rst),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_1 _06875_ (.A0(_02998_),
    .A1(_01061_),
    .S(rst),
    .X(_02999_));
 sky130_fd_sc_hd__mux2_1 _06876_ (.A0(_03000_),
    .A1(_01060_),
    .S(rst),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _06877_ (.A0(_03002_),
    .A1(_01059_),
    .S(rst),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _06878_ (.A0(_03004_),
    .A1(_01058_),
    .S(rst),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_1 _06879_ (.A0(_03006_),
    .A1(_01057_),
    .S(rst),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _06880_ (.A0(_03008_),
    .A1(_01056_),
    .S(rst),
    .X(_03009_));
 sky130_fd_sc_hd__mux2_1 _06881_ (.A0(_03010_),
    .A1(_01055_),
    .S(rst),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _06882_ (.A0(_03012_),
    .A1(_01054_),
    .S(rst),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _06883_ (.A0(_03014_),
    .A1(_01053_),
    .S(rst),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _06884_ (.A0(_03016_),
    .A1(_01052_),
    .S(rst),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _06885_ (.A0(_03018_),
    .A1(_01051_),
    .S(rst),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _06886_ (.A0(_03020_),
    .A1(_01050_),
    .S(rst),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_1 _06887_ (.A0(_03022_),
    .A1(_01049_),
    .S(rst),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _06888_ (.A0(_03024_),
    .A1(_01048_),
    .S(rst),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _06889_ (.A0(_03026_),
    .A1(_01047_),
    .S(rst),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _06890_ (.A0(_03028_),
    .A1(_01046_),
    .S(rst),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _06891_ (.A0(_03030_),
    .A1(_01045_),
    .S(rst),
    .X(_03031_));
 sky130_fd_sc_hd__mux2_1 _06892_ (.A0(_03032_),
    .A1(_01044_),
    .S(rst),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _06893_ (.A0(_03034_),
    .A1(_01043_),
    .S(rst),
    .X(_03035_));
 sky130_fd_sc_hd__mux2_1 _06894_ (.A0(_03036_),
    .A1(_01042_),
    .S(rst),
    .X(_03037_));
 sky130_fd_sc_hd__mux2_1 _06895_ (.A0(_03038_),
    .A1(_01041_),
    .S(rst),
    .X(_03039_));
 sky130_fd_sc_hd__mux2_1 _06896_ (.A0(_03040_),
    .A1(_01040_),
    .S(rst),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _06897_ (.A0(_03042_),
    .A1(_01039_),
    .S(rst),
    .X(_03043_));
 sky130_fd_sc_hd__mux2_1 _06898_ (.A0(_03044_),
    .A1(_01038_),
    .S(rst),
    .X(_03045_));
 sky130_fd_sc_hd__mux2_1 _06899_ (.A0(_03046_),
    .A1(_01037_),
    .S(rst),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_1 _06900_ (.A0(_03048_),
    .A1(_01036_),
    .S(rst),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _06901_ (.A0(_03050_),
    .A1(_01035_),
    .S(rst),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _06902_ (.A0(_03052_),
    .A1(_01034_),
    .S(rst),
    .X(_03053_));
 sky130_fd_sc_hd__mux2_1 _06903_ (.A0(_03054_),
    .A1(_01033_),
    .S(rst),
    .X(_03055_));
 sky130_fd_sc_hd__mux2_1 _06904_ (.A0(_03056_),
    .A1(_01032_),
    .S(rst),
    .X(_03057_));
 sky130_fd_sc_hd__mux2_1 _06905_ (.A0(_03058_),
    .A1(_01031_),
    .S(rst),
    .X(_03059_));
 sky130_fd_sc_hd__mux2_1 _06906_ (.A0(_03060_),
    .A1(_01030_),
    .S(rst),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _06907_ (.A0(_03062_),
    .A1(_01029_),
    .S(rst),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _06908_ (.A0(_03064_),
    .A1(_01028_),
    .S(rst),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _06909_ (.A0(_03066_),
    .A1(_01027_),
    .S(rst),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _06910_ (.A0(_03068_),
    .A1(_01026_),
    .S(rst),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _06911_ (.A0(_03070_),
    .A1(_01025_),
    .S(rst),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _06912_ (.A0(_03072_),
    .A1(_01024_),
    .S(rst),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _06913_ (.A0(_03074_),
    .A1(_01023_),
    .S(rst),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _06914_ (.A0(_03076_),
    .A1(_01022_),
    .S(rst),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _06915_ (.A0(_03078_),
    .A1(_01021_),
    .S(rst),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _06916_ (.A0(_03080_),
    .A1(_01020_),
    .S(rst),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _06917_ (.A0(_03082_),
    .A1(_01019_),
    .S(rst),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _06918_ (.A0(_03084_),
    .A1(_01018_),
    .S(rst),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _06919_ (.A0(_03086_),
    .A1(_01017_),
    .S(rst),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _06920_ (.A0(_03088_),
    .A1(_01016_),
    .S(rst),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _06921_ (.A0(_03090_),
    .A1(_01015_),
    .S(rst),
    .X(_03091_));
 sky130_fd_sc_hd__mux2_1 _06922_ (.A0(_03092_),
    .A1(_01014_),
    .S(rst),
    .X(_03093_));
 sky130_fd_sc_hd__mux2_1 _06923_ (.A0(_03094_),
    .A1(_01013_),
    .S(rst),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _06924_ (.A0(_03096_),
    .A1(_01012_),
    .S(rst),
    .X(_03097_));
 sky130_fd_sc_hd__mux2_1 _06925_ (.A0(_03098_),
    .A1(_01011_),
    .S(rst),
    .X(_03099_));
 sky130_fd_sc_hd__mux2_1 _06926_ (.A0(_03100_),
    .A1(_01010_),
    .S(rst),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _06927_ (.A0(_03102_),
    .A1(_01009_),
    .S(rst),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _06928_ (.A0(_03104_),
    .A1(_01008_),
    .S(rst),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _06929_ (.A0(_03106_),
    .A1(_01007_),
    .S(rst),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _06930_ (.A0(_03108_),
    .A1(_01006_),
    .S(rst),
    .X(_03109_));
 sky130_fd_sc_hd__mux2_1 _06931_ (.A0(_03110_),
    .A1(_01005_),
    .S(rst),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _06932_ (.A0(_03112_),
    .A1(_01004_),
    .S(rst),
    .X(_03113_));
 sky130_fd_sc_hd__mux2_1 _06933_ (.A0(_03114_),
    .A1(_01003_),
    .S(rst),
    .X(_03115_));
 sky130_fd_sc_hd__mux2_1 _06934_ (.A0(_03116_),
    .A1(_01002_),
    .S(rst),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _06935_ (.A0(_03118_),
    .A1(_01001_),
    .S(rst),
    .X(_03119_));
 sky130_fd_sc_hd__mux2_1 _06936_ (.A0(_03120_),
    .A1(_01000_),
    .S(rst),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_1 _06937_ (.A0(_03122_),
    .A1(_00999_),
    .S(rst),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _06938_ (.A0(_03124_),
    .A1(_00998_),
    .S(rst),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _06939_ (.A0(_03126_),
    .A1(_00997_),
    .S(rst),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_1 _06940_ (.A0(_03128_),
    .A1(_00996_),
    .S(rst),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_1 _06941_ (.A0(_03130_),
    .A1(_00995_),
    .S(rst),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_1 _06942_ (.A0(_03132_),
    .A1(_00994_),
    .S(rst),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_1 _06943_ (.A0(_03134_),
    .A1(_00993_),
    .S(rst),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_1 _06944_ (.A0(_03136_),
    .A1(_00992_),
    .S(rst),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_1 _06945_ (.A0(_03138_),
    .A1(_00991_),
    .S(rst),
    .X(_03139_));
 sky130_fd_sc_hd__mux2_1 _06946_ (.A0(_03140_),
    .A1(_00990_),
    .S(rst),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _06947_ (.A0(_03142_),
    .A1(_00989_),
    .S(rst),
    .X(_03143_));
 sky130_fd_sc_hd__mux2_1 _06948_ (.A0(_03144_),
    .A1(_00988_),
    .S(rst),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _06949_ (.A0(_03146_),
    .A1(_00987_),
    .S(rst),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_1 _06950_ (.A0(_03148_),
    .A1(_00986_),
    .S(rst),
    .X(_03149_));
 sky130_fd_sc_hd__mux2_1 _06951_ (.A0(_03150_),
    .A1(_00985_),
    .S(rst),
    .X(_03151_));
 sky130_fd_sc_hd__mux2_1 _06952_ (.A0(_03152_),
    .A1(_00984_),
    .S(rst),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_1 _06953_ (.A0(_03154_),
    .A1(_00983_),
    .S(rst),
    .X(_03155_));
 sky130_fd_sc_hd__mux2_1 _06954_ (.A0(_03156_),
    .A1(_00982_),
    .S(rst),
    .X(_03157_));
 sky130_fd_sc_hd__mux2_1 _06955_ (.A0(_03158_),
    .A1(_02022_),
    .S(rst),
    .X(_03159_));
 sky130_fd_sc_hd__mux2_1 _06956_ (.A0(_03160_),
    .A1(_02021_),
    .S(rst),
    .X(_03161_));
 sky130_fd_sc_hd__mux2_1 _06957_ (.A0(_03162_),
    .A1(_02020_),
    .S(rst),
    .X(_03163_));
 sky130_fd_sc_hd__mux2_1 _06958_ (.A0(_03164_),
    .A1(_02019_),
    .S(rst),
    .X(_03165_));
 sky130_fd_sc_hd__mux2_1 _06959_ (.A0(_03166_),
    .A1(_02018_),
    .S(rst),
    .X(_03167_));
 sky130_fd_sc_hd__mux2_1 _06960_ (.A0(_03168_),
    .A1(_02017_),
    .S(rst),
    .X(_03169_));
 sky130_fd_sc_hd__mux2_1 _06961_ (.A0(_03170_),
    .A1(_02016_),
    .S(rst),
    .X(_03171_));
 sky130_fd_sc_hd__mux2_1 _06962_ (.A0(_03172_),
    .A1(_02015_),
    .S(rst),
    .X(_03173_));
 sky130_fd_sc_hd__mux2_1 _06963_ (.A0(_03174_),
    .A1(_02014_),
    .S(rst),
    .X(_03175_));
 sky130_fd_sc_hd__mux2_1 _06964_ (.A0(_03176_),
    .A1(_02013_),
    .S(rst),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _06965_ (.A0(_03178_),
    .A1(_02012_),
    .S(rst),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_1 _06966_ (.A0(_03180_),
    .A1(_02011_),
    .S(rst),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _06967_ (.A0(_03182_),
    .A1(_02010_),
    .S(rst),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _06968_ (.A0(_03184_),
    .A1(_02009_),
    .S(rst),
    .X(_03185_));
 sky130_fd_sc_hd__mux2_1 _06969_ (.A0(_03186_),
    .A1(_02008_),
    .S(rst),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_1 _06970_ (.A0(_03188_),
    .A1(_02007_),
    .S(rst),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _06971_ (.A0(_03190_),
    .A1(_02006_),
    .S(rst),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _06972_ (.A0(_03192_),
    .A1(_02005_),
    .S(rst),
    .X(_03193_));
 sky130_fd_sc_hd__mux2_1 _06973_ (.A0(_03194_),
    .A1(_02004_),
    .S(rst),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _06974_ (.A0(_03196_),
    .A1(_02003_),
    .S(rst),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _06975_ (.A0(_03198_),
    .A1(_02002_),
    .S(rst),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_1 _06976_ (.A0(_03200_),
    .A1(_02001_),
    .S(rst),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _06977_ (.A0(_03202_),
    .A1(_02000_),
    .S(rst),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _06978_ (.A0(_03204_),
    .A1(_01999_),
    .S(rst),
    .X(_03205_));
 sky130_fd_sc_hd__mux2_1 _06979_ (.A0(_03206_),
    .A1(_01998_),
    .S(rst),
    .X(_03207_));
 sky130_fd_sc_hd__mux2_1 _06980_ (.A0(_03208_),
    .A1(_01997_),
    .S(rst),
    .X(_03209_));
 sky130_fd_sc_hd__mux2_1 _06981_ (.A0(_03210_),
    .A1(_01996_),
    .S(rst),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _06982_ (.A0(_03212_),
    .A1(_01995_),
    .S(rst),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _06983_ (.A0(_03214_),
    .A1(_01994_),
    .S(rst),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _06984_ (.A0(_03216_),
    .A1(_01993_),
    .S(rst),
    .X(_03217_));
 sky130_fd_sc_hd__mux2_1 _06985_ (.A0(_03218_),
    .A1(_01992_),
    .S(rst),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _06986_ (.A0(_03220_),
    .A1(_01991_),
    .S(rst),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _06987_ (.A0(_03222_),
    .A1(_01990_),
    .S(rst),
    .X(_03223_));
 sky130_fd_sc_hd__mux2_1 _06988_ (.A0(_03224_),
    .A1(_01989_),
    .S(rst),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _06989_ (.A0(_03226_),
    .A1(_01988_),
    .S(rst),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _06990_ (.A0(_03228_),
    .A1(_01987_),
    .S(rst),
    .X(_03229_));
 sky130_fd_sc_hd__mux2_1 _06991_ (.A0(_03230_),
    .A1(_01986_),
    .S(rst),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _06992_ (.A0(_03232_),
    .A1(_01985_),
    .S(rst),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _06993_ (.A0(_03234_),
    .A1(_01984_),
    .S(rst),
    .X(_03235_));
 sky130_fd_sc_hd__mux2_1 _06994_ (.A0(_03236_),
    .A1(_01983_),
    .S(rst),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _06995_ (.A0(_03238_),
    .A1(_01982_),
    .S(rst),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _06996_ (.A0(_03240_),
    .A1(_01981_),
    .S(rst),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _06997_ (.A0(_03242_),
    .A1(_01980_),
    .S(rst),
    .X(_03243_));
 sky130_fd_sc_hd__mux2_1 _06998_ (.A0(_03244_),
    .A1(_01979_),
    .S(rst),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _06999_ (.A0(_03246_),
    .A1(_01978_),
    .S(rst),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _07000_ (.A0(_03248_),
    .A1(_01977_),
    .S(rst),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_1 _07001_ (.A0(_03250_),
    .A1(_01976_),
    .S(rst),
    .X(_03251_));
 sky130_fd_sc_hd__mux2_1 _07002_ (.A0(_03252_),
    .A1(_01975_),
    .S(rst),
    .X(_03253_));
 sky130_fd_sc_hd__mux2_1 _07003_ (.A0(_03254_),
    .A1(_01974_),
    .S(rst),
    .X(_03255_));
 sky130_fd_sc_hd__mux2_1 _07004_ (.A0(_03256_),
    .A1(_01973_),
    .S(rst),
    .X(_03257_));
 sky130_fd_sc_hd__mux2_1 _07005_ (.A0(_03258_),
    .A1(_01972_),
    .S(rst),
    .X(_03259_));
 sky130_fd_sc_hd__mux2_1 _07006_ (.A0(_03260_),
    .A1(_01971_),
    .S(rst),
    .X(_03261_));
 sky130_fd_sc_hd__mux2_1 _07007_ (.A0(_03262_),
    .A1(_01970_),
    .S(rst),
    .X(_03263_));
 sky130_fd_sc_hd__mux2_1 _07008_ (.A0(_03264_),
    .A1(_01969_),
    .S(rst),
    .X(_03265_));
 sky130_fd_sc_hd__mux2_1 _07009_ (.A0(_03266_),
    .A1(_01968_),
    .S(rst),
    .X(_03267_));
 sky130_fd_sc_hd__mux2_1 _07010_ (.A0(_03268_),
    .A1(_01967_),
    .S(rst),
    .X(_03269_));
 sky130_fd_sc_hd__mux2_1 _07011_ (.A0(_03270_),
    .A1(_01966_),
    .S(rst),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _07012_ (.A0(_03272_),
    .A1(_01965_),
    .S(rst),
    .X(_03273_));
 sky130_fd_sc_hd__mux2_1 _07013_ (.A0(_03274_),
    .A1(_01964_),
    .S(rst),
    .X(_03275_));
 sky130_fd_sc_hd__mux2_1 _07014_ (.A0(_03276_),
    .A1(_01963_),
    .S(rst),
    .X(_03277_));
 sky130_fd_sc_hd__mux2_1 _07015_ (.A0(_03278_),
    .A1(_01962_),
    .S(rst),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_1 _07016_ (.A0(_03280_),
    .A1(_01961_),
    .S(rst),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(_03282_),
    .A1(_01960_),
    .S(rst),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _07018_ (.A0(_03284_),
    .A1(_01959_),
    .S(rst),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _07019_ (.A0(_03286_),
    .A1(_01958_),
    .S(rst),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(_03288_),
    .A1(_01957_),
    .S(rst),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _07021_ (.A0(_03290_),
    .A1(_01956_),
    .S(rst),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _07022_ (.A0(_03292_),
    .A1(_01955_),
    .S(rst),
    .X(_03293_));
 sky130_fd_sc_hd__mux2_1 _07023_ (.A0(_03294_),
    .A1(_01954_),
    .S(rst),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(_03296_),
    .A1(_01953_),
    .S(rst),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _07025_ (.A0(_03298_),
    .A1(_01952_),
    .S(rst),
    .X(_03299_));
 sky130_fd_sc_hd__mux2_1 _07026_ (.A0(_03300_),
    .A1(_01951_),
    .S(rst),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(_03302_),
    .A1(_01950_),
    .S(rst),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _07028_ (.A0(_03304_),
    .A1(_01949_),
    .S(rst),
    .X(_03305_));
 sky130_fd_sc_hd__mux2_1 _07029_ (.A0(_03306_),
    .A1(_01948_),
    .S(rst),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _07030_ (.A0(_03308_),
    .A1(_01947_),
    .S(rst),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _07031_ (.A0(_03310_),
    .A1(_01946_),
    .S(rst),
    .X(_03311_));
 sky130_fd_sc_hd__mux2_1 _07032_ (.A0(_03312_),
    .A1(_01945_),
    .S(rst),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _07033_ (.A0(_03314_),
    .A1(_01944_),
    .S(rst),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _07034_ (.A0(_03316_),
    .A1(_01943_),
    .S(rst),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(_03318_),
    .A1(_01942_),
    .S(rst),
    .X(_03319_));
 sky130_fd_sc_hd__mux2_1 _07036_ (.A0(_03320_),
    .A1(_01941_),
    .S(rst),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(_03322_),
    .A1(_01940_),
    .S(rst),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _07038_ (.A0(_03324_),
    .A1(_01939_),
    .S(rst),
    .X(_03325_));
 sky130_fd_sc_hd__mux2_1 _07039_ (.A0(_03326_),
    .A1(_01938_),
    .S(rst),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _07040_ (.A0(_03328_),
    .A1(_01937_),
    .S(rst),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _07041_ (.A0(_03330_),
    .A1(_01936_),
    .S(rst),
    .X(_03331_));
 sky130_fd_sc_hd__mux2_1 _07042_ (.A0(_03332_),
    .A1(_01935_),
    .S(rst),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _07043_ (.A0(_03334_),
    .A1(_01934_),
    .S(rst),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(_03336_),
    .A1(_01933_),
    .S(rst),
    .X(_03337_));
 sky130_fd_sc_hd__mux2_1 _07045_ (.A0(_03338_),
    .A1(_01932_),
    .S(rst),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(_03340_),
    .A1(_01931_),
    .S(rst),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(_03342_),
    .A1(_01930_),
    .S(rst),
    .X(_03343_));
 sky130_fd_sc_hd__mux2_1 _07048_ (.A0(_03344_),
    .A1(_01929_),
    .S(rst),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _07049_ (.A0(_03346_),
    .A1(_01928_),
    .S(rst),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(_03348_),
    .A1(_01927_),
    .S(rst),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(_03350_),
    .A1(_01926_),
    .S(rst),
    .X(_03351_));
 sky130_fd_sc_hd__mux2_1 _07052_ (.A0(_03352_),
    .A1(_01925_),
    .S(rst),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _07053_ (.A0(_03354_),
    .A1(_01924_),
    .S(rst),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _07054_ (.A0(_03356_),
    .A1(_01923_),
    .S(rst),
    .X(_03357_));
 sky130_fd_sc_hd__mux2_1 _07055_ (.A0(_03358_),
    .A1(_01922_),
    .S(rst),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _07056_ (.A0(_03360_),
    .A1(_01921_),
    .S(rst),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _07057_ (.A0(_03362_),
    .A1(_01920_),
    .S(rst),
    .X(_03363_));
 sky130_fd_sc_hd__mux2_1 _07058_ (.A0(_03364_),
    .A1(_01919_),
    .S(rst),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _07059_ (.A0(_03366_),
    .A1(_01918_),
    .S(rst),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _07060_ (.A0(_03368_),
    .A1(_01917_),
    .S(rst),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_1 _07061_ (.A0(_03370_),
    .A1(_01916_),
    .S(rst),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _07062_ (.A0(_03372_),
    .A1(_01915_),
    .S(rst),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _07063_ (.A0(_03374_),
    .A1(_01914_),
    .S(rst),
    .X(_03375_));
 sky130_fd_sc_hd__mux2_1 _07064_ (.A0(_03376_),
    .A1(_01913_),
    .S(rst),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _07065_ (.A0(_03378_),
    .A1(_01912_),
    .S(rst),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _07066_ (.A0(_03380_),
    .A1(_01911_),
    .S(rst),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _07067_ (.A0(_03382_),
    .A1(_01910_),
    .S(rst),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _07068_ (.A0(_03384_),
    .A1(_01909_),
    .S(rst),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_1 _07069_ (.A0(_03386_),
    .A1(_01908_),
    .S(rst),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _07070_ (.A0(_03388_),
    .A1(_01907_),
    .S(rst),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_1 _07071_ (.A0(_03390_),
    .A1(_01906_),
    .S(rst),
    .X(_03391_));
 sky130_fd_sc_hd__mux2_1 _07072_ (.A0(_03392_),
    .A1(_01905_),
    .S(rst),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _07073_ (.A0(_03394_),
    .A1(_01904_),
    .S(rst),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_1 _07074_ (.A0(_03396_),
    .A1(_01903_),
    .S(rst),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _07075_ (.A0(_03398_),
    .A1(_01902_),
    .S(rst),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _07076_ (.A0(_03400_),
    .A1(_01901_),
    .S(rst),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_1 _07077_ (.A0(_03402_),
    .A1(_01900_),
    .S(rst),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _07078_ (.A0(_03404_),
    .A1(_01899_),
    .S(rst),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_1 _07079_ (.A0(_03406_),
    .A1(_01898_),
    .S(rst),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _07080_ (.A0(_03408_),
    .A1(_01897_),
    .S(rst),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _07081_ (.A0(_03410_),
    .A1(_01896_),
    .S(rst),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _07082_ (.A0(_03412_),
    .A1(_01895_),
    .S(rst),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _07083_ (.A0(_03414_),
    .A1(_01894_),
    .S(rst),
    .X(_03415_));
 sky130_fd_sc_hd__mux2_1 _07084_ (.A0(_03416_),
    .A1(_01893_),
    .S(rst),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _07085_ (.A0(_03418_),
    .A1(_01892_),
    .S(rst),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _07086_ (.A0(_03420_),
    .A1(_01891_),
    .S(rst),
    .X(_03421_));
 sky130_fd_sc_hd__mux2_1 _07087_ (.A0(_03422_),
    .A1(_01890_),
    .S(rst),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _07088_ (.A0(_03424_),
    .A1(_01889_),
    .S(rst),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(_03426_),
    .A1(_01888_),
    .S(rst),
    .X(_03427_));
 sky130_fd_sc_hd__mux2_1 _07090_ (.A0(_03428_),
    .A1(_01887_),
    .S(rst),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _07091_ (.A0(_03430_),
    .A1(_01886_),
    .S(rst),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _07092_ (.A0(_03432_),
    .A1(_01885_),
    .S(rst),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _07093_ (.A0(_03434_),
    .A1(_01884_),
    .S(rst),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _07094_ (.A0(_03436_),
    .A1(_01883_),
    .S(rst),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _07095_ (.A0(_03438_),
    .A1(_01882_),
    .S(rst),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(_03440_),
    .A1(_01881_),
    .S(rst),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _07097_ (.A0(_03442_),
    .A1(_01880_),
    .S(rst),
    .X(_03443_));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(_03444_),
    .A1(_01879_),
    .S(rst),
    .X(_03445_));
 sky130_fd_sc_hd__mux2_1 _07099_ (.A0(_03446_),
    .A1(_01878_),
    .S(rst),
    .X(_03447_));
 sky130_fd_sc_hd__mux2_1 _07100_ (.A0(_03448_),
    .A1(_01877_),
    .S(rst),
    .X(_03449_));
 sky130_fd_sc_hd__mux2_1 _07101_ (.A0(_03450_),
    .A1(_01876_),
    .S(rst),
    .X(_03451_));
 sky130_fd_sc_hd__mux2_1 _07102_ (.A0(_03452_),
    .A1(_01875_),
    .S(rst),
    .X(_03453_));
 sky130_fd_sc_hd__mux2_1 _07103_ (.A0(_03454_),
    .A1(_01874_),
    .S(rst),
    .X(_03455_));
 sky130_fd_sc_hd__mux2_1 _07104_ (.A0(_03456_),
    .A1(_01873_),
    .S(rst),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_1 _07105_ (.A0(_03458_),
    .A1(_01872_),
    .S(rst),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _07106_ (.A0(_03460_),
    .A1(_01871_),
    .S(rst),
    .X(_03461_));
 sky130_fd_sc_hd__mux2_1 _07107_ (.A0(_03462_),
    .A1(_01870_),
    .S(rst),
    .X(_03463_));
 sky130_fd_sc_hd__mux2_1 _07108_ (.A0(_03464_),
    .A1(_01869_),
    .S(rst),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_1 _07109_ (.A0(_03466_),
    .A1(_01868_),
    .S(rst),
    .X(_03467_));
 sky130_fd_sc_hd__mux2_1 _07110_ (.A0(_03468_),
    .A1(_01867_),
    .S(rst),
    .X(_03469_));
 sky130_fd_sc_hd__mux2_1 _07111_ (.A0(_03470_),
    .A1(_01866_),
    .S(rst),
    .X(_03471_));
 sky130_fd_sc_hd__mux2_1 _07112_ (.A0(_03472_),
    .A1(_01865_),
    .S(rst),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_1 _07113_ (.A0(_03474_),
    .A1(_01864_),
    .S(rst),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_1 _07114_ (.A0(_03476_),
    .A1(_01863_),
    .S(rst),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _07115_ (.A0(_03478_),
    .A1(_01862_),
    .S(rst),
    .X(_03479_));
 sky130_fd_sc_hd__mux2_1 _07116_ (.A0(_03480_),
    .A1(_01861_),
    .S(rst),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _07117_ (.A0(_03482_),
    .A1(_01860_),
    .S(rst),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _07118_ (.A0(_03484_),
    .A1(_01859_),
    .S(rst),
    .X(_03485_));
 sky130_fd_sc_hd__mux2_1 _07119_ (.A0(_03486_),
    .A1(_01858_),
    .S(rst),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _07120_ (.A0(_03488_),
    .A1(_01857_),
    .S(rst),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _07121_ (.A0(_03490_),
    .A1(_01856_),
    .S(rst),
    .X(_03491_));
 sky130_fd_sc_hd__mux2_1 _07122_ (.A0(_03492_),
    .A1(_01855_),
    .S(rst),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _07123_ (.A0(_03494_),
    .A1(_01854_),
    .S(rst),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _07124_ (.A0(_03496_),
    .A1(_01853_),
    .S(rst),
    .X(_03497_));
 sky130_fd_sc_hd__mux2_1 _07125_ (.A0(_03498_),
    .A1(_01852_),
    .S(rst),
    .X(_03499_));
 sky130_fd_sc_hd__mux2_1 _07126_ (.A0(_03500_),
    .A1(_01851_),
    .S(rst),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _07127_ (.A0(_03502_),
    .A1(_01850_),
    .S(rst),
    .X(_03503_));
 sky130_fd_sc_hd__mux2_1 _07128_ (.A0(_03504_),
    .A1(_01849_),
    .S(rst),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _07129_ (.A0(_03506_),
    .A1(_01848_),
    .S(rst),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _07130_ (.A0(_03508_),
    .A1(_01847_),
    .S(rst),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _07131_ (.A0(_03510_),
    .A1(_01846_),
    .S(rst),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _07132_ (.A0(_03512_),
    .A1(_01845_),
    .S(rst),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _07133_ (.A0(_03514_),
    .A1(_01844_),
    .S(rst),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _07134_ (.A0(_03516_),
    .A1(_01843_),
    .S(rst),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _07135_ (.A0(_03518_),
    .A1(_01842_),
    .S(rst),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _07136_ (.A0(_03520_),
    .A1(_01841_),
    .S(rst),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _07137_ (.A0(_03522_),
    .A1(_01840_),
    .S(rst),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _07138_ (.A0(_03524_),
    .A1(_01839_),
    .S(rst),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_1 _07139_ (.A0(_03526_),
    .A1(_01838_),
    .S(rst),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _07140_ (.A0(_03528_),
    .A1(_01837_),
    .S(rst),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_1 _07141_ (.A0(_03530_),
    .A1(_01836_),
    .S(rst),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_1 _07142_ (.A0(_03532_),
    .A1(_01835_),
    .S(rst),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _07143_ (.A0(_03534_),
    .A1(_01834_),
    .S(rst),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _07144_ (.A0(_03536_),
    .A1(_01833_),
    .S(rst),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _07145_ (.A0(_03538_),
    .A1(_01832_),
    .S(rst),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _07146_ (.A0(_03540_),
    .A1(_01831_),
    .S(rst),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _07147_ (.A0(_03542_),
    .A1(_01830_),
    .S(rst),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _07148_ (.A0(_03544_),
    .A1(_01829_),
    .S(rst),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_1 _07149_ (.A0(_03546_),
    .A1(_01828_),
    .S(rst),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _07150_ (.A0(_03548_),
    .A1(_01827_),
    .S(rst),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _07151_ (.A0(_03550_),
    .A1(_01826_),
    .S(rst),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_1 _07152_ (.A0(_03552_),
    .A1(_01825_),
    .S(rst),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_1 _07153_ (.A0(_03554_),
    .A1(_01824_),
    .S(rst),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _07154_ (.A0(_03556_),
    .A1(_01823_),
    .S(rst),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _07155_ (.A0(_03558_),
    .A1(_01822_),
    .S(rst),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _07156_ (.A0(_03560_),
    .A1(_01542_),
    .S(rst),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _07157_ (.A0(_03562_),
    .A1(_01821_),
    .S(rst),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _07158_ (.A0(_03564_),
    .A1(_01820_),
    .S(rst),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _07159_ (.A0(_03566_),
    .A1(_01819_),
    .S(rst),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _07160_ (.A0(_03568_),
    .A1(_01818_),
    .S(rst),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _07161_ (.A0(_03570_),
    .A1(_01817_),
    .S(rst),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _07162_ (.A0(_03572_),
    .A1(_01816_),
    .S(rst),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _07163_ (.A0(_03574_),
    .A1(_01815_),
    .S(rst),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _07164_ (.A0(_03576_),
    .A1(_01814_),
    .S(rst),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _07165_ (.A0(_03578_),
    .A1(_01813_),
    .S(rst),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(_03580_),
    .A1(_01812_),
    .S(rst),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _07167_ (.A0(_03582_),
    .A1(_01811_),
    .S(rst),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _07168_ (.A0(_03584_),
    .A1(_01810_),
    .S(rst),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _07169_ (.A0(_03586_),
    .A1(_01809_),
    .S(rst),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _07170_ (.A0(_03588_),
    .A1(_01808_),
    .S(rst),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _07171_ (.A0(_03590_),
    .A1(_01807_),
    .S(rst),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _07172_ (.A0(_03592_),
    .A1(_01806_),
    .S(rst),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _07173_ (.A0(_03594_),
    .A1(_01805_),
    .S(rst),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _07174_ (.A0(_03596_),
    .A1(_01804_),
    .S(rst),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _07175_ (.A0(_03598_),
    .A1(_01803_),
    .S(rst),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _07176_ (.A0(_03600_),
    .A1(_01802_),
    .S(rst),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _07177_ (.A0(_03602_),
    .A1(_01801_),
    .S(rst),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _07178_ (.A0(_03604_),
    .A1(_01800_),
    .S(rst),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _07179_ (.A0(_03606_),
    .A1(_01799_),
    .S(rst),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(_03608_),
    .A1(_01798_),
    .S(rst),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _07181_ (.A0(_03610_),
    .A1(_01797_),
    .S(rst),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _07182_ (.A0(_03612_),
    .A1(_01796_),
    .S(rst),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _07183_ (.A0(_03614_),
    .A1(_01795_),
    .S(rst),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _07184_ (.A0(_03616_),
    .A1(_01794_),
    .S(rst),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_1 _07185_ (.A0(_03618_),
    .A1(_01793_),
    .S(rst),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _07186_ (.A0(_03620_),
    .A1(_01792_),
    .S(rst),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_1 _07187_ (.A0(_03622_),
    .A1(_01791_),
    .S(rst),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _07188_ (.A0(_03624_),
    .A1(_01790_),
    .S(rst),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _07189_ (.A0(_03626_),
    .A1(_01789_),
    .S(rst),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _07190_ (.A0(_03628_),
    .A1(_01788_),
    .S(rst),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _07191_ (.A0(_03630_),
    .A1(_01787_),
    .S(rst),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _07192_ (.A0(_03632_),
    .A1(_01786_),
    .S(rst),
    .X(_03633_));
 sky130_fd_sc_hd__mux2_1 _07193_ (.A0(_03634_),
    .A1(_01785_),
    .S(rst),
    .X(_03635_));
 sky130_fd_sc_hd__mux2_1 _07194_ (.A0(_03636_),
    .A1(_01784_),
    .S(rst),
    .X(_03637_));
 sky130_fd_sc_hd__mux2_1 _07195_ (.A0(_03638_),
    .A1(_01783_),
    .S(rst),
    .X(_03639_));
 sky130_fd_sc_hd__mux2_1 _07196_ (.A0(_03640_),
    .A1(_01782_),
    .S(rst),
    .X(_03641_));
 sky130_fd_sc_hd__mux2_1 _07197_ (.A0(_03642_),
    .A1(_01781_),
    .S(rst),
    .X(_03643_));
 sky130_fd_sc_hd__mux2_1 _07198_ (.A0(_03644_),
    .A1(_01780_),
    .S(rst),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _07199_ (.A0(_03646_),
    .A1(_01779_),
    .S(rst),
    .X(_03647_));
 sky130_fd_sc_hd__mux2_1 _07200_ (.A0(_03648_),
    .A1(_01778_),
    .S(rst),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _07201_ (.A0(_03650_),
    .A1(_01777_),
    .S(rst),
    .X(_03651_));
 sky130_fd_sc_hd__mux2_1 _07202_ (.A0(_03652_),
    .A1(_01776_),
    .S(rst),
    .X(_03653_));
 sky130_fd_sc_hd__mux2_1 _07203_ (.A0(_03654_),
    .A1(_01775_),
    .S(rst),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_1 _07204_ (.A0(_03656_),
    .A1(_01774_),
    .S(rst),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _07205_ (.A0(_03658_),
    .A1(_01773_),
    .S(rst),
    .X(_03659_));
 sky130_fd_sc_hd__mux2_1 _07206_ (.A0(_03660_),
    .A1(_01772_),
    .S(rst),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_1 _07207_ (.A0(_03662_),
    .A1(_01770_),
    .S(rst),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _07208_ (.A0(_03664_),
    .A1(_01769_),
    .S(rst),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _07209_ (.A0(_03666_),
    .A1(_01768_),
    .S(rst),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _07210_ (.A0(_03668_),
    .A1(_01767_),
    .S(rst),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _07211_ (.A0(_03670_),
    .A1(_01766_),
    .S(rst),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _07212_ (.A0(_03672_),
    .A1(_01765_),
    .S(rst),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _07213_ (.A0(_03674_),
    .A1(_01764_),
    .S(rst),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _07214_ (.A0(_03676_),
    .A1(_01763_),
    .S(rst),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _07215_ (.A0(_03678_),
    .A1(_01762_),
    .S(rst),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _07216_ (.A0(_03680_),
    .A1(_01761_),
    .S(rst),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _07217_ (.A0(_03682_),
    .A1(_01760_),
    .S(rst),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _07218_ (.A0(_03684_),
    .A1(_01759_),
    .S(rst),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _07219_ (.A0(_03686_),
    .A1(_01758_),
    .S(rst),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _07220_ (.A0(_03688_),
    .A1(_01757_),
    .S(rst),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _07221_ (.A0(_03690_),
    .A1(_01756_),
    .S(rst),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _07222_ (.A0(_03692_),
    .A1(_01755_),
    .S(rst),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _07223_ (.A0(_03694_),
    .A1(_01754_),
    .S(rst),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _07224_ (.A0(_03696_),
    .A1(_01753_),
    .S(rst),
    .X(_03697_));
 sky130_fd_sc_hd__mux2_1 _07225_ (.A0(_03698_),
    .A1(_01752_),
    .S(rst),
    .X(_03699_));
 sky130_fd_sc_hd__mux2_1 _07226_ (.A0(_03700_),
    .A1(_01751_),
    .S(rst),
    .X(_03701_));
 sky130_fd_sc_hd__mux2_1 _07227_ (.A0(_03702_),
    .A1(_01750_),
    .S(rst),
    .X(_03703_));
 sky130_fd_sc_hd__mux2_1 _07228_ (.A0(_03704_),
    .A1(_01749_),
    .S(rst),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _07229_ (.A0(_03706_),
    .A1(_01748_),
    .S(rst),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _07230_ (.A0(_03708_),
    .A1(_01747_),
    .S(rst),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _07231_ (.A0(_03710_),
    .A1(_01746_),
    .S(rst),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _07232_ (.A0(_03712_),
    .A1(_01745_),
    .S(rst),
    .X(_03713_));
 sky130_fd_sc_hd__mux2_1 _07233_ (.A0(_03714_),
    .A1(_01744_),
    .S(rst),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _07234_ (.A0(_03716_),
    .A1(_01743_),
    .S(rst),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _07235_ (.A0(_03718_),
    .A1(_01742_),
    .S(rst),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _07236_ (.A0(_03720_),
    .A1(_01741_),
    .S(rst),
    .X(_03721_));
 sky130_fd_sc_hd__mux2_1 _07237_ (.A0(_03722_),
    .A1(_01740_),
    .S(rst),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _07238_ (.A0(_03724_),
    .A1(_01739_),
    .S(rst),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_1 _07239_ (.A0(_03726_),
    .A1(_01738_),
    .S(rst),
    .X(_03727_));
 sky130_fd_sc_hd__mux2_1 _07240_ (.A0(_03728_),
    .A1(_01737_),
    .S(rst),
    .X(_03729_));
 sky130_fd_sc_hd__mux2_1 _07241_ (.A0(_03730_),
    .A1(_01736_),
    .S(rst),
    .X(_03731_));
 sky130_fd_sc_hd__mux2_1 _07242_ (.A0(_03732_),
    .A1(_01735_),
    .S(rst),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_1 _07243_ (.A0(_03734_),
    .A1(_01734_),
    .S(rst),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _07244_ (.A0(_03736_),
    .A1(_01733_),
    .S(rst),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _07245_ (.A0(_03738_),
    .A1(_01732_),
    .S(rst),
    .X(_03739_));
 sky130_fd_sc_hd__mux2_1 _07246_ (.A0(_03740_),
    .A1(_01731_),
    .S(rst),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _07247_ (.A0(_03742_),
    .A1(_01730_),
    .S(rst),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _07248_ (.A0(_03744_),
    .A1(_01729_),
    .S(rst),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _07249_ (.A0(_03746_),
    .A1(_01728_),
    .S(rst),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _07250_ (.A0(_03748_),
    .A1(_01727_),
    .S(rst),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_1 _07251_ (.A0(_03750_),
    .A1(_01726_),
    .S(rst),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _07252_ (.A0(_03752_),
    .A1(_01725_),
    .S(rst),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _07253_ (.A0(_03754_),
    .A1(_01724_),
    .S(rst),
    .X(_03755_));
 sky130_fd_sc_hd__mux2_1 _07254_ (.A0(_03756_),
    .A1(_01723_),
    .S(rst),
    .X(_03757_));
 sky130_fd_sc_hd__mux2_1 _07255_ (.A0(_03758_),
    .A1(_01722_),
    .S(rst),
    .X(_03759_));
 sky130_fd_sc_hd__mux2_1 _07256_ (.A0(_03760_),
    .A1(_01721_),
    .S(rst),
    .X(_03761_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(_03762_),
    .A1(_01720_),
    .S(rst),
    .X(_03763_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(_03764_),
    .A1(_01719_),
    .S(rst),
    .X(_03765_));
 sky130_fd_sc_hd__mux2_1 _07259_ (.A0(_03766_),
    .A1(_01718_),
    .S(rst),
    .X(_03767_));
 sky130_fd_sc_hd__mux2_1 _07260_ (.A0(_03768_),
    .A1(_01717_),
    .S(rst),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _07261_ (.A0(_03770_),
    .A1(_01716_),
    .S(rst),
    .X(_03771_));
 sky130_fd_sc_hd__mux2_1 _07262_ (.A0(_03772_),
    .A1(_01715_),
    .S(rst),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _07263_ (.A0(_03774_),
    .A1(_01714_),
    .S(rst),
    .X(_03775_));
 sky130_fd_sc_hd__mux2_1 _07264_ (.A0(_03776_),
    .A1(_01713_),
    .S(rst),
    .X(_03777_));
 sky130_fd_sc_hd__mux2_1 _07265_ (.A0(_03778_),
    .A1(_01712_),
    .S(rst),
    .X(_03779_));
 sky130_fd_sc_hd__mux2_1 _07266_ (.A0(_03780_),
    .A1(_01711_),
    .S(rst),
    .X(_03781_));
 sky130_fd_sc_hd__mux2_1 _07267_ (.A0(_03782_),
    .A1(_01710_),
    .S(rst),
    .X(_03783_));
 sky130_fd_sc_hd__mux2_1 _07268_ (.A0(_03784_),
    .A1(_01709_),
    .S(rst),
    .X(_03785_));
 sky130_fd_sc_hd__mux2_1 _07269_ (.A0(_03786_),
    .A1(_01708_),
    .S(rst),
    .X(_03787_));
 sky130_fd_sc_hd__mux2_1 _07270_ (.A0(_03788_),
    .A1(_01707_),
    .S(rst),
    .X(_03789_));
 sky130_fd_sc_hd__mux2_1 _07271_ (.A0(_03790_),
    .A1(_01706_),
    .S(rst),
    .X(_03791_));
 sky130_fd_sc_hd__mux2_1 _07272_ (.A0(_03792_),
    .A1(_01705_),
    .S(rst),
    .X(_03793_));
 sky130_fd_sc_hd__mux2_1 _07273_ (.A0(_03794_),
    .A1(_01704_),
    .S(rst),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _07274_ (.A0(_03796_),
    .A1(_01703_),
    .S(rst),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_1 _07275_ (.A0(_03798_),
    .A1(_01702_),
    .S(rst),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _07276_ (.A0(_03800_),
    .A1(_01701_),
    .S(rst),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _07277_ (.A0(_03802_),
    .A1(_01700_),
    .S(rst),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_1 _07278_ (.A0(_03804_),
    .A1(_01699_),
    .S(rst),
    .X(_03805_));
 sky130_fd_sc_hd__mux2_1 _07279_ (.A0(_03806_),
    .A1(_01698_),
    .S(rst),
    .X(_03807_));
 sky130_fd_sc_hd__mux2_1 _07280_ (.A0(_03808_),
    .A1(_01697_),
    .S(rst),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_1 _07281_ (.A0(_03810_),
    .A1(_01696_),
    .S(rst),
    .X(_03811_));
 sky130_fd_sc_hd__mux2_1 _07282_ (.A0(_03812_),
    .A1(_01695_),
    .S(rst),
    .X(_03813_));
 sky130_fd_sc_hd__mux2_1 _07283_ (.A0(_03814_),
    .A1(_01694_),
    .S(rst),
    .X(_03815_));
 sky130_fd_sc_hd__mux2_1 _07284_ (.A0(_03816_),
    .A1(_01693_),
    .S(rst),
    .X(_03817_));
 sky130_fd_sc_hd__mux2_1 _07285_ (.A0(_03818_),
    .A1(_01692_),
    .S(rst),
    .X(_03819_));
 sky130_fd_sc_hd__mux2_1 _07286_ (.A0(_03820_),
    .A1(_01691_),
    .S(rst),
    .X(_03821_));
 sky130_fd_sc_hd__mux2_1 _07287_ (.A0(_03822_),
    .A1(_01690_),
    .S(rst),
    .X(_03823_));
 sky130_fd_sc_hd__mux2_1 _07288_ (.A0(_03824_),
    .A1(_01689_),
    .S(rst),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_1 _07289_ (.A0(_03826_),
    .A1(_01688_),
    .S(rst),
    .X(_03827_));
 sky130_fd_sc_hd__mux2_1 _07290_ (.A0(_03828_),
    .A1(_01687_),
    .S(rst),
    .X(_03829_));
 sky130_fd_sc_hd__mux2_1 _07291_ (.A0(_03830_),
    .A1(_01686_),
    .S(rst),
    .X(_03831_));
 sky130_fd_sc_hd__mux2_1 _07292_ (.A0(_03832_),
    .A1(_01685_),
    .S(rst),
    .X(_03833_));
 sky130_fd_sc_hd__mux2_1 _07293_ (.A0(_03834_),
    .A1(_01684_),
    .S(rst),
    .X(_03835_));
 sky130_fd_sc_hd__mux2_1 _07294_ (.A0(_03836_),
    .A1(_01683_),
    .S(rst),
    .X(_03837_));
 sky130_fd_sc_hd__mux2_1 _07295_ (.A0(_03838_),
    .A1(_01682_),
    .S(rst),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(_03840_),
    .A1(_01681_),
    .S(rst),
    .X(_03841_));
 sky130_fd_sc_hd__mux2_1 _07297_ (.A0(_03842_),
    .A1(_01680_),
    .S(rst),
    .X(_03843_));
 sky130_fd_sc_hd__mux2_1 _07298_ (.A0(_03844_),
    .A1(_01679_),
    .S(rst),
    .X(_03845_));
 sky130_fd_sc_hd__mux2_1 _07299_ (.A0(_03846_),
    .A1(_01678_),
    .S(rst),
    .X(_03847_));
 sky130_fd_sc_hd__mux2_1 _07300_ (.A0(_03848_),
    .A1(_01677_),
    .S(rst),
    .X(_03849_));
 sky130_fd_sc_hd__mux2_1 _07301_ (.A0(_03850_),
    .A1(_01676_),
    .S(rst),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_1 _07302_ (.A0(_03852_),
    .A1(_01675_),
    .S(rst),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _07303_ (.A0(_03854_),
    .A1(_01674_),
    .S(rst),
    .X(_03855_));
 sky130_fd_sc_hd__mux2_1 _07304_ (.A0(_03856_),
    .A1(_01673_),
    .S(rst),
    .X(_03857_));
 sky130_fd_sc_hd__mux2_1 _07305_ (.A0(_03858_),
    .A1(_01672_),
    .S(rst),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_1 _07306_ (.A0(_03860_),
    .A1(_01671_),
    .S(rst),
    .X(_03861_));
 sky130_fd_sc_hd__mux2_1 _07307_ (.A0(_03862_),
    .A1(_01670_),
    .S(rst),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _07308_ (.A0(_03864_),
    .A1(_01669_),
    .S(rst),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _07309_ (.A0(_03866_),
    .A1(_01668_),
    .S(rst),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _07310_ (.A0(_03868_),
    .A1(_01667_),
    .S(rst),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_1 _07311_ (.A0(_03870_),
    .A1(_01666_),
    .S(rst),
    .X(_03871_));
 sky130_fd_sc_hd__mux2_1 _07312_ (.A0(_03872_),
    .A1(_01665_),
    .S(rst),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _07313_ (.A0(_03874_),
    .A1(_01664_),
    .S(rst),
    .X(_03875_));
 sky130_fd_sc_hd__mux2_1 _07314_ (.A0(_03876_),
    .A1(_01663_),
    .S(rst),
    .X(_03877_));
 sky130_fd_sc_hd__mux2_1 _07315_ (.A0(_03878_),
    .A1(_01662_),
    .S(rst),
    .X(_03879_));
 sky130_fd_sc_hd__mux2_1 _07316_ (.A0(_03880_),
    .A1(_01661_),
    .S(rst),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_1 _07317_ (.A0(_03882_),
    .A1(_01660_),
    .S(rst),
    .X(_03883_));
 sky130_fd_sc_hd__mux2_1 _07318_ (.A0(_03884_),
    .A1(_01659_),
    .S(rst),
    .X(_03885_));
 sky130_fd_sc_hd__mux2_1 _07319_ (.A0(_03886_),
    .A1(_01658_),
    .S(rst),
    .X(_03887_));
 sky130_fd_sc_hd__mux2_1 _07320_ (.A0(_03888_),
    .A1(_01657_),
    .S(rst),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _07321_ (.A0(_03890_),
    .A1(_01656_),
    .S(rst),
    .X(_03891_));
 sky130_fd_sc_hd__mux2_1 _07322_ (.A0(_03892_),
    .A1(_01655_),
    .S(rst),
    .X(_03893_));
 sky130_fd_sc_hd__mux2_1 _07323_ (.A0(_03894_),
    .A1(_01654_),
    .S(rst),
    .X(_03895_));
 sky130_fd_sc_hd__mux2_1 _07324_ (.A0(_03896_),
    .A1(_01653_),
    .S(rst),
    .X(_03897_));
 sky130_fd_sc_hd__mux2_1 _07325_ (.A0(_03898_),
    .A1(_01652_),
    .S(rst),
    .X(_03899_));
 sky130_fd_sc_hd__mux2_1 _07326_ (.A0(_03900_),
    .A1(_01651_),
    .S(rst),
    .X(_03901_));
 sky130_fd_sc_hd__mux2_1 _07327_ (.A0(_03902_),
    .A1(_01650_),
    .S(rst),
    .X(_03903_));
 sky130_fd_sc_hd__mux2_1 _07328_ (.A0(_03904_),
    .A1(_01649_),
    .S(rst),
    .X(_03905_));
 sky130_fd_sc_hd__mux2_1 _07329_ (.A0(_03906_),
    .A1(_01648_),
    .S(rst),
    .X(_03907_));
 sky130_fd_sc_hd__mux2_1 _07330_ (.A0(_03908_),
    .A1(_01647_),
    .S(rst),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _07331_ (.A0(_03910_),
    .A1(_01646_),
    .S(rst),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _07332_ (.A0(_03912_),
    .A1(_01645_),
    .S(rst),
    .X(_03913_));
 sky130_fd_sc_hd__mux2_1 _07333_ (.A0(_03914_),
    .A1(_01644_),
    .S(rst),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _07334_ (.A0(_03916_),
    .A1(_01643_),
    .S(rst),
    .X(_03917_));
 sky130_fd_sc_hd__mux2_1 _07335_ (.A0(_03918_),
    .A1(_01642_),
    .S(rst),
    .X(_03919_));
 sky130_fd_sc_hd__mux2_1 _07336_ (.A0(_03920_),
    .A1(_01641_),
    .S(rst),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _07337_ (.A0(_03922_),
    .A1(_01640_),
    .S(rst),
    .X(_03923_));
 sky130_fd_sc_hd__mux2_1 _07338_ (.A0(_03924_),
    .A1(_01639_),
    .S(rst),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _07339_ (.A0(_03926_),
    .A1(_01638_),
    .S(rst),
    .X(_03927_));
 sky130_fd_sc_hd__mux2_1 _07340_ (.A0(_03928_),
    .A1(_01637_),
    .S(rst),
    .X(_03929_));
 sky130_fd_sc_hd__mux2_1 _07341_ (.A0(_03930_),
    .A1(_01636_),
    .S(rst),
    .X(_03931_));
 sky130_fd_sc_hd__mux2_1 _07342_ (.A0(_03932_),
    .A1(_01635_),
    .S(rst),
    .X(_03933_));
 sky130_fd_sc_hd__mux2_1 _07343_ (.A0(_03934_),
    .A1(_01634_),
    .S(rst),
    .X(_03935_));
 sky130_fd_sc_hd__mux2_1 _07344_ (.A0(_03936_),
    .A1(_01633_),
    .S(rst),
    .X(_03937_));
 sky130_fd_sc_hd__mux2_1 _07345_ (.A0(_03938_),
    .A1(_01632_),
    .S(rst),
    .X(_03939_));
 sky130_fd_sc_hd__mux2_1 _07346_ (.A0(_03940_),
    .A1(_01631_),
    .S(rst),
    .X(_03941_));
 sky130_fd_sc_hd__mux2_1 _07347_ (.A0(_03942_),
    .A1(_01630_),
    .S(rst),
    .X(_03943_));
 sky130_fd_sc_hd__mux2_1 _07348_ (.A0(_03944_),
    .A1(_01629_),
    .S(rst),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _07349_ (.A0(_03946_),
    .A1(_01628_),
    .S(rst),
    .X(_03947_));
 sky130_fd_sc_hd__mux2_1 _07350_ (.A0(_03948_),
    .A1(_01627_),
    .S(rst),
    .X(_03949_));
 sky130_fd_sc_hd__mux2_1 _07351_ (.A0(_03950_),
    .A1(_01626_),
    .S(rst),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_1 _07352_ (.A0(_03952_),
    .A1(_01625_),
    .S(rst),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _07353_ (.A0(_03954_),
    .A1(_01624_),
    .S(rst),
    .X(_03955_));
 sky130_fd_sc_hd__mux2_1 _07354_ (.A0(_03956_),
    .A1(_01623_),
    .S(rst),
    .X(_03957_));
 sky130_fd_sc_hd__mux2_1 _07355_ (.A0(_03958_),
    .A1(_01622_),
    .S(rst),
    .X(_03959_));
 sky130_fd_sc_hd__mux2_1 _07356_ (.A0(_03960_),
    .A1(_01621_),
    .S(rst),
    .X(_03961_));
 sky130_fd_sc_hd__mux2_1 _07357_ (.A0(_03962_),
    .A1(_01620_),
    .S(rst),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_1 _07358_ (.A0(_03964_),
    .A1(_01619_),
    .S(rst),
    .X(_03965_));
 sky130_fd_sc_hd__mux2_1 _07359_ (.A0(_03966_),
    .A1(_01618_),
    .S(rst),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _07360_ (.A0(_03968_),
    .A1(_01617_),
    .S(rst),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_1 _07361_ (.A0(_03970_),
    .A1(_01771_),
    .S(rst),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_1 _07362_ (.A0(_03972_),
    .A1(_01616_),
    .S(rst),
    .X(_03973_));
 sky130_fd_sc_hd__mux2_1 _07363_ (.A0(_03974_),
    .A1(_01615_),
    .S(rst),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _07364_ (.A0(_03976_),
    .A1(_01614_),
    .S(rst),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _07365_ (.A0(_03978_),
    .A1(_01613_),
    .S(rst),
    .X(_03979_));
 sky130_fd_sc_hd__mux2_1 _07366_ (.A0(_03980_),
    .A1(_01612_),
    .S(rst),
    .X(_03981_));
 sky130_fd_sc_hd__mux2_1 _07367_ (.A0(_03982_),
    .A1(_01611_),
    .S(rst),
    .X(_03983_));
 sky130_fd_sc_hd__mux2_1 _07368_ (.A0(_03984_),
    .A1(_01610_),
    .S(rst),
    .X(_03985_));
 sky130_fd_sc_hd__mux2_1 _07369_ (.A0(_03986_),
    .A1(_01609_),
    .S(rst),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _07370_ (.A0(_03988_),
    .A1(_01608_),
    .S(rst),
    .X(_03989_));
 sky130_fd_sc_hd__mux2_1 _07371_ (.A0(_03990_),
    .A1(_01607_),
    .S(rst),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _07372_ (.A0(_03992_),
    .A1(_01606_),
    .S(rst),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _07373_ (.A0(_03994_),
    .A1(_01605_),
    .S(rst),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _07374_ (.A0(_03996_),
    .A1(_01604_),
    .S(rst),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _07375_ (.A0(_03998_),
    .A1(_01603_),
    .S(rst),
    .X(_03999_));
 sky130_fd_sc_hd__mux2_1 _07376_ (.A0(_04000_),
    .A1(_01602_),
    .S(rst),
    .X(_04001_));
 sky130_fd_sc_hd__mux2_1 _07377_ (.A0(_04002_),
    .A1(_01601_),
    .S(rst),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _07378_ (.A0(_04004_),
    .A1(_01600_),
    .S(rst),
    .X(_04005_));
 sky130_fd_sc_hd__mux2_1 _07379_ (.A0(_04006_),
    .A1(_01599_),
    .S(rst),
    .X(_04007_));
 sky130_fd_sc_hd__mux2_1 _07380_ (.A0(_04008_),
    .A1(_01598_),
    .S(rst),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_1 _07381_ (.A0(_04010_),
    .A1(_01597_),
    .S(rst),
    .X(_04011_));
 sky130_fd_sc_hd__mux2_1 _07382_ (.A0(_04012_),
    .A1(_01596_),
    .S(rst),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_1 _07383_ (.A0(_04014_),
    .A1(_01595_),
    .S(rst),
    .X(_04015_));
 sky130_fd_sc_hd__mux2_1 _07384_ (.A0(_04016_),
    .A1(_01594_),
    .S(rst),
    .X(_04017_));
 sky130_fd_sc_hd__mux2_1 _07385_ (.A0(_04018_),
    .A1(_01593_),
    .S(rst),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _07386_ (.A0(_04020_),
    .A1(_01592_),
    .S(rst),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _07387_ (.A0(_04022_),
    .A1(_01591_),
    .S(rst),
    .X(_04023_));
 sky130_fd_sc_hd__mux2_1 _07388_ (.A0(_04024_),
    .A1(_01590_),
    .S(rst),
    .X(_04025_));
 sky130_fd_sc_hd__mux2_1 _07389_ (.A0(_04026_),
    .A1(_01589_),
    .S(rst),
    .X(_04027_));
 sky130_fd_sc_hd__mux2_1 _07390_ (.A0(_04028_),
    .A1(_01550_),
    .S(rst),
    .X(_04029_));
 sky130_fd_sc_hd__mux2_1 _07391_ (.A0(_04030_),
    .A1(_01549_),
    .S(rst),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_1 _07392_ (.A0(_04032_),
    .A1(_01588_),
    .S(rst),
    .X(_04033_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(_04034_),
    .A1(_01551_),
    .S(rst),
    .X(_04035_));
 sky130_fd_sc_hd__mux2_1 _07394_ (.A0(_04036_),
    .A1(_01548_),
    .S(rst),
    .X(_04037_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(_04038_),
    .A1(_01587_),
    .S(rst),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_1 _07396_ (.A0(_04040_),
    .A1(_01552_),
    .S(rst),
    .X(_04041_));
 sky130_fd_sc_hd__mux2_1 _07397_ (.A0(_04042_),
    .A1(_01546_),
    .S(rst),
    .X(_04043_));
 sky130_fd_sc_hd__mux2_1 _07398_ (.A0(_04044_),
    .A1(_01586_),
    .S(rst),
    .X(_04045_));
 sky130_fd_sc_hd__mux2_1 _07399_ (.A0(_04046_),
    .A1(_01543_),
    .S(rst),
    .X(_04047_));
 sky130_fd_sc_hd__mux2_1 _07400_ (.A0(_04048_),
    .A1(_01585_),
    .S(rst),
    .X(_04049_));
 sky130_fd_sc_hd__mux2_1 _07401_ (.A0(_04050_),
    .A1(_01553_),
    .S(rst),
    .X(_04051_));
 sky130_fd_sc_hd__mux2_1 _07402_ (.A0(_04052_),
    .A1(_01545_),
    .S(rst),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_1 _07403_ (.A0(_04054_),
    .A1(_01584_),
    .S(rst),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _07404_ (.A0(_04056_),
    .A1(_01583_),
    .S(rst),
    .X(_04057_));
 sky130_fd_sc_hd__mux2_1 _07405_ (.A0(_04058_),
    .A1(_01582_),
    .S(rst),
    .X(_04059_));
 sky130_fd_sc_hd__mux2_1 _07406_ (.A0(_04060_),
    .A1(_01581_),
    .S(rst),
    .X(_04061_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(_04062_),
    .A1(_01580_),
    .S(rst),
    .X(_04063_));
 sky130_fd_sc_hd__mux2_1 _07408_ (.A0(_04064_),
    .A1(_01579_),
    .S(rst),
    .X(_04065_));
 sky130_fd_sc_hd__mux2_1 _07409_ (.A0(_04066_),
    .A1(_01578_),
    .S(rst),
    .X(_04067_));
 sky130_fd_sc_hd__mux2_1 _07410_ (.A0(_04068_),
    .A1(_01577_),
    .S(rst),
    .X(_04069_));
 sky130_fd_sc_hd__mux2_1 _07411_ (.A0(_04070_),
    .A1(_01576_),
    .S(rst),
    .X(_04071_));
 sky130_fd_sc_hd__mux2_1 _07412_ (.A0(_04072_),
    .A1(_01575_),
    .S(rst),
    .X(_04073_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(_04074_),
    .A1(_01574_),
    .S(rst),
    .X(_04075_));
 sky130_fd_sc_hd__mux2_1 _07414_ (.A0(_04076_),
    .A1(_01573_),
    .S(rst),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_1 _07415_ (.A0(_04078_),
    .A1(_01572_),
    .S(rst),
    .X(_04079_));
 sky130_fd_sc_hd__mux2_1 _07416_ (.A0(_04080_),
    .A1(_01571_),
    .S(rst),
    .X(_04081_));
 sky130_fd_sc_hd__mux2_1 _07417_ (.A0(_04082_),
    .A1(_01570_),
    .S(rst),
    .X(_04083_));
 sky130_fd_sc_hd__mux2_1 _07418_ (.A0(_04084_),
    .A1(_01569_),
    .S(rst),
    .X(_04085_));
 sky130_fd_sc_hd__mux2_1 _07419_ (.A0(_04086_),
    .A1(_01568_),
    .S(rst),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _07420_ (.A0(_04088_),
    .A1(_01567_),
    .S(rst),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _07421_ (.A0(_04090_),
    .A1(_01566_),
    .S(rst),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _07422_ (.A0(_04092_),
    .A1(_01565_),
    .S(rst),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _07423_ (.A0(_04094_),
    .A1(_01564_),
    .S(rst),
    .X(_04095_));
 sky130_fd_sc_hd__mux2_1 _07424_ (.A0(_04096_),
    .A1(_01563_),
    .S(rst),
    .X(_04097_));
 sky130_fd_sc_hd__mux2_1 _07425_ (.A0(_04098_),
    .A1(_01562_),
    .S(rst),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _07426_ (.A0(_04100_),
    .A1(_01561_),
    .S(rst),
    .X(_04101_));
 sky130_fd_sc_hd__mux2_1 _07427_ (.A0(_04102_),
    .A1(_01560_),
    .S(rst),
    .X(_04103_));
 sky130_fd_sc_hd__mux2_1 _07428_ (.A0(_04104_),
    .A1(_01559_),
    .S(rst),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _07429_ (.A0(_04106_),
    .A1(_01558_),
    .S(rst),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _07430_ (.A0(_04108_),
    .A1(_01557_),
    .S(rst),
    .X(_04109_));
 sky130_fd_sc_hd__mux2_1 _07431_ (.A0(_04110_),
    .A1(_01556_),
    .S(rst),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _07432_ (.A0(_04112_),
    .A1(_01555_),
    .S(rst),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_1 _07433_ (.A0(_04114_),
    .A1(_01554_),
    .S(rst),
    .X(_04115_));
 sky130_fd_sc_hd__mux2_1 _07434_ (.A0(_04116_),
    .A1(_01547_),
    .S(rst),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _07435_ (.A0(_04118_),
    .A1(_01544_),
    .S(rst),
    .X(_04119_));
 sky130_fd_sc_hd__conb_1 _07436_ (.LO(_00982_));
 sky130_fd_sc_hd__conb_1 _07437_ (.LO(_00983_));
 sky130_fd_sc_hd__conb_1 _07438_ (.LO(_00984_));
 sky130_fd_sc_hd__conb_1 _07439_ (.LO(_00985_));
 sky130_fd_sc_hd__conb_1 _07440_ (.LO(_00986_));
 sky130_fd_sc_hd__conb_1 _07441_ (.LO(_00987_));
 sky130_fd_sc_hd__conb_1 _07442_ (.LO(_00988_));
 sky130_fd_sc_hd__conb_1 _07443_ (.LO(_00989_));
 sky130_fd_sc_hd__conb_1 _07444_ (.LO(_00990_));
 sky130_fd_sc_hd__conb_1 _07445_ (.LO(_00991_));
 sky130_fd_sc_hd__conb_1 _07446_ (.LO(_00992_));
 sky130_fd_sc_hd__conb_1 _07447_ (.LO(_00993_));
 sky130_fd_sc_hd__conb_1 _07448_ (.LO(_00994_));
 sky130_fd_sc_hd__conb_1 _07449_ (.LO(_00995_));
 sky130_fd_sc_hd__conb_1 _07450_ (.LO(_00996_));
 sky130_fd_sc_hd__conb_1 _07451_ (.LO(_00997_));
 sky130_fd_sc_hd__conb_1 _07452_ (.LO(_00998_));
 sky130_fd_sc_hd__conb_1 _07453_ (.LO(_00999_));
 sky130_fd_sc_hd__conb_1 _07454_ (.LO(_01000_));
 sky130_fd_sc_hd__conb_1 _07455_ (.LO(_01001_));
 sky130_fd_sc_hd__conb_1 _07456_ (.LO(_01002_));
 sky130_fd_sc_hd__conb_1 _07457_ (.LO(_01003_));
 sky130_fd_sc_hd__conb_1 _07458_ (.LO(_01004_));
 sky130_fd_sc_hd__conb_1 _07459_ (.LO(_01005_));
 sky130_fd_sc_hd__conb_1 _07460_ (.LO(_01006_));
 sky130_fd_sc_hd__conb_1 _07461_ (.LO(_01007_));
 sky130_fd_sc_hd__conb_1 _07462_ (.LO(_01008_));
 sky130_fd_sc_hd__conb_1 _07463_ (.LO(_01009_));
 sky130_fd_sc_hd__conb_1 _07464_ (.LO(_01010_));
 sky130_fd_sc_hd__conb_1 _07465_ (.LO(_01011_));
 sky130_fd_sc_hd__conb_1 _07466_ (.LO(_01012_));
 sky130_fd_sc_hd__conb_1 _07467_ (.LO(_01013_));
 sky130_fd_sc_hd__conb_1 _07468_ (.LO(_01014_));
 sky130_fd_sc_hd__conb_1 _07469_ (.LO(_01015_));
 sky130_fd_sc_hd__conb_1 _07470_ (.LO(_01016_));
 sky130_fd_sc_hd__conb_1 _07471_ (.LO(_01017_));
 sky130_fd_sc_hd__conb_1 _07472_ (.LO(_01018_));
 sky130_fd_sc_hd__conb_1 _07473_ (.LO(_01019_));
 sky130_fd_sc_hd__conb_1 _07474_ (.LO(_01020_));
 sky130_fd_sc_hd__conb_1 _07475_ (.LO(_01021_));
 sky130_fd_sc_hd__conb_1 _07476_ (.LO(_01022_));
 sky130_fd_sc_hd__conb_1 _07477_ (.LO(_01023_));
 sky130_fd_sc_hd__conb_1 _07478_ (.LO(_01024_));
 sky130_fd_sc_hd__conb_1 _07479_ (.LO(_01025_));
 sky130_fd_sc_hd__conb_1 _07480_ (.LO(_01026_));
 sky130_fd_sc_hd__conb_1 _07481_ (.LO(_01027_));
 sky130_fd_sc_hd__conb_1 _07482_ (.LO(_01028_));
 sky130_fd_sc_hd__conb_1 _07483_ (.LO(_01029_));
 sky130_fd_sc_hd__conb_1 _07484_ (.LO(_01030_));
 sky130_fd_sc_hd__conb_1 _07485_ (.LO(_01031_));
 sky130_fd_sc_hd__conb_1 _07486_ (.LO(_01032_));
 sky130_fd_sc_hd__conb_1 _07487_ (.LO(_01033_));
 sky130_fd_sc_hd__conb_1 _07488_ (.LO(_01034_));
 sky130_fd_sc_hd__conb_1 _07489_ (.LO(_01035_));
 sky130_fd_sc_hd__conb_1 _07490_ (.LO(_01036_));
 sky130_fd_sc_hd__conb_1 _07491_ (.LO(_01037_));
 sky130_fd_sc_hd__conb_1 _07492_ (.LO(_01038_));
 sky130_fd_sc_hd__conb_1 _07493_ (.LO(_01039_));
 sky130_fd_sc_hd__conb_1 _07494_ (.LO(_01040_));
 sky130_fd_sc_hd__conb_1 _07495_ (.LO(_01041_));
 sky130_fd_sc_hd__conb_1 _07496_ (.LO(_01042_));
 sky130_fd_sc_hd__conb_1 _07497_ (.LO(_01043_));
 sky130_fd_sc_hd__conb_1 _07498_ (.LO(_01044_));
 sky130_fd_sc_hd__conb_1 _07499_ (.LO(_01045_));
 sky130_fd_sc_hd__conb_1 _07500_ (.LO(_01046_));
 sky130_fd_sc_hd__conb_1 _07501_ (.LO(_01047_));
 sky130_fd_sc_hd__conb_1 _07502_ (.LO(_01048_));
 sky130_fd_sc_hd__conb_1 _07503_ (.LO(_01049_));
 sky130_fd_sc_hd__conb_1 _07504_ (.LO(_01050_));
 sky130_fd_sc_hd__conb_1 _07505_ (.LO(_01051_));
 sky130_fd_sc_hd__conb_1 _07506_ (.LO(_01052_));
 sky130_fd_sc_hd__conb_1 _07507_ (.LO(_01053_));
 sky130_fd_sc_hd__conb_1 _07508_ (.LO(_01054_));
 sky130_fd_sc_hd__conb_1 _07509_ (.LO(_01055_));
 sky130_fd_sc_hd__conb_1 _07510_ (.LO(_01056_));
 sky130_fd_sc_hd__conb_1 _07511_ (.LO(_01057_));
 sky130_fd_sc_hd__conb_1 _07512_ (.LO(_01058_));
 sky130_fd_sc_hd__conb_1 _07513_ (.LO(_01059_));
 sky130_fd_sc_hd__conb_1 _07514_ (.LO(_01060_));
 sky130_fd_sc_hd__conb_1 _07515_ (.LO(_01061_));
 sky130_fd_sc_hd__conb_1 _07516_ (.LO(_01062_));
 sky130_fd_sc_hd__conb_1 _07517_ (.LO(_01063_));
 sky130_fd_sc_hd__conb_1 _07518_ (.LO(_01064_));
 sky130_fd_sc_hd__conb_1 _07519_ (.LO(_01065_));
 sky130_fd_sc_hd__conb_1 _07520_ (.LO(_01066_));
 sky130_fd_sc_hd__conb_1 _07521_ (.LO(_01067_));
 sky130_fd_sc_hd__conb_1 _07522_ (.LO(_01068_));
 sky130_fd_sc_hd__conb_1 _07523_ (.LO(_01069_));
 sky130_fd_sc_hd__conb_1 _07524_ (.LO(_01070_));
 sky130_fd_sc_hd__conb_1 _07525_ (.LO(_01071_));
 sky130_fd_sc_hd__conb_1 _07526_ (.LO(_01072_));
 sky130_fd_sc_hd__conb_1 _07527_ (.LO(_01073_));
 sky130_fd_sc_hd__conb_1 _07528_ (.LO(_01074_));
 sky130_fd_sc_hd__conb_1 _07529_ (.LO(_01075_));
 sky130_fd_sc_hd__conb_1 _07530_ (.LO(_01076_));
 sky130_fd_sc_hd__conb_1 _07531_ (.LO(_01077_));
 sky130_fd_sc_hd__conb_1 _07532_ (.LO(_01078_));
 sky130_fd_sc_hd__conb_1 _07533_ (.LO(_01079_));
 sky130_fd_sc_hd__conb_1 _07534_ (.LO(_01080_));
 sky130_fd_sc_hd__conb_1 _07535_ (.LO(_01081_));
 sky130_fd_sc_hd__conb_1 _07536_ (.LO(_01082_));
 sky130_fd_sc_hd__conb_1 _07537_ (.LO(_01083_));
 sky130_fd_sc_hd__conb_1 _07538_ (.LO(_01084_));
 sky130_fd_sc_hd__conb_1 _07539_ (.LO(_01085_));
 sky130_fd_sc_hd__conb_1 _07540_ (.LO(_01086_));
 sky130_fd_sc_hd__conb_1 _07541_ (.LO(_01087_));
 sky130_fd_sc_hd__conb_1 _07542_ (.LO(_01088_));
 sky130_fd_sc_hd__conb_1 _07543_ (.LO(_01089_));
 sky130_fd_sc_hd__conb_1 _07544_ (.LO(_01090_));
 sky130_fd_sc_hd__conb_1 _07545_ (.LO(_01091_));
 sky130_fd_sc_hd__conb_1 _07546_ (.LO(_01092_));
 sky130_fd_sc_hd__conb_1 _07547_ (.LO(_01093_));
 sky130_fd_sc_hd__conb_1 _07548_ (.LO(_01094_));
 sky130_fd_sc_hd__conb_1 _07549_ (.LO(_01095_));
 sky130_fd_sc_hd__conb_1 _07550_ (.LO(_01096_));
 sky130_fd_sc_hd__conb_1 _07551_ (.LO(_01097_));
 sky130_fd_sc_hd__conb_1 _07552_ (.LO(_01098_));
 sky130_fd_sc_hd__conb_1 _07553_ (.LO(_01099_));
 sky130_fd_sc_hd__conb_1 _07554_ (.LO(_01100_));
 sky130_fd_sc_hd__conb_1 _07555_ (.LO(_01101_));
 sky130_fd_sc_hd__conb_1 _07556_ (.LO(_01102_));
 sky130_fd_sc_hd__conb_1 _07557_ (.LO(_01103_));
 sky130_fd_sc_hd__conb_1 _07558_ (.LO(_01104_));
 sky130_fd_sc_hd__conb_1 _07559_ (.LO(_01105_));
 sky130_fd_sc_hd__conb_1 _07560_ (.LO(_01106_));
 sky130_fd_sc_hd__conb_1 _07561_ (.LO(_01107_));
 sky130_fd_sc_hd__conb_1 _07562_ (.LO(_01108_));
 sky130_fd_sc_hd__conb_1 _07563_ (.LO(_01109_));
 sky130_fd_sc_hd__conb_1 _07564_ (.LO(_01110_));
 sky130_fd_sc_hd__conb_1 _07565_ (.LO(_01111_));
 sky130_fd_sc_hd__conb_1 _07566_ (.LO(_01112_));
 sky130_fd_sc_hd__conb_1 _07567_ (.LO(_01113_));
 sky130_fd_sc_hd__conb_1 _07568_ (.LO(_01114_));
 sky130_fd_sc_hd__conb_1 _07569_ (.LO(_01115_));
 sky130_fd_sc_hd__conb_1 _07570_ (.LO(_01116_));
 sky130_fd_sc_hd__conb_1 _07571_ (.LO(_01117_));
 sky130_fd_sc_hd__conb_1 _07572_ (.LO(_01118_));
 sky130_fd_sc_hd__conb_1 _07573_ (.LO(_01119_));
 sky130_fd_sc_hd__conb_1 _07574_ (.LO(_01120_));
 sky130_fd_sc_hd__conb_1 _07575_ (.LO(_01121_));
 sky130_fd_sc_hd__conb_1 _07576_ (.LO(_01122_));
 sky130_fd_sc_hd__conb_1 _07577_ (.LO(_01123_));
 sky130_fd_sc_hd__conb_1 _07578_ (.LO(_01124_));
 sky130_fd_sc_hd__conb_1 _07579_ (.LO(_01125_));
 sky130_fd_sc_hd__conb_1 _07580_ (.LO(_01126_));
 sky130_fd_sc_hd__conb_1 _07581_ (.LO(_01127_));
 sky130_fd_sc_hd__conb_1 _07582_ (.LO(_01128_));
 sky130_fd_sc_hd__conb_1 _07583_ (.LO(_01129_));
 sky130_fd_sc_hd__conb_1 _07584_ (.LO(_01130_));
 sky130_fd_sc_hd__conb_1 _07585_ (.LO(_01131_));
 sky130_fd_sc_hd__conb_1 _07586_ (.LO(_01132_));
 sky130_fd_sc_hd__conb_1 _07587_ (.LO(_01133_));
 sky130_fd_sc_hd__conb_1 _07588_ (.LO(_01134_));
 sky130_fd_sc_hd__conb_1 _07589_ (.LO(_01135_));
 sky130_fd_sc_hd__conb_1 _07590_ (.LO(_01136_));
 sky130_fd_sc_hd__conb_1 _07591_ (.LO(_01137_));
 sky130_fd_sc_hd__conb_1 _07592_ (.LO(_01138_));
 sky130_fd_sc_hd__conb_1 _07593_ (.LO(_01139_));
 sky130_fd_sc_hd__conb_1 _07594_ (.LO(_01140_));
 sky130_fd_sc_hd__conb_1 _07595_ (.LO(_01141_));
 sky130_fd_sc_hd__conb_1 _07596_ (.LO(_01142_));
 sky130_fd_sc_hd__conb_1 _07597_ (.LO(_01143_));
 sky130_fd_sc_hd__conb_1 _07598_ (.LO(_01144_));
 sky130_fd_sc_hd__conb_1 _07599_ (.LO(_01145_));
 sky130_fd_sc_hd__conb_1 _07600_ (.LO(_01146_));
 sky130_fd_sc_hd__conb_1 _07601_ (.LO(_01147_));
 sky130_fd_sc_hd__conb_1 _07602_ (.LO(_01148_));
 sky130_fd_sc_hd__conb_1 _07603_ (.LO(_01149_));
 sky130_fd_sc_hd__conb_1 _07604_ (.LO(_01150_));
 sky130_fd_sc_hd__conb_1 _07605_ (.LO(_01151_));
 sky130_fd_sc_hd__conb_1 _07606_ (.LO(_01152_));
 sky130_fd_sc_hd__conb_1 _07607_ (.LO(_01153_));
 sky130_fd_sc_hd__conb_1 _07608_ (.LO(_01154_));
 sky130_fd_sc_hd__conb_1 _07609_ (.LO(_01155_));
 sky130_fd_sc_hd__conb_1 _07610_ (.LO(_01156_));
 sky130_fd_sc_hd__conb_1 _07611_ (.LO(_01157_));
 sky130_fd_sc_hd__conb_1 _07612_ (.LO(_01158_));
 sky130_fd_sc_hd__conb_1 _07613_ (.LO(_01159_));
 sky130_fd_sc_hd__conb_1 _07614_ (.LO(_01160_));
 sky130_fd_sc_hd__conb_1 _07615_ (.LO(_01161_));
 sky130_fd_sc_hd__conb_1 _07616_ (.LO(_01162_));
 sky130_fd_sc_hd__conb_1 _07617_ (.LO(_01163_));
 sky130_fd_sc_hd__conb_1 _07618_ (.LO(_01164_));
 sky130_fd_sc_hd__conb_1 _07619_ (.LO(_01165_));
 sky130_fd_sc_hd__conb_1 _07620_ (.LO(_01166_));
 sky130_fd_sc_hd__conb_1 _07621_ (.LO(_01167_));
 sky130_fd_sc_hd__conb_1 _07622_ (.LO(_01168_));
 sky130_fd_sc_hd__conb_1 _07623_ (.LO(_01169_));
 sky130_fd_sc_hd__conb_1 _07624_ (.LO(_01170_));
 sky130_fd_sc_hd__conb_1 _07625_ (.LO(_01171_));
 sky130_fd_sc_hd__conb_1 _07626_ (.LO(_01172_));
 sky130_fd_sc_hd__conb_1 _07627_ (.LO(_01173_));
 sky130_fd_sc_hd__conb_1 _07628_ (.LO(_01174_));
 sky130_fd_sc_hd__conb_1 _07629_ (.LO(_01175_));
 sky130_fd_sc_hd__conb_1 _07630_ (.LO(_01176_));
 sky130_fd_sc_hd__conb_1 _07631_ (.LO(_01177_));
 sky130_fd_sc_hd__conb_1 _07632_ (.LO(_01178_));
 sky130_fd_sc_hd__conb_1 _07633_ (.LO(_01179_));
 sky130_fd_sc_hd__conb_1 _07634_ (.LO(_01180_));
 sky130_fd_sc_hd__conb_1 _07635_ (.LO(_01181_));
 sky130_fd_sc_hd__conb_1 _07636_ (.LO(_01182_));
 sky130_fd_sc_hd__conb_1 _07637_ (.LO(_01183_));
 sky130_fd_sc_hd__conb_1 _07638_ (.LO(_01184_));
 sky130_fd_sc_hd__conb_1 _07639_ (.LO(_01185_));
 sky130_fd_sc_hd__conb_1 _07640_ (.LO(_01186_));
 sky130_fd_sc_hd__conb_1 _07641_ (.LO(_01187_));
 sky130_fd_sc_hd__conb_1 _07642_ (.LO(_01188_));
 sky130_fd_sc_hd__conb_1 _07643_ (.LO(_01189_));
 sky130_fd_sc_hd__conb_1 _07644_ (.LO(_01190_));
 sky130_fd_sc_hd__conb_1 _07645_ (.LO(_01191_));
 sky130_fd_sc_hd__conb_1 _07646_ (.LO(_01192_));
 sky130_fd_sc_hd__conb_1 _07647_ (.LO(_01193_));
 sky130_fd_sc_hd__conb_1 _07648_ (.LO(_01194_));
 sky130_fd_sc_hd__conb_1 _07649_ (.LO(_01195_));
 sky130_fd_sc_hd__conb_1 _07650_ (.LO(_01196_));
 sky130_fd_sc_hd__conb_1 _07651_ (.LO(_01197_));
 sky130_fd_sc_hd__conb_1 _07652_ (.LO(_01198_));
 sky130_fd_sc_hd__conb_1 _07653_ (.LO(_01199_));
 sky130_fd_sc_hd__conb_1 _07654_ (.LO(_01200_));
 sky130_fd_sc_hd__conb_1 _07655_ (.LO(_01201_));
 sky130_fd_sc_hd__conb_1 _07656_ (.LO(_01202_));
 sky130_fd_sc_hd__conb_1 _07657_ (.LO(_01203_));
 sky130_fd_sc_hd__conb_1 _07658_ (.LO(_01204_));
 sky130_fd_sc_hd__conb_1 _07659_ (.LO(_01205_));
 sky130_fd_sc_hd__conb_1 _07660_ (.LO(_01206_));
 sky130_fd_sc_hd__conb_1 _07661_ (.LO(_01207_));
 sky130_fd_sc_hd__conb_1 _07662_ (.LO(_01208_));
 sky130_fd_sc_hd__conb_1 _07663_ (.LO(_01209_));
 sky130_fd_sc_hd__conb_1 _07664_ (.LO(_01210_));
 sky130_fd_sc_hd__conb_1 _07665_ (.LO(_01211_));
 sky130_fd_sc_hd__conb_1 _07666_ (.LO(_01212_));
 sky130_fd_sc_hd__conb_1 _07667_ (.LO(_01213_));
 sky130_fd_sc_hd__conb_1 _07668_ (.LO(_01214_));
 sky130_fd_sc_hd__conb_1 _07669_ (.LO(_01215_));
 sky130_fd_sc_hd__conb_1 _07670_ (.LO(_01216_));
 sky130_fd_sc_hd__conb_1 _07671_ (.LO(_01217_));
 sky130_fd_sc_hd__conb_1 _07672_ (.LO(_01218_));
 sky130_fd_sc_hd__conb_1 _07673_ (.LO(_01219_));
 sky130_fd_sc_hd__conb_1 _07674_ (.LO(_01220_));
 sky130_fd_sc_hd__conb_1 _07675_ (.LO(_01221_));
 sky130_fd_sc_hd__conb_1 _07676_ (.LO(_01222_));
 sky130_fd_sc_hd__conb_1 _07677_ (.LO(_01223_));
 sky130_fd_sc_hd__conb_1 _07678_ (.LO(_01224_));
 sky130_fd_sc_hd__conb_1 _07679_ (.LO(_01225_));
 sky130_fd_sc_hd__conb_1 _07680_ (.LO(_01226_));
 sky130_fd_sc_hd__conb_1 _07681_ (.LO(_01227_));
 sky130_fd_sc_hd__conb_1 _07682_ (.LO(_01228_));
 sky130_fd_sc_hd__conb_1 _07683_ (.LO(_01229_));
 sky130_fd_sc_hd__conb_1 _07684_ (.LO(_01230_));
 sky130_fd_sc_hd__conb_1 _07685_ (.LO(_01231_));
 sky130_fd_sc_hd__conb_1 _07686_ (.LO(_01232_));
 sky130_fd_sc_hd__conb_1 _07687_ (.LO(_01233_));
 sky130_fd_sc_hd__conb_1 _07688_ (.LO(_01234_));
 sky130_fd_sc_hd__conb_1 _07689_ (.LO(_01235_));
 sky130_fd_sc_hd__conb_1 _07690_ (.LO(_01236_));
 sky130_fd_sc_hd__conb_1 _07691_ (.LO(_01237_));
 sky130_fd_sc_hd__conb_1 _07692_ (.LO(_01238_));
 sky130_fd_sc_hd__conb_1 _07693_ (.LO(_01239_));
 sky130_fd_sc_hd__conb_1 _07694_ (.LO(_01240_));
 sky130_fd_sc_hd__conb_1 _07695_ (.LO(_01241_));
 sky130_fd_sc_hd__conb_1 _07696_ (.LO(_01242_));
 sky130_fd_sc_hd__conb_1 _07697_ (.LO(_01243_));
 sky130_fd_sc_hd__conb_1 _07698_ (.LO(_01244_));
 sky130_fd_sc_hd__conb_1 _07699_ (.LO(_01245_));
 sky130_fd_sc_hd__conb_1 _07700_ (.LO(_01246_));
 sky130_fd_sc_hd__conb_1 _07701_ (.LO(_01247_));
 sky130_fd_sc_hd__conb_1 _07702_ (.LO(_01248_));
 sky130_fd_sc_hd__conb_1 _07703_ (.LO(_01249_));
 sky130_fd_sc_hd__conb_1 _07704_ (.LO(_01250_));
 sky130_fd_sc_hd__conb_1 _07705_ (.LO(_01251_));
 sky130_fd_sc_hd__conb_1 _07706_ (.LO(_01252_));
 sky130_fd_sc_hd__conb_1 _07707_ (.LO(_01253_));
 sky130_fd_sc_hd__conb_1 _07708_ (.LO(_01254_));
 sky130_fd_sc_hd__conb_1 _07709_ (.LO(_01255_));
 sky130_fd_sc_hd__conb_1 _07710_ (.LO(_01256_));
 sky130_fd_sc_hd__conb_1 _07711_ (.LO(_01257_));
 sky130_fd_sc_hd__conb_1 _07712_ (.LO(_01258_));
 sky130_fd_sc_hd__conb_1 _07713_ (.LO(_01259_));
 sky130_fd_sc_hd__conb_1 _07714_ (.LO(_01260_));
 sky130_fd_sc_hd__conb_1 _07715_ (.LO(_01261_));
 sky130_fd_sc_hd__conb_1 _07716_ (.LO(_01262_));
 sky130_fd_sc_hd__conb_1 _07717_ (.LO(_01263_));
 sky130_fd_sc_hd__conb_1 _07718_ (.LO(_01264_));
 sky130_fd_sc_hd__conb_1 _07719_ (.LO(_01265_));
 sky130_fd_sc_hd__conb_1 _07720_ (.LO(_01266_));
 sky130_fd_sc_hd__conb_1 _07721_ (.LO(_01267_));
 sky130_fd_sc_hd__conb_1 _07722_ (.LO(_01268_));
 sky130_fd_sc_hd__conb_1 _07723_ (.LO(_01269_));
 sky130_fd_sc_hd__conb_1 _07724_ (.LO(_01270_));
 sky130_fd_sc_hd__conb_1 _07725_ (.LO(_01271_));
 sky130_fd_sc_hd__conb_1 _07726_ (.LO(_01272_));
 sky130_fd_sc_hd__conb_1 _07727_ (.LO(_01273_));
 sky130_fd_sc_hd__conb_1 _07728_ (.LO(_01274_));
 sky130_fd_sc_hd__conb_1 _07729_ (.LO(_01275_));
 sky130_fd_sc_hd__conb_1 _07730_ (.LO(_01276_));
 sky130_fd_sc_hd__conb_1 _07731_ (.LO(_01277_));
 sky130_fd_sc_hd__conb_1 _07732_ (.LO(_01278_));
 sky130_fd_sc_hd__conb_1 _07733_ (.LO(_01279_));
 sky130_fd_sc_hd__conb_1 _07734_ (.LO(_01280_));
 sky130_fd_sc_hd__conb_1 _07735_ (.LO(_01281_));
 sky130_fd_sc_hd__conb_1 _07736_ (.LO(_01282_));
 sky130_fd_sc_hd__conb_1 _07737_ (.LO(_01283_));
 sky130_fd_sc_hd__conb_1 _07738_ (.LO(_01284_));
 sky130_fd_sc_hd__conb_1 _07739_ (.LO(_01285_));
 sky130_fd_sc_hd__conb_1 _07740_ (.LO(_01286_));
 sky130_fd_sc_hd__conb_1 _07741_ (.LO(_01287_));
 sky130_fd_sc_hd__conb_1 _07742_ (.LO(_01288_));
 sky130_fd_sc_hd__conb_1 _07743_ (.LO(_01289_));
 sky130_fd_sc_hd__conb_1 _07744_ (.LO(_01290_));
 sky130_fd_sc_hd__conb_1 _07745_ (.LO(_01291_));
 sky130_fd_sc_hd__conb_1 _07746_ (.LO(_01292_));
 sky130_fd_sc_hd__conb_1 _07747_ (.LO(_01293_));
 sky130_fd_sc_hd__conb_1 _07748_ (.LO(_01294_));
 sky130_fd_sc_hd__conb_1 _07749_ (.LO(_01295_));
 sky130_fd_sc_hd__conb_1 _07750_ (.LO(_01296_));
 sky130_fd_sc_hd__conb_1 _07751_ (.LO(_01297_));
 sky130_fd_sc_hd__conb_1 _07752_ (.LO(_01298_));
 sky130_fd_sc_hd__conb_1 _07753_ (.LO(_01299_));
 sky130_fd_sc_hd__conb_1 _07754_ (.LO(_01300_));
 sky130_fd_sc_hd__conb_1 _07755_ (.LO(_01301_));
 sky130_fd_sc_hd__conb_1 _07756_ (.LO(_01302_));
 sky130_fd_sc_hd__conb_1 _07757_ (.LO(_01303_));
 sky130_fd_sc_hd__conb_1 _07758_ (.LO(_01304_));
 sky130_fd_sc_hd__conb_1 _07759_ (.LO(_01305_));
 sky130_fd_sc_hd__conb_1 _07760_ (.LO(_01306_));
 sky130_fd_sc_hd__conb_1 _07761_ (.LO(_01307_));
 sky130_fd_sc_hd__conb_1 _07762_ (.LO(_01308_));
 sky130_fd_sc_hd__conb_1 _07763_ (.LO(_01309_));
 sky130_fd_sc_hd__conb_1 _07764_ (.LO(_01310_));
 sky130_fd_sc_hd__conb_1 _07765_ (.LO(_01311_));
 sky130_fd_sc_hd__conb_1 _07766_ (.LO(_01312_));
 sky130_fd_sc_hd__conb_1 _07767_ (.LO(_01313_));
 sky130_fd_sc_hd__conb_1 _07768_ (.LO(_01314_));
 sky130_fd_sc_hd__conb_1 _07769_ (.LO(_01315_));
 sky130_fd_sc_hd__conb_1 _07770_ (.LO(_01316_));
 sky130_fd_sc_hd__conb_1 _07771_ (.LO(_01317_));
 sky130_fd_sc_hd__conb_1 _07772_ (.LO(_01318_));
 sky130_fd_sc_hd__conb_1 _07773_ (.LO(_01319_));
 sky130_fd_sc_hd__conb_1 _07774_ (.LO(_01320_));
 sky130_fd_sc_hd__conb_1 _07775_ (.LO(_01321_));
 sky130_fd_sc_hd__conb_1 _07776_ (.LO(_01322_));
 sky130_fd_sc_hd__conb_1 _07777_ (.LO(_01323_));
 sky130_fd_sc_hd__conb_1 _07778_ (.LO(_01324_));
 sky130_fd_sc_hd__conb_1 _07779_ (.LO(_01325_));
 sky130_fd_sc_hd__conb_1 _07780_ (.LO(_01326_));
 sky130_fd_sc_hd__conb_1 _07781_ (.LO(_01327_));
 sky130_fd_sc_hd__conb_1 _07782_ (.LO(_01328_));
 sky130_fd_sc_hd__conb_1 _07783_ (.LO(_01329_));
 sky130_fd_sc_hd__conb_1 _07784_ (.LO(_01330_));
 sky130_fd_sc_hd__conb_1 _07785_ (.LO(_01331_));
 sky130_fd_sc_hd__conb_1 _07786_ (.LO(_01332_));
 sky130_fd_sc_hd__conb_1 _07787_ (.LO(_01333_));
 sky130_fd_sc_hd__conb_1 _07788_ (.LO(_01334_));
 sky130_fd_sc_hd__conb_1 _07789_ (.LO(_01335_));
 sky130_fd_sc_hd__conb_1 _07790_ (.LO(_01336_));
 sky130_fd_sc_hd__conb_1 _07791_ (.LO(_01337_));
 sky130_fd_sc_hd__conb_1 _07792_ (.LO(_01338_));
 sky130_fd_sc_hd__conb_1 _07793_ (.LO(_01339_));
 sky130_fd_sc_hd__conb_1 _07794_ (.LO(_01340_));
 sky130_fd_sc_hd__conb_1 _07795_ (.LO(_01341_));
 sky130_fd_sc_hd__conb_1 _07796_ (.LO(_01342_));
 sky130_fd_sc_hd__conb_1 _07797_ (.LO(_01343_));
 sky130_fd_sc_hd__conb_1 _07798_ (.LO(_01344_));
 sky130_fd_sc_hd__conb_1 _07799_ (.LO(_01345_));
 sky130_fd_sc_hd__conb_1 _07800_ (.LO(_01346_));
 sky130_fd_sc_hd__conb_1 _07801_ (.LO(_01347_));
 sky130_fd_sc_hd__conb_1 _07802_ (.LO(_01348_));
 sky130_fd_sc_hd__conb_1 _07803_ (.LO(_01349_));
 sky130_fd_sc_hd__conb_1 _07804_ (.LO(_01350_));
 sky130_fd_sc_hd__conb_1 _07805_ (.LO(_01351_));
 sky130_fd_sc_hd__conb_1 _07806_ (.LO(_01352_));
 sky130_fd_sc_hd__conb_1 _07807_ (.LO(_01353_));
 sky130_fd_sc_hd__conb_1 _07808_ (.LO(_01354_));
 sky130_fd_sc_hd__conb_1 _07809_ (.LO(_01355_));
 sky130_fd_sc_hd__conb_1 _07810_ (.LO(_01356_));
 sky130_fd_sc_hd__conb_1 _07811_ (.LO(_01357_));
 sky130_fd_sc_hd__conb_1 _07812_ (.LO(_01358_));
 sky130_fd_sc_hd__conb_1 _07813_ (.LO(_01359_));
 sky130_fd_sc_hd__conb_1 _07814_ (.LO(_01360_));
 sky130_fd_sc_hd__conb_1 _07815_ (.LO(_01361_));
 sky130_fd_sc_hd__conb_1 _07816_ (.LO(_01362_));
 sky130_fd_sc_hd__conb_1 _07817_ (.LO(_01363_));
 sky130_fd_sc_hd__conb_1 _07818_ (.LO(_01364_));
 sky130_fd_sc_hd__conb_1 _07819_ (.LO(_01365_));
 sky130_fd_sc_hd__conb_1 _07820_ (.LO(_01366_));
 sky130_fd_sc_hd__conb_1 _07821_ (.LO(_01367_));
 sky130_fd_sc_hd__conb_1 _07822_ (.LO(_01368_));
 sky130_fd_sc_hd__conb_1 _07823_ (.LO(_01369_));
 sky130_fd_sc_hd__conb_1 _07824_ (.LO(_01370_));
 sky130_fd_sc_hd__conb_1 _07825_ (.LO(_01371_));
 sky130_fd_sc_hd__conb_1 _07826_ (.LO(_01372_));
 sky130_fd_sc_hd__conb_1 _07827_ (.LO(_01373_));
 sky130_fd_sc_hd__conb_1 _07828_ (.LO(_01374_));
 sky130_fd_sc_hd__conb_1 _07829_ (.LO(_01375_));
 sky130_fd_sc_hd__conb_1 _07830_ (.LO(_01376_));
 sky130_fd_sc_hd__conb_1 _07831_ (.LO(_01377_));
 sky130_fd_sc_hd__conb_1 _07832_ (.LO(_01378_));
 sky130_fd_sc_hd__conb_1 _07833_ (.LO(_01379_));
 sky130_fd_sc_hd__conb_1 _07834_ (.LO(_01380_));
 sky130_fd_sc_hd__conb_1 _07835_ (.LO(_01381_));
 sky130_fd_sc_hd__conb_1 _07836_ (.LO(_01382_));
 sky130_fd_sc_hd__conb_1 _07837_ (.LO(_01383_));
 sky130_fd_sc_hd__conb_1 _07838_ (.LO(_01384_));
 sky130_fd_sc_hd__conb_1 _07839_ (.LO(_01385_));
 sky130_fd_sc_hd__conb_1 _07840_ (.LO(_01386_));
 sky130_fd_sc_hd__conb_1 _07841_ (.LO(_01387_));
 sky130_fd_sc_hd__conb_1 _07842_ (.LO(_01388_));
 sky130_fd_sc_hd__conb_1 _07843_ (.LO(_01389_));
 sky130_fd_sc_hd__conb_1 _07844_ (.LO(_01390_));
 sky130_fd_sc_hd__conb_1 _07845_ (.LO(_01391_));
 sky130_fd_sc_hd__conb_1 _07846_ (.LO(_01392_));
 sky130_fd_sc_hd__conb_1 _07847_ (.LO(_01393_));
 sky130_fd_sc_hd__conb_1 _07848_ (.LO(_01394_));
 sky130_fd_sc_hd__conb_1 _07849_ (.LO(_01395_));
 sky130_fd_sc_hd__conb_1 _07850_ (.LO(_01396_));
 sky130_fd_sc_hd__conb_1 _07851_ (.LO(_01397_));
 sky130_fd_sc_hd__conb_1 _07852_ (.LO(_01398_));
 sky130_fd_sc_hd__conb_1 _07853_ (.LO(_01399_));
 sky130_fd_sc_hd__conb_1 _07854_ (.LO(_01400_));
 sky130_fd_sc_hd__conb_1 _07855_ (.LO(_01401_));
 sky130_fd_sc_hd__conb_1 _07856_ (.LO(_01402_));
 sky130_fd_sc_hd__conb_1 _07857_ (.LO(_01403_));
 sky130_fd_sc_hd__conb_1 _07858_ (.LO(_01404_));
 sky130_fd_sc_hd__conb_1 _07859_ (.LO(_01405_));
 sky130_fd_sc_hd__conb_1 _07860_ (.LO(_01406_));
 sky130_fd_sc_hd__conb_1 _07861_ (.LO(_01407_));
 sky130_fd_sc_hd__conb_1 _07862_ (.LO(_01408_));
 sky130_fd_sc_hd__conb_1 _07863_ (.LO(_01409_));
 sky130_fd_sc_hd__conb_1 _07864_ (.LO(_01410_));
 sky130_fd_sc_hd__conb_1 _07865_ (.LO(_01411_));
 sky130_fd_sc_hd__conb_1 _07866_ (.LO(_01412_));
 sky130_fd_sc_hd__conb_1 _07867_ (.LO(_01413_));
 sky130_fd_sc_hd__conb_1 _07868_ (.LO(_01414_));
 sky130_fd_sc_hd__conb_1 _07869_ (.LO(_01415_));
 sky130_fd_sc_hd__conb_1 _07870_ (.LO(_01416_));
 sky130_fd_sc_hd__conb_1 _07871_ (.LO(_01417_));
 sky130_fd_sc_hd__conb_1 _07872_ (.LO(_01418_));
 sky130_fd_sc_hd__conb_1 _07873_ (.LO(_01419_));
 sky130_fd_sc_hd__conb_1 _07874_ (.LO(_01420_));
 sky130_fd_sc_hd__conb_1 _07875_ (.LO(_01421_));
 sky130_fd_sc_hd__conb_1 _07876_ (.LO(_01422_));
 sky130_fd_sc_hd__conb_1 _07877_ (.LO(_01423_));
 sky130_fd_sc_hd__conb_1 _07878_ (.LO(_01424_));
 sky130_fd_sc_hd__conb_1 _07879_ (.LO(_01425_));
 sky130_fd_sc_hd__conb_1 _07880_ (.LO(_01426_));
 sky130_fd_sc_hd__conb_1 _07881_ (.LO(_01427_));
 sky130_fd_sc_hd__conb_1 _07882_ (.LO(_01428_));
 sky130_fd_sc_hd__conb_1 _07883_ (.LO(_01429_));
 sky130_fd_sc_hd__conb_1 _07884_ (.LO(_01430_));
 sky130_fd_sc_hd__conb_1 _07885_ (.LO(_01431_));
 sky130_fd_sc_hd__conb_1 _07886_ (.LO(_01432_));
 sky130_fd_sc_hd__conb_1 _07887_ (.LO(_01433_));
 sky130_fd_sc_hd__conb_1 _07888_ (.LO(_01434_));
 sky130_fd_sc_hd__conb_1 _07889_ (.LO(_01435_));
 sky130_fd_sc_hd__conb_1 _07890_ (.LO(_01436_));
 sky130_fd_sc_hd__conb_1 _07891_ (.LO(_01437_));
 sky130_fd_sc_hd__conb_1 _07892_ (.LO(_01438_));
 sky130_fd_sc_hd__conb_1 _07893_ (.LO(_01439_));
 sky130_fd_sc_hd__conb_1 _07894_ (.LO(_01440_));
 sky130_fd_sc_hd__conb_1 _07895_ (.LO(_01441_));
 sky130_fd_sc_hd__conb_1 _07896_ (.LO(_01442_));
 sky130_fd_sc_hd__conb_1 _07897_ (.LO(_01443_));
 sky130_fd_sc_hd__conb_1 _07898_ (.LO(_01444_));
 sky130_fd_sc_hd__conb_1 _07899_ (.LO(_01445_));
 sky130_fd_sc_hd__conb_1 _07900_ (.LO(_01446_));
 sky130_fd_sc_hd__conb_1 _07901_ (.LO(_01447_));
 sky130_fd_sc_hd__conb_1 _07902_ (.LO(_01448_));
 sky130_fd_sc_hd__conb_1 _07903_ (.LO(_01449_));
 sky130_fd_sc_hd__conb_1 _07904_ (.LO(_01450_));
 sky130_fd_sc_hd__conb_1 _07905_ (.LO(_01451_));
 sky130_fd_sc_hd__conb_1 _07906_ (.LO(_01452_));
 sky130_fd_sc_hd__conb_1 _07907_ (.LO(_01453_));
 sky130_fd_sc_hd__conb_1 _07908_ (.LO(_01454_));
 sky130_fd_sc_hd__conb_1 _07909_ (.LO(_01455_));
 sky130_fd_sc_hd__conb_1 _07910_ (.LO(_01456_));
 sky130_fd_sc_hd__conb_1 _07911_ (.LO(_01457_));
 sky130_fd_sc_hd__conb_1 _07912_ (.LO(_01458_));
 sky130_fd_sc_hd__conb_1 _07913_ (.LO(_01459_));
 sky130_fd_sc_hd__conb_1 _07914_ (.LO(_01460_));
 sky130_fd_sc_hd__conb_1 _07915_ (.LO(_01461_));
 sky130_fd_sc_hd__conb_1 _07916_ (.LO(_01462_));
 sky130_fd_sc_hd__conb_1 _07917_ (.LO(_01463_));
 sky130_fd_sc_hd__conb_1 _07918_ (.LO(_01464_));
 sky130_fd_sc_hd__conb_1 _07919_ (.LO(_01465_));
 sky130_fd_sc_hd__conb_1 _07920_ (.LO(_01466_));
 sky130_fd_sc_hd__conb_1 _07921_ (.LO(_01467_));
 sky130_fd_sc_hd__conb_1 _07922_ (.LO(_01468_));
 sky130_fd_sc_hd__conb_1 _07923_ (.LO(_01469_));
 sky130_fd_sc_hd__conb_1 _07924_ (.LO(_01470_));
 sky130_fd_sc_hd__conb_1 _07925_ (.LO(_01471_));
 sky130_fd_sc_hd__conb_1 _07926_ (.LO(_01472_));
 sky130_fd_sc_hd__conb_1 _07927_ (.LO(_01473_));
 sky130_fd_sc_hd__conb_1 _07928_ (.LO(_01474_));
 sky130_fd_sc_hd__conb_1 _07929_ (.LO(_01475_));
 sky130_fd_sc_hd__conb_1 _07930_ (.LO(_01476_));
 sky130_fd_sc_hd__conb_1 _07931_ (.LO(_01477_));
 sky130_fd_sc_hd__conb_1 _07932_ (.LO(_01478_));
 sky130_fd_sc_hd__conb_1 _07933_ (.LO(_01479_));
 sky130_fd_sc_hd__conb_1 _07934_ (.LO(_01480_));
 sky130_fd_sc_hd__conb_1 _07935_ (.LO(_01481_));
 sky130_fd_sc_hd__conb_1 _07936_ (.LO(_01482_));
 sky130_fd_sc_hd__conb_1 _07937_ (.LO(_01483_));
 sky130_fd_sc_hd__conb_1 _07938_ (.LO(_01484_));
 sky130_fd_sc_hd__conb_1 _07939_ (.LO(_01485_));
 sky130_fd_sc_hd__conb_1 _07940_ (.LO(_01486_));
 sky130_fd_sc_hd__conb_1 _07941_ (.LO(_01487_));
 sky130_fd_sc_hd__conb_1 _07942_ (.LO(_01488_));
 sky130_fd_sc_hd__conb_1 _07943_ (.LO(_01489_));
 sky130_fd_sc_hd__conb_1 _07944_ (.LO(_01490_));
 sky130_fd_sc_hd__conb_1 _07945_ (.LO(_01491_));
 sky130_fd_sc_hd__conb_1 _07946_ (.LO(_01492_));
 sky130_fd_sc_hd__conb_1 _07947_ (.LO(_01493_));
 sky130_fd_sc_hd__conb_1 _07948_ (.LO(_01494_));
 sky130_fd_sc_hd__conb_1 _07949_ (.LO(_01495_));
 sky130_fd_sc_hd__conb_1 _07950_ (.LO(_01496_));
 sky130_fd_sc_hd__conb_1 _07951_ (.LO(_01497_));
 sky130_fd_sc_hd__conb_1 _07952_ (.LO(_01498_));
 sky130_fd_sc_hd__conb_1 _07953_ (.LO(_01499_));
 sky130_fd_sc_hd__conb_1 _07954_ (.LO(_01500_));
 sky130_fd_sc_hd__conb_1 _07955_ (.LO(_01501_));
 sky130_fd_sc_hd__conb_1 _07956_ (.LO(_01502_));
 sky130_fd_sc_hd__conb_1 _07957_ (.LO(_01503_));
 sky130_fd_sc_hd__conb_1 _07958_ (.LO(_01504_));
 sky130_fd_sc_hd__conb_1 _07959_ (.LO(_01505_));
 sky130_fd_sc_hd__conb_1 _07960_ (.LO(_01506_));
 sky130_fd_sc_hd__conb_1 _07961_ (.LO(_01507_));
 sky130_fd_sc_hd__conb_1 _07962_ (.LO(_01508_));
 sky130_fd_sc_hd__conb_1 _07963_ (.LO(_01509_));
 sky130_fd_sc_hd__conb_1 _07964_ (.LO(_01510_));
 sky130_fd_sc_hd__conb_1 _07965_ (.LO(_01511_));
 sky130_fd_sc_hd__conb_1 _07966_ (.LO(_01512_));
 sky130_fd_sc_hd__conb_1 _07967_ (.LO(_01513_));
 sky130_fd_sc_hd__conb_1 _07968_ (.LO(_01514_));
 sky130_fd_sc_hd__conb_1 _07969_ (.LO(_01515_));
 sky130_fd_sc_hd__conb_1 _07970_ (.LO(_01516_));
 sky130_fd_sc_hd__conb_1 _07971_ (.LO(_01517_));
 sky130_fd_sc_hd__conb_1 _07972_ (.LO(_01518_));
 sky130_fd_sc_hd__conb_1 _07973_ (.LO(_01519_));
 sky130_fd_sc_hd__conb_1 _07974_ (.LO(_01520_));
 sky130_fd_sc_hd__conb_1 _07975_ (.LO(_01521_));
 sky130_fd_sc_hd__conb_1 _07976_ (.LO(_01522_));
 sky130_fd_sc_hd__conb_1 _07977_ (.LO(_01523_));
 sky130_fd_sc_hd__conb_1 _07978_ (.LO(_01524_));
 sky130_fd_sc_hd__conb_1 _07979_ (.LO(_01525_));
 sky130_fd_sc_hd__conb_1 _07980_ (.LO(_01526_));
 sky130_fd_sc_hd__conb_1 _07981_ (.LO(_01527_));
 sky130_fd_sc_hd__conb_1 _07982_ (.LO(_01528_));
 sky130_fd_sc_hd__conb_1 _07983_ (.LO(_01529_));
 sky130_fd_sc_hd__conb_1 _07984_ (.LO(_01530_));
 sky130_fd_sc_hd__conb_1 _07985_ (.LO(_01531_));
 sky130_fd_sc_hd__conb_1 _07986_ (.LO(_01532_));
 sky130_fd_sc_hd__conb_1 _07987_ (.LO(_01533_));
 sky130_fd_sc_hd__conb_1 _07988_ (.LO(_01534_));
 sky130_fd_sc_hd__conb_1 _07989_ (.LO(_01535_));
 sky130_fd_sc_hd__conb_1 _07990_ (.LO(_01536_));
 sky130_fd_sc_hd__conb_1 _07991_ (.LO(_01537_));
 sky130_fd_sc_hd__conb_1 _07992_ (.LO(_01538_));
 sky130_fd_sc_hd__conb_1 _07993_ (.LO(_01539_));
 sky130_fd_sc_hd__conb_1 _07994_ (.LO(_01540_));
 sky130_fd_sc_hd__conb_1 _07995_ (.LO(_01541_));
 sky130_fd_sc_hd__conb_1 _07996_ (.LO(_01542_));
 sky130_fd_sc_hd__conb_1 _07997_ (.LO(_01543_));
 sky130_fd_sc_hd__conb_1 _07998_ (.LO(_01544_));
 sky130_fd_sc_hd__conb_1 _07999_ (.LO(_01545_));
 sky130_fd_sc_hd__conb_1 _08000_ (.LO(_01546_));
 sky130_fd_sc_hd__conb_1 _08001_ (.LO(_01547_));
 sky130_fd_sc_hd__conb_1 _08002_ (.LO(_01548_));
 sky130_fd_sc_hd__conb_1 _08003_ (.LO(_01549_));
 sky130_fd_sc_hd__conb_1 _08004_ (.LO(_01550_));
 sky130_fd_sc_hd__conb_1 _08005_ (.LO(_01551_));
 sky130_fd_sc_hd__conb_1 _08006_ (.LO(_01552_));
 sky130_fd_sc_hd__conb_1 _08007_ (.LO(_01553_));
 sky130_fd_sc_hd__conb_1 _08008_ (.LO(_01554_));
 sky130_fd_sc_hd__conb_1 _08009_ (.LO(_01555_));
 sky130_fd_sc_hd__conb_1 _08010_ (.LO(_01556_));
 sky130_fd_sc_hd__conb_1 _08011_ (.LO(_01557_));
 sky130_fd_sc_hd__conb_1 _08012_ (.LO(_01558_));
 sky130_fd_sc_hd__conb_1 _08013_ (.LO(_01559_));
 sky130_fd_sc_hd__conb_1 _08014_ (.LO(_01560_));
 sky130_fd_sc_hd__conb_1 _08015_ (.LO(_01561_));
 sky130_fd_sc_hd__conb_1 _08016_ (.LO(_01562_));
 sky130_fd_sc_hd__conb_1 _08017_ (.LO(_01563_));
 sky130_fd_sc_hd__conb_1 _08018_ (.LO(_01564_));
 sky130_fd_sc_hd__conb_1 _08019_ (.LO(_01565_));
 sky130_fd_sc_hd__conb_1 _08020_ (.LO(_01566_));
 sky130_fd_sc_hd__conb_1 _08021_ (.LO(_01567_));
 sky130_fd_sc_hd__conb_1 _08022_ (.LO(_01568_));
 sky130_fd_sc_hd__conb_1 _08023_ (.LO(_01569_));
 sky130_fd_sc_hd__conb_1 _08024_ (.LO(_01570_));
 sky130_fd_sc_hd__conb_1 _08025_ (.LO(_01571_));
 sky130_fd_sc_hd__conb_1 _08026_ (.LO(_01572_));
 sky130_fd_sc_hd__conb_1 _08027_ (.LO(_01573_));
 sky130_fd_sc_hd__conb_1 _08028_ (.LO(_01574_));
 sky130_fd_sc_hd__conb_1 _08029_ (.LO(_01575_));
 sky130_fd_sc_hd__conb_1 _08030_ (.LO(_01576_));
 sky130_fd_sc_hd__conb_1 _08031_ (.LO(_01577_));
 sky130_fd_sc_hd__conb_1 _08032_ (.LO(_01578_));
 sky130_fd_sc_hd__conb_1 _08033_ (.LO(_01579_));
 sky130_fd_sc_hd__conb_1 _08034_ (.LO(_01580_));
 sky130_fd_sc_hd__conb_1 _08035_ (.LO(_01581_));
 sky130_fd_sc_hd__conb_1 _08036_ (.LO(_01582_));
 sky130_fd_sc_hd__conb_1 _08037_ (.LO(_01583_));
 sky130_fd_sc_hd__conb_1 _08038_ (.LO(_01584_));
 sky130_fd_sc_hd__conb_1 _08039_ (.LO(_01585_));
 sky130_fd_sc_hd__conb_1 _08040_ (.LO(_01586_));
 sky130_fd_sc_hd__conb_1 _08041_ (.LO(_01587_));
 sky130_fd_sc_hd__conb_1 _08042_ (.LO(_01588_));
 sky130_fd_sc_hd__conb_1 _08043_ (.LO(_01589_));
 sky130_fd_sc_hd__conb_1 _08044_ (.LO(_01590_));
 sky130_fd_sc_hd__conb_1 _08045_ (.LO(_01591_));
 sky130_fd_sc_hd__conb_1 _08046_ (.LO(_01592_));
 sky130_fd_sc_hd__conb_1 _08047_ (.LO(_01593_));
 sky130_fd_sc_hd__conb_1 _08048_ (.LO(_01594_));
 sky130_fd_sc_hd__conb_1 _08049_ (.LO(_01595_));
 sky130_fd_sc_hd__conb_1 _08050_ (.LO(_01596_));
 sky130_fd_sc_hd__conb_1 _08051_ (.LO(_01597_));
 sky130_fd_sc_hd__conb_1 _08052_ (.LO(_01598_));
 sky130_fd_sc_hd__conb_1 _08053_ (.LO(_01599_));
 sky130_fd_sc_hd__conb_1 _08054_ (.LO(_01600_));
 sky130_fd_sc_hd__conb_1 _08055_ (.LO(_01601_));
 sky130_fd_sc_hd__conb_1 _08056_ (.LO(_01602_));
 sky130_fd_sc_hd__conb_1 _08057_ (.LO(_01603_));
 sky130_fd_sc_hd__conb_1 _08058_ (.LO(_01604_));
 sky130_fd_sc_hd__conb_1 _08059_ (.LO(_01605_));
 sky130_fd_sc_hd__conb_1 _08060_ (.LO(_01606_));
 sky130_fd_sc_hd__conb_1 _08061_ (.LO(_01607_));
 sky130_fd_sc_hd__conb_1 _08062_ (.LO(_01608_));
 sky130_fd_sc_hd__conb_1 _08063_ (.LO(_01609_));
 sky130_fd_sc_hd__conb_1 _08064_ (.LO(_01610_));
 sky130_fd_sc_hd__conb_1 _08065_ (.LO(_01611_));
 sky130_fd_sc_hd__conb_1 _08066_ (.LO(_01612_));
 sky130_fd_sc_hd__conb_1 _08067_ (.LO(_01613_));
 sky130_fd_sc_hd__conb_1 _08068_ (.LO(_01614_));
 sky130_fd_sc_hd__conb_1 _08069_ (.LO(_01615_));
 sky130_fd_sc_hd__conb_1 _08070_ (.LO(_01616_));
 sky130_fd_sc_hd__conb_1 _08071_ (.LO(_01617_));
 sky130_fd_sc_hd__conb_1 _08072_ (.LO(_01618_));
 sky130_fd_sc_hd__conb_1 _08073_ (.LO(_01619_));
 sky130_fd_sc_hd__conb_1 _08074_ (.LO(_01620_));
 sky130_fd_sc_hd__conb_1 _08075_ (.LO(_01621_));
 sky130_fd_sc_hd__conb_1 _08076_ (.LO(_01622_));
 sky130_fd_sc_hd__conb_1 _08077_ (.LO(_01623_));
 sky130_fd_sc_hd__conb_1 _08078_ (.LO(_01624_));
 sky130_fd_sc_hd__conb_1 _08079_ (.LO(_01625_));
 sky130_fd_sc_hd__conb_1 _08080_ (.LO(_01626_));
 sky130_fd_sc_hd__conb_1 _08081_ (.LO(_01627_));
 sky130_fd_sc_hd__conb_1 _08082_ (.LO(_01628_));
 sky130_fd_sc_hd__conb_1 _08083_ (.LO(_01629_));
 sky130_fd_sc_hd__conb_1 _08084_ (.LO(_01630_));
 sky130_fd_sc_hd__conb_1 _08085_ (.LO(_01631_));
 sky130_fd_sc_hd__conb_1 _08086_ (.LO(_01632_));
 sky130_fd_sc_hd__conb_1 _08087_ (.LO(_01633_));
 sky130_fd_sc_hd__conb_1 _08088_ (.LO(_01634_));
 sky130_fd_sc_hd__conb_1 _08089_ (.LO(_01635_));
 sky130_fd_sc_hd__conb_1 _08090_ (.LO(_01636_));
 sky130_fd_sc_hd__conb_1 _08091_ (.LO(_01637_));
 sky130_fd_sc_hd__conb_1 _08092_ (.LO(_01638_));
 sky130_fd_sc_hd__conb_1 _08093_ (.LO(_01639_));
 sky130_fd_sc_hd__conb_1 _08094_ (.LO(_01640_));
 sky130_fd_sc_hd__conb_1 _08095_ (.LO(_01641_));
 sky130_fd_sc_hd__conb_1 _08096_ (.LO(_01642_));
 sky130_fd_sc_hd__conb_1 _08097_ (.LO(_01643_));
 sky130_fd_sc_hd__conb_1 _08098_ (.LO(_01644_));
 sky130_fd_sc_hd__conb_1 _08099_ (.LO(_01645_));
 sky130_fd_sc_hd__conb_1 _08100_ (.LO(_01646_));
 sky130_fd_sc_hd__conb_1 _08101_ (.LO(_01647_));
 sky130_fd_sc_hd__conb_1 _08102_ (.LO(_01648_));
 sky130_fd_sc_hd__conb_1 _08103_ (.LO(_01649_));
 sky130_fd_sc_hd__conb_1 _08104_ (.LO(_01650_));
 sky130_fd_sc_hd__conb_1 _08105_ (.LO(_01651_));
 sky130_fd_sc_hd__conb_1 _08106_ (.LO(_01652_));
 sky130_fd_sc_hd__conb_1 _08107_ (.LO(_01653_));
 sky130_fd_sc_hd__conb_1 _08108_ (.LO(_01654_));
 sky130_fd_sc_hd__conb_1 _08109_ (.LO(_01655_));
 sky130_fd_sc_hd__conb_1 _08110_ (.LO(_01656_));
 sky130_fd_sc_hd__conb_1 _08111_ (.LO(_01657_));
 sky130_fd_sc_hd__conb_1 _08112_ (.LO(_01658_));
 sky130_fd_sc_hd__conb_1 _08113_ (.LO(_01659_));
 sky130_fd_sc_hd__conb_1 _08114_ (.LO(_01660_));
 sky130_fd_sc_hd__conb_1 _08115_ (.LO(_01661_));
 sky130_fd_sc_hd__conb_1 _08116_ (.LO(_01662_));
 sky130_fd_sc_hd__conb_1 _08117_ (.LO(_01663_));
 sky130_fd_sc_hd__conb_1 _08118_ (.LO(_01664_));
 sky130_fd_sc_hd__conb_1 _08119_ (.LO(_01665_));
 sky130_fd_sc_hd__conb_1 _08120_ (.LO(_01666_));
 sky130_fd_sc_hd__conb_1 _08121_ (.LO(_01667_));
 sky130_fd_sc_hd__conb_1 _08122_ (.LO(_01668_));
 sky130_fd_sc_hd__conb_1 _08123_ (.LO(_01669_));
 sky130_fd_sc_hd__conb_1 _08124_ (.LO(_01670_));
 sky130_fd_sc_hd__conb_1 _08125_ (.LO(_01671_));
 sky130_fd_sc_hd__conb_1 _08126_ (.LO(_01672_));
 sky130_fd_sc_hd__conb_1 _08127_ (.LO(_01673_));
 sky130_fd_sc_hd__conb_1 _08128_ (.LO(_01674_));
 sky130_fd_sc_hd__conb_1 _08129_ (.LO(_01675_));
 sky130_fd_sc_hd__conb_1 _08130_ (.LO(_01676_));
 sky130_fd_sc_hd__conb_1 _08131_ (.LO(_01677_));
 sky130_fd_sc_hd__conb_1 _08132_ (.LO(_01678_));
 sky130_fd_sc_hd__conb_1 _08133_ (.LO(_01679_));
 sky130_fd_sc_hd__conb_1 _08134_ (.LO(_01680_));
 sky130_fd_sc_hd__conb_1 _08135_ (.LO(_01681_));
 sky130_fd_sc_hd__conb_1 _08136_ (.LO(_01682_));
 sky130_fd_sc_hd__conb_1 _08137_ (.LO(_01683_));
 sky130_fd_sc_hd__conb_1 _08138_ (.LO(_01684_));
 sky130_fd_sc_hd__conb_1 _08139_ (.LO(_01685_));
 sky130_fd_sc_hd__conb_1 _08140_ (.LO(_01686_));
 sky130_fd_sc_hd__conb_1 _08141_ (.LO(_01687_));
 sky130_fd_sc_hd__conb_1 _08142_ (.LO(_01688_));
 sky130_fd_sc_hd__conb_1 _08143_ (.LO(_01689_));
 sky130_fd_sc_hd__conb_1 _08144_ (.LO(_01690_));
 sky130_fd_sc_hd__conb_1 _08145_ (.LO(_01691_));
 sky130_fd_sc_hd__conb_1 _08146_ (.LO(_01692_));
 sky130_fd_sc_hd__conb_1 _08147_ (.LO(_01693_));
 sky130_fd_sc_hd__conb_1 _08148_ (.LO(_01694_));
 sky130_fd_sc_hd__conb_1 _08149_ (.LO(_01695_));
 sky130_fd_sc_hd__conb_1 _08150_ (.LO(_01696_));
 sky130_fd_sc_hd__conb_1 _08151_ (.LO(_01697_));
 sky130_fd_sc_hd__conb_1 _08152_ (.LO(_01698_));
 sky130_fd_sc_hd__conb_1 _08153_ (.LO(_01699_));
 sky130_fd_sc_hd__conb_1 _08154_ (.LO(_01700_));
 sky130_fd_sc_hd__conb_1 _08155_ (.LO(_01701_));
 sky130_fd_sc_hd__conb_1 _08156_ (.LO(_01702_));
 sky130_fd_sc_hd__conb_1 _08157_ (.LO(_01703_));
 sky130_fd_sc_hd__conb_1 _08158_ (.LO(_01704_));
 sky130_fd_sc_hd__conb_1 _08159_ (.LO(_01705_));
 sky130_fd_sc_hd__conb_1 _08160_ (.LO(_01706_));
 sky130_fd_sc_hd__conb_1 _08161_ (.LO(_01707_));
 sky130_fd_sc_hd__conb_1 _08162_ (.LO(_01708_));
 sky130_fd_sc_hd__conb_1 _08163_ (.LO(_01709_));
 sky130_fd_sc_hd__conb_1 _08164_ (.LO(_01710_));
 sky130_fd_sc_hd__conb_1 _08165_ (.LO(_01711_));
 sky130_fd_sc_hd__conb_1 _08166_ (.LO(_01712_));
 sky130_fd_sc_hd__conb_1 _08167_ (.LO(_01713_));
 sky130_fd_sc_hd__conb_1 _08168_ (.LO(_01714_));
 sky130_fd_sc_hd__conb_1 _08169_ (.LO(_01715_));
 sky130_fd_sc_hd__conb_1 _08170_ (.LO(_01716_));
 sky130_fd_sc_hd__conb_1 _08171_ (.LO(_01717_));
 sky130_fd_sc_hd__conb_1 _08172_ (.LO(_01718_));
 sky130_fd_sc_hd__conb_1 _08173_ (.LO(_01719_));
 sky130_fd_sc_hd__conb_1 _08174_ (.LO(_01720_));
 sky130_fd_sc_hd__conb_1 _08175_ (.LO(_01721_));
 sky130_fd_sc_hd__conb_1 _08176_ (.LO(_01722_));
 sky130_fd_sc_hd__conb_1 _08177_ (.LO(_01723_));
 sky130_fd_sc_hd__conb_1 _08178_ (.LO(_01724_));
 sky130_fd_sc_hd__conb_1 _08179_ (.LO(_01725_));
 sky130_fd_sc_hd__conb_1 _08180_ (.LO(_01726_));
 sky130_fd_sc_hd__conb_1 _08181_ (.LO(_01727_));
 sky130_fd_sc_hd__conb_1 _08182_ (.LO(_01728_));
 sky130_fd_sc_hd__conb_1 _08183_ (.LO(_01729_));
 sky130_fd_sc_hd__conb_1 _08184_ (.LO(_01730_));
 sky130_fd_sc_hd__conb_1 _08185_ (.LO(_01731_));
 sky130_fd_sc_hd__conb_1 _08186_ (.LO(_01732_));
 sky130_fd_sc_hd__conb_1 _08187_ (.LO(_01733_));
 sky130_fd_sc_hd__conb_1 _08188_ (.LO(_01734_));
 sky130_fd_sc_hd__conb_1 _08189_ (.LO(_01735_));
 sky130_fd_sc_hd__conb_1 _08190_ (.LO(_01736_));
 sky130_fd_sc_hd__conb_1 _08191_ (.LO(_01737_));
 sky130_fd_sc_hd__conb_1 _08192_ (.LO(_01738_));
 sky130_fd_sc_hd__conb_1 _08193_ (.LO(_01739_));
 sky130_fd_sc_hd__conb_1 _08194_ (.LO(_01740_));
 sky130_fd_sc_hd__conb_1 _08195_ (.LO(_01741_));
 sky130_fd_sc_hd__conb_1 _08196_ (.LO(_01742_));
 sky130_fd_sc_hd__conb_1 _08197_ (.LO(_01743_));
 sky130_fd_sc_hd__conb_1 _08198_ (.LO(_01744_));
 sky130_fd_sc_hd__conb_1 _08199_ (.LO(_01745_));
 sky130_fd_sc_hd__conb_1 _08200_ (.LO(_01746_));
 sky130_fd_sc_hd__conb_1 _08201_ (.LO(_01747_));
 sky130_fd_sc_hd__conb_1 _08202_ (.LO(_01748_));
 sky130_fd_sc_hd__conb_1 _08203_ (.LO(_01749_));
 sky130_fd_sc_hd__conb_1 _08204_ (.LO(_01750_));
 sky130_fd_sc_hd__conb_1 _08205_ (.LO(_01751_));
 sky130_fd_sc_hd__conb_1 _08206_ (.LO(_01752_));
 sky130_fd_sc_hd__conb_1 _08207_ (.LO(_01753_));
 sky130_fd_sc_hd__conb_1 _08208_ (.LO(_01754_));
 sky130_fd_sc_hd__conb_1 _08209_ (.LO(_01755_));
 sky130_fd_sc_hd__conb_1 _08210_ (.LO(_01756_));
 sky130_fd_sc_hd__conb_1 _08211_ (.LO(_01757_));
 sky130_fd_sc_hd__conb_1 _08212_ (.LO(_01758_));
 sky130_fd_sc_hd__conb_1 _08213_ (.LO(_01759_));
 sky130_fd_sc_hd__conb_1 _08214_ (.LO(_01760_));
 sky130_fd_sc_hd__conb_1 _08215_ (.LO(_01761_));
 sky130_fd_sc_hd__conb_1 _08216_ (.LO(_01762_));
 sky130_fd_sc_hd__conb_1 _08217_ (.LO(_01763_));
 sky130_fd_sc_hd__conb_1 _08218_ (.LO(_01764_));
 sky130_fd_sc_hd__conb_1 _08219_ (.LO(_01765_));
 sky130_fd_sc_hd__conb_1 _08220_ (.LO(_01766_));
 sky130_fd_sc_hd__conb_1 _08221_ (.LO(_01767_));
 sky130_fd_sc_hd__conb_1 _08222_ (.LO(_01768_));
 sky130_fd_sc_hd__conb_1 _08223_ (.LO(_01769_));
 sky130_fd_sc_hd__conb_1 _08224_ (.LO(_01770_));
 sky130_fd_sc_hd__conb_1 _08225_ (.LO(_01771_));
 sky130_fd_sc_hd__conb_1 _08226_ (.LO(_01772_));
 sky130_fd_sc_hd__conb_1 _08227_ (.LO(_01773_));
 sky130_fd_sc_hd__conb_1 _08228_ (.LO(_01774_));
 sky130_fd_sc_hd__conb_1 _08229_ (.LO(_01775_));
 sky130_fd_sc_hd__conb_1 _08230_ (.LO(_01776_));
 sky130_fd_sc_hd__conb_1 _08231_ (.LO(_01777_));
 sky130_fd_sc_hd__conb_1 _08232_ (.LO(_01778_));
 sky130_fd_sc_hd__conb_1 _08233_ (.LO(_01779_));
 sky130_fd_sc_hd__conb_1 _08234_ (.LO(_01780_));
 sky130_fd_sc_hd__conb_1 _08235_ (.LO(_01781_));
 sky130_fd_sc_hd__conb_1 _08236_ (.LO(_01782_));
 sky130_fd_sc_hd__conb_1 _08237_ (.LO(_01783_));
 sky130_fd_sc_hd__conb_1 _08238_ (.LO(_01784_));
 sky130_fd_sc_hd__conb_1 _08239_ (.LO(_01785_));
 sky130_fd_sc_hd__conb_1 _08240_ (.LO(_01786_));
 sky130_fd_sc_hd__conb_1 _08241_ (.LO(_01787_));
 sky130_fd_sc_hd__conb_1 _08242_ (.LO(_01788_));
 sky130_fd_sc_hd__conb_1 _08243_ (.LO(_01789_));
 sky130_fd_sc_hd__conb_1 _08244_ (.LO(_01790_));
 sky130_fd_sc_hd__conb_1 _08245_ (.LO(_01791_));
 sky130_fd_sc_hd__conb_1 _08246_ (.LO(_01792_));
 sky130_fd_sc_hd__conb_1 _08247_ (.LO(_01793_));
 sky130_fd_sc_hd__conb_1 _08248_ (.LO(_01794_));
 sky130_fd_sc_hd__conb_1 _08249_ (.LO(_01795_));
 sky130_fd_sc_hd__conb_1 _08250_ (.LO(_01796_));
 sky130_fd_sc_hd__conb_1 _08251_ (.LO(_01797_));
 sky130_fd_sc_hd__conb_1 _08252_ (.LO(_01798_));
 sky130_fd_sc_hd__conb_1 _08253_ (.LO(_01799_));
 sky130_fd_sc_hd__conb_1 _08254_ (.LO(_01800_));
 sky130_fd_sc_hd__conb_1 _08255_ (.LO(_01801_));
 sky130_fd_sc_hd__conb_1 _08256_ (.LO(_01802_));
 sky130_fd_sc_hd__conb_1 _08257_ (.LO(_01803_));
 sky130_fd_sc_hd__conb_1 _08258_ (.LO(_01804_));
 sky130_fd_sc_hd__conb_1 _08259_ (.LO(_01805_));
 sky130_fd_sc_hd__conb_1 _08260_ (.LO(_01806_));
 sky130_fd_sc_hd__conb_1 _08261_ (.LO(_01807_));
 sky130_fd_sc_hd__conb_1 _08262_ (.LO(_01808_));
 sky130_fd_sc_hd__conb_1 _08263_ (.LO(_01809_));
 sky130_fd_sc_hd__conb_1 _08264_ (.LO(_01810_));
 sky130_fd_sc_hd__conb_1 _08265_ (.LO(_01811_));
 sky130_fd_sc_hd__conb_1 _08266_ (.LO(_01812_));
 sky130_fd_sc_hd__conb_1 _08267_ (.LO(_01813_));
 sky130_fd_sc_hd__conb_1 _08268_ (.LO(_01814_));
 sky130_fd_sc_hd__conb_1 _08269_ (.LO(_01815_));
 sky130_fd_sc_hd__conb_1 _08270_ (.LO(_01816_));
 sky130_fd_sc_hd__conb_1 _08271_ (.LO(_01817_));
 sky130_fd_sc_hd__conb_1 _08272_ (.LO(_01818_));
 sky130_fd_sc_hd__conb_1 _08273_ (.LO(_01819_));
 sky130_fd_sc_hd__conb_1 _08274_ (.LO(_01820_));
 sky130_fd_sc_hd__conb_1 _08275_ (.LO(_01821_));
 sky130_fd_sc_hd__conb_1 _08276_ (.LO(_01822_));
 sky130_fd_sc_hd__conb_1 _08277_ (.LO(_01823_));
 sky130_fd_sc_hd__conb_1 _08278_ (.LO(_01824_));
 sky130_fd_sc_hd__conb_1 _08279_ (.LO(_01825_));
 sky130_fd_sc_hd__conb_1 _08280_ (.LO(_01826_));
 sky130_fd_sc_hd__conb_1 _08281_ (.LO(_01827_));
 sky130_fd_sc_hd__conb_1 _08282_ (.LO(_01828_));
 sky130_fd_sc_hd__conb_1 _08283_ (.LO(_01829_));
 sky130_fd_sc_hd__conb_1 _08284_ (.LO(_01830_));
 sky130_fd_sc_hd__conb_1 _08285_ (.LO(_01831_));
 sky130_fd_sc_hd__conb_1 _08286_ (.LO(_01832_));
 sky130_fd_sc_hd__conb_1 _08287_ (.LO(_01833_));
 sky130_fd_sc_hd__conb_1 _08288_ (.LO(_01834_));
 sky130_fd_sc_hd__conb_1 _08289_ (.LO(_01835_));
 sky130_fd_sc_hd__conb_1 _08290_ (.LO(_01836_));
 sky130_fd_sc_hd__conb_1 _08291_ (.LO(_01837_));
 sky130_fd_sc_hd__conb_1 _08292_ (.LO(_01838_));
 sky130_fd_sc_hd__conb_1 _08293_ (.LO(_01839_));
 sky130_fd_sc_hd__conb_1 _08294_ (.LO(_01840_));
 sky130_fd_sc_hd__conb_1 _08295_ (.LO(_01841_));
 sky130_fd_sc_hd__conb_1 _08296_ (.LO(_01842_));
 sky130_fd_sc_hd__conb_1 _08297_ (.LO(_01843_));
 sky130_fd_sc_hd__conb_1 _08298_ (.LO(_01844_));
 sky130_fd_sc_hd__conb_1 _08299_ (.LO(_01845_));
 sky130_fd_sc_hd__conb_1 _08300_ (.LO(_01846_));
 sky130_fd_sc_hd__conb_1 _08301_ (.LO(_01847_));
 sky130_fd_sc_hd__conb_1 _08302_ (.LO(_01848_));
 sky130_fd_sc_hd__conb_1 _08303_ (.LO(_01849_));
 sky130_fd_sc_hd__conb_1 _08304_ (.LO(_01850_));
 sky130_fd_sc_hd__conb_1 _08305_ (.LO(_01851_));
 sky130_fd_sc_hd__conb_1 _08306_ (.LO(_01852_));
 sky130_fd_sc_hd__conb_1 _08307_ (.LO(_01853_));
 sky130_fd_sc_hd__conb_1 _08308_ (.LO(_01854_));
 sky130_fd_sc_hd__conb_1 _08309_ (.LO(_01855_));
 sky130_fd_sc_hd__conb_1 _08310_ (.LO(_01856_));
 sky130_fd_sc_hd__conb_1 _08311_ (.LO(_01857_));
 sky130_fd_sc_hd__conb_1 _08312_ (.LO(_01858_));
 sky130_fd_sc_hd__conb_1 _08313_ (.LO(_01859_));
 sky130_fd_sc_hd__conb_1 _08314_ (.LO(_01860_));
 sky130_fd_sc_hd__conb_1 _08315_ (.LO(_01861_));
 sky130_fd_sc_hd__conb_1 _08316_ (.LO(_01862_));
 sky130_fd_sc_hd__conb_1 _08317_ (.LO(_01863_));
 sky130_fd_sc_hd__conb_1 _08318_ (.LO(_01864_));
 sky130_fd_sc_hd__conb_1 _08319_ (.LO(_01865_));
 sky130_fd_sc_hd__conb_1 _08320_ (.LO(_01866_));
 sky130_fd_sc_hd__conb_1 _08321_ (.LO(_01867_));
 sky130_fd_sc_hd__conb_1 _08322_ (.LO(_01868_));
 sky130_fd_sc_hd__conb_1 _08323_ (.LO(_01869_));
 sky130_fd_sc_hd__conb_1 _08324_ (.LO(_01870_));
 sky130_fd_sc_hd__conb_1 _08325_ (.LO(_01871_));
 sky130_fd_sc_hd__conb_1 _08326_ (.LO(_01872_));
 sky130_fd_sc_hd__conb_1 _08327_ (.LO(_01873_));
 sky130_fd_sc_hd__conb_1 _08328_ (.LO(_01874_));
 sky130_fd_sc_hd__conb_1 _08329_ (.LO(_01875_));
 sky130_fd_sc_hd__conb_1 _08330_ (.LO(_01876_));
 sky130_fd_sc_hd__conb_1 _08331_ (.LO(_01877_));
 sky130_fd_sc_hd__conb_1 _08332_ (.LO(_01878_));
 sky130_fd_sc_hd__conb_1 _08333_ (.LO(_01879_));
 sky130_fd_sc_hd__conb_1 _08334_ (.LO(_01880_));
 sky130_fd_sc_hd__conb_1 _08335_ (.LO(_01881_));
 sky130_fd_sc_hd__conb_1 _08336_ (.LO(_01882_));
 sky130_fd_sc_hd__conb_1 _08337_ (.LO(_01883_));
 sky130_fd_sc_hd__conb_1 _08338_ (.LO(_01884_));
 sky130_fd_sc_hd__conb_1 _08339_ (.LO(_01885_));
 sky130_fd_sc_hd__conb_1 _08340_ (.LO(_01886_));
 sky130_fd_sc_hd__conb_1 _08341_ (.LO(_01887_));
 sky130_fd_sc_hd__conb_1 _08342_ (.LO(_01888_));
 sky130_fd_sc_hd__conb_1 _08343_ (.LO(_01889_));
 sky130_fd_sc_hd__conb_1 _08344_ (.LO(_01890_));
 sky130_fd_sc_hd__conb_1 _08345_ (.LO(_01891_));
 sky130_fd_sc_hd__conb_1 _08346_ (.LO(_01892_));
 sky130_fd_sc_hd__conb_1 _08347_ (.LO(_01893_));
 sky130_fd_sc_hd__conb_1 _08348_ (.LO(_01894_));
 sky130_fd_sc_hd__conb_1 _08349_ (.LO(_01895_));
 sky130_fd_sc_hd__conb_1 _08350_ (.LO(_01896_));
 sky130_fd_sc_hd__conb_1 _08351_ (.LO(_01897_));
 sky130_fd_sc_hd__conb_1 _08352_ (.LO(_01898_));
 sky130_fd_sc_hd__conb_1 _08353_ (.LO(_01899_));
 sky130_fd_sc_hd__conb_1 _08354_ (.LO(_01900_));
 sky130_fd_sc_hd__conb_1 _08355_ (.LO(_01901_));
 sky130_fd_sc_hd__conb_1 _08356_ (.LO(_01902_));
 sky130_fd_sc_hd__conb_1 _08357_ (.LO(_01903_));
 sky130_fd_sc_hd__conb_1 _08358_ (.LO(_01904_));
 sky130_fd_sc_hd__conb_1 _08359_ (.LO(_01905_));
 sky130_fd_sc_hd__conb_1 _08360_ (.LO(_01906_));
 sky130_fd_sc_hd__conb_1 _08361_ (.LO(_01907_));
 sky130_fd_sc_hd__conb_1 _08362_ (.LO(_01908_));
 sky130_fd_sc_hd__conb_1 _08363_ (.LO(_01909_));
 sky130_fd_sc_hd__conb_1 _08364_ (.LO(_01910_));
 sky130_fd_sc_hd__conb_1 _08365_ (.LO(_01911_));
 sky130_fd_sc_hd__conb_1 _08366_ (.LO(_01912_));
 sky130_fd_sc_hd__conb_1 _08367_ (.LO(_01913_));
 sky130_fd_sc_hd__conb_1 _08368_ (.LO(_01914_));
 sky130_fd_sc_hd__conb_1 _08369_ (.LO(_01915_));
 sky130_fd_sc_hd__conb_1 _08370_ (.LO(_01916_));
 sky130_fd_sc_hd__conb_1 _08371_ (.LO(_01917_));
 sky130_fd_sc_hd__conb_1 _08372_ (.LO(_01918_));
 sky130_fd_sc_hd__conb_1 _08373_ (.LO(_01919_));
 sky130_fd_sc_hd__conb_1 _08374_ (.LO(_01920_));
 sky130_fd_sc_hd__conb_1 _08375_ (.LO(_01921_));
 sky130_fd_sc_hd__conb_1 _08376_ (.LO(_01922_));
 sky130_fd_sc_hd__conb_1 _08377_ (.LO(_01923_));
 sky130_fd_sc_hd__conb_1 _08378_ (.LO(_01924_));
 sky130_fd_sc_hd__conb_1 _08379_ (.LO(_01925_));
 sky130_fd_sc_hd__conb_1 _08380_ (.LO(_01926_));
 sky130_fd_sc_hd__conb_1 _08381_ (.LO(_01927_));
 sky130_fd_sc_hd__conb_1 _08382_ (.LO(_01928_));
 sky130_fd_sc_hd__conb_1 _08383_ (.LO(_01929_));
 sky130_fd_sc_hd__conb_1 _08384_ (.LO(_01930_));
 sky130_fd_sc_hd__conb_1 _08385_ (.LO(_01931_));
 sky130_fd_sc_hd__conb_1 _08386_ (.LO(_01932_));
 sky130_fd_sc_hd__conb_1 _08387_ (.LO(_01933_));
 sky130_fd_sc_hd__conb_1 _08388_ (.LO(_01934_));
 sky130_fd_sc_hd__conb_1 _08389_ (.LO(_01935_));
 sky130_fd_sc_hd__conb_1 _08390_ (.LO(_01936_));
 sky130_fd_sc_hd__conb_1 _08391_ (.LO(_01937_));
 sky130_fd_sc_hd__conb_1 _08392_ (.LO(_01938_));
 sky130_fd_sc_hd__conb_1 _08393_ (.LO(_01939_));
 sky130_fd_sc_hd__conb_1 _08394_ (.LO(_01940_));
 sky130_fd_sc_hd__conb_1 _08395_ (.LO(_01941_));
 sky130_fd_sc_hd__conb_1 _08396_ (.LO(_01942_));
 sky130_fd_sc_hd__conb_1 _08397_ (.LO(_01943_));
 sky130_fd_sc_hd__conb_1 _08398_ (.LO(_01944_));
 sky130_fd_sc_hd__conb_1 _08399_ (.LO(_01945_));
 sky130_fd_sc_hd__conb_1 _08400_ (.LO(_01946_));
 sky130_fd_sc_hd__conb_1 _08401_ (.LO(_01947_));
 sky130_fd_sc_hd__conb_1 _08402_ (.LO(_01948_));
 sky130_fd_sc_hd__conb_1 _08403_ (.LO(_01949_));
 sky130_fd_sc_hd__conb_1 _08404_ (.LO(_01950_));
 sky130_fd_sc_hd__conb_1 _08405_ (.LO(_01951_));
 sky130_fd_sc_hd__conb_1 _08406_ (.LO(_01952_));
 sky130_fd_sc_hd__conb_1 _08407_ (.LO(_01953_));
 sky130_fd_sc_hd__conb_1 _08408_ (.LO(_01954_));
 sky130_fd_sc_hd__conb_1 _08409_ (.LO(_01955_));
 sky130_fd_sc_hd__conb_1 _08410_ (.LO(_01956_));
 sky130_fd_sc_hd__conb_1 _08411_ (.LO(_01957_));
 sky130_fd_sc_hd__conb_1 _08412_ (.LO(_01958_));
 sky130_fd_sc_hd__conb_1 _08413_ (.LO(_01959_));
 sky130_fd_sc_hd__conb_1 _08414_ (.LO(_01960_));
 sky130_fd_sc_hd__conb_1 _08415_ (.LO(_01961_));
 sky130_fd_sc_hd__conb_1 _08416_ (.LO(_01962_));
 sky130_fd_sc_hd__conb_1 _08417_ (.LO(_01963_));
 sky130_fd_sc_hd__conb_1 _08418_ (.LO(_01964_));
 sky130_fd_sc_hd__conb_1 _08419_ (.LO(_01965_));
 sky130_fd_sc_hd__conb_1 _08420_ (.LO(_01966_));
 sky130_fd_sc_hd__conb_1 _08421_ (.LO(_01967_));
 sky130_fd_sc_hd__conb_1 _08422_ (.LO(_01968_));
 sky130_fd_sc_hd__conb_1 _08423_ (.LO(_01969_));
 sky130_fd_sc_hd__conb_1 _08424_ (.LO(_01970_));
 sky130_fd_sc_hd__conb_1 _08425_ (.LO(_01971_));
 sky130_fd_sc_hd__conb_1 _08426_ (.LO(_01972_));
 sky130_fd_sc_hd__conb_1 _08427_ (.LO(_01973_));
 sky130_fd_sc_hd__conb_1 _08428_ (.LO(_01974_));
 sky130_fd_sc_hd__conb_1 _08429_ (.LO(_01975_));
 sky130_fd_sc_hd__conb_1 _08430_ (.LO(_01976_));
 sky130_fd_sc_hd__conb_1 _08431_ (.LO(_01977_));
 sky130_fd_sc_hd__conb_1 _08432_ (.LO(_01978_));
 sky130_fd_sc_hd__conb_1 _08433_ (.LO(_01979_));
 sky130_fd_sc_hd__conb_1 _08434_ (.LO(_01980_));
 sky130_fd_sc_hd__conb_1 _08435_ (.LO(_01981_));
 sky130_fd_sc_hd__conb_1 _08436_ (.LO(_01982_));
 sky130_fd_sc_hd__conb_1 _08437_ (.LO(_01983_));
 sky130_fd_sc_hd__conb_1 _08438_ (.LO(_01984_));
 sky130_fd_sc_hd__conb_1 _08439_ (.LO(_01985_));
 sky130_fd_sc_hd__conb_1 _08440_ (.LO(_01986_));
 sky130_fd_sc_hd__conb_1 _08441_ (.LO(_01987_));
 sky130_fd_sc_hd__conb_1 _08442_ (.LO(_01988_));
 sky130_fd_sc_hd__conb_1 _08443_ (.LO(_01989_));
 sky130_fd_sc_hd__conb_1 _08444_ (.LO(_01990_));
 sky130_fd_sc_hd__conb_1 _08445_ (.LO(_01991_));
 sky130_fd_sc_hd__conb_1 _08446_ (.LO(_01992_));
 sky130_fd_sc_hd__conb_1 _08447_ (.LO(_01993_));
 sky130_fd_sc_hd__conb_1 _08448_ (.LO(_01994_));
 sky130_fd_sc_hd__conb_1 _08449_ (.LO(_01995_));
 sky130_fd_sc_hd__conb_1 _08450_ (.LO(_01996_));
 sky130_fd_sc_hd__conb_1 _08451_ (.LO(_01997_));
 sky130_fd_sc_hd__conb_1 _08452_ (.LO(_01998_));
 sky130_fd_sc_hd__conb_1 _08453_ (.LO(_01999_));
 sky130_fd_sc_hd__conb_1 _08454_ (.LO(_02000_));
 sky130_fd_sc_hd__conb_1 _08455_ (.LO(_02001_));
 sky130_fd_sc_hd__conb_1 _08456_ (.LO(_02002_));
 sky130_fd_sc_hd__conb_1 _08457_ (.LO(_02003_));
 sky130_fd_sc_hd__conb_1 _08458_ (.LO(_02004_));
 sky130_fd_sc_hd__conb_1 _08459_ (.LO(_02005_));
 sky130_fd_sc_hd__conb_1 _08460_ (.LO(_02006_));
 sky130_fd_sc_hd__conb_1 _08461_ (.LO(_02007_));
 sky130_fd_sc_hd__conb_1 _08462_ (.LO(_02008_));
 sky130_fd_sc_hd__conb_1 _08463_ (.LO(_02009_));
 sky130_fd_sc_hd__conb_1 _08464_ (.LO(_02010_));
 sky130_fd_sc_hd__conb_1 _08465_ (.LO(_02011_));
 sky130_fd_sc_hd__conb_1 _08466_ (.LO(_02012_));
 sky130_fd_sc_hd__conb_1 _08467_ (.LO(_02013_));
 sky130_fd_sc_hd__conb_1 _08468_ (.LO(_02014_));
 sky130_fd_sc_hd__conb_1 _08469_ (.LO(_02015_));
 sky130_fd_sc_hd__conb_1 _08470_ (.LO(_02016_));
 sky130_fd_sc_hd__conb_1 _08471_ (.LO(_02017_));
 sky130_fd_sc_hd__conb_1 _08472_ (.LO(_02018_));
 sky130_fd_sc_hd__conb_1 _08473_ (.LO(_02019_));
 sky130_fd_sc_hd__conb_1 _08474_ (.LO(_02020_));
 sky130_fd_sc_hd__conb_1 _08475_ (.LO(_02021_));
 sky130_fd_sc_hd__conb_1 _08476_ (.LO(_02022_));
 sky130_fd_sc_hd__buf_2 _08477_ (.A(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ),
    .X(cb_east_out[0]));
 sky130_fd_sc_hd__buf_2 _08478_ (.A(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ),
    .X(cb_east_out[1]));
 sky130_fd_sc_hd__buf_2 _08479_ (.A(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ),
    .X(cb_east_out[2]));
 sky130_fd_sc_hd__buf_2 _08480_ (.A(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ),
    .X(cb_east_out[3]));
 sky130_fd_sc_hd__buf_2 _08481_ (.A(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ),
    .X(cb_east_out[4]));
 sky130_fd_sc_hd__buf_2 _08482_ (.A(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ),
    .X(cb_east_out[5]));
 sky130_fd_sc_hd__buf_2 _08483_ (.A(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ),
    .X(cb_east_out[6]));
 sky130_fd_sc_hd__buf_2 _08484_ (.A(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ),
    .X(cb_east_out[7]));
 sky130_fd_sc_hd__buf_2 _08485_ (.A(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ),
    .X(cb_east_out[8]));
 sky130_fd_sc_hd__buf_2 _08486_ (.A(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ),
    .X(cb_east_out[9]));
 sky130_fd_sc_hd__buf_2 _08487_ (.A(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ),
    .X(cb_north_out[0]));
 sky130_fd_sc_hd__buf_2 _08488_ (.A(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ),
    .X(cb_north_out[1]));
 sky130_fd_sc_hd__buf_2 _08489_ (.A(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ),
    .X(cb_north_out[2]));
 sky130_fd_sc_hd__buf_2 _08490_ (.A(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ),
    .X(cb_north_out[3]));
 sky130_fd_sc_hd__buf_2 _08491_ (.A(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ),
    .X(cb_north_out[4]));
 sky130_fd_sc_hd__buf_2 _08492_ (.A(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ),
    .X(cb_north_out[5]));
 sky130_fd_sc_hd__buf_2 _08493_ (.A(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ),
    .X(cb_north_out[6]));
 sky130_fd_sc_hd__buf_2 _08494_ (.A(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ),
    .X(cb_north_out[7]));
 sky130_fd_sc_hd__buf_2 _08495_ (.A(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ),
    .X(cb_north_out[8]));
 sky130_fd_sc_hd__buf_2 _08496_ (.A(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ),
    .X(cb_north_out[9]));
 sky130_fd_sc_hd__buf_2 _08497_ (.A(set_out_hard),
    .X(clb_south_out[4]));
 sky130_fd_sc_hd__buf_2 _08498_ (.A(shift_out_hard),
    .X(clb_west_out[4]));
 sky130_fd_sc_hd__buf_2 _08499_ (.A(north_double[4]),
    .X(south_double[0]));
 sky130_fd_sc_hd__buf_2 _08500_ (.A(north_double[5]),
    .X(south_double[1]));
 sky130_fd_sc_hd__buf_2 _08501_ (.A(north_double[6]),
    .X(south_double[2]));
 sky130_fd_sc_hd__buf_2 _08502_ (.A(north_double[7]),
    .X(south_double[3]));
 sky130_fd_sc_hd__buf_2 _08503_ (.A(east_double[0]),
    .X(west_double[4]));
 sky130_fd_sc_hd__buf_2 _08504_ (.A(east_double[1]),
    .X(west_double[5]));
 sky130_fd_sc_hd__buf_2 _08505_ (.A(east_double[2]),
    .X(west_double[6]));
 sky130_fd_sc_hd__buf_2 _08506_ (.A(east_double[3]),
    .X(west_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08507_ (.A(north_double[5]),
    .TE_B(_00687_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08508_ (.A(north_double[4]),
    .TE_B(_00688_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08509_ (.A(south_single[3]),
    .TE_B(_00689_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08510_ (.A(south_single[2]),
    .TE_B(_00690_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08511_ (.A(south_single[1]),
    .TE_B(_00691_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08512_ (.A(south_single[0]),
    .TE_B(_00692_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08513_ (.A(shift_out_hard),
    .TE_B(_00693_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08514_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00694_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08515_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00695_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08516_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00696_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08517_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00697_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08518_ (.A(south_double[7]),
    .TE_B(_00698_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08519_ (.A(south_double[6]),
    .TE_B(_00699_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08520_ (.A(south_double[5]),
    .TE_B(_00700_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08521_ (.A(south_double[4]),
    .TE_B(_00701_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08522_ (.A(north_double[7]),
    .TE_B(_00702_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08523_ (.A(north_double[6]),
    .TE_B(_00703_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08524_ (.A(north_double[5]),
    .TE_B(_00704_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08525_ (.A(north_double[4]),
    .TE_B(_00705_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08526_ (.A(south_single[3]),
    .TE_B(_00706_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08527_ (.A(south_single[2]),
    .TE_B(_00707_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08528_ (.A(south_single[1]),
    .TE_B(_00708_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08529_ (.A(south_single[0]),
    .TE_B(_00709_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08530_ (.A(shift_out_hard),
    .TE_B(_00710_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08531_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00711_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08532_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00712_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08533_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00713_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08534_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00714_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08535_ (.A(south_double[7]),
    .TE_B(_00715_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08536_ (.A(south_double[6]),
    .TE_B(_00716_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08537_ (.A(south_double[5]),
    .TE_B(_00717_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08538_ (.A(south_double[4]),
    .TE_B(_00718_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08539_ (.A(north_double[7]),
    .TE_B(_00719_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08540_ (.A(north_double[6]),
    .TE_B(_00720_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08541_ (.A(north_double[5]),
    .TE_B(_00721_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08542_ (.A(north_double[4]),
    .TE_B(_00722_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08543_ (.A(south_single[3]),
    .TE_B(_00723_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08544_ (.A(south_single[2]),
    .TE_B(_00724_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08545_ (.A(south_single[1]),
    .TE_B(_00725_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08546_ (.A(south_single[0]),
    .TE_B(_00726_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08547_ (.A(shift_out_hard),
    .TE_B(_00727_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08548_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00728_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08549_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00729_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08550_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00730_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08551_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00731_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08552_ (.A(south_double[7]),
    .TE_B(_00732_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08553_ (.A(south_double[6]),
    .TE_B(_00733_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08554_ (.A(south_double[5]),
    .TE_B(_00734_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08555_ (.A(south_double[4]),
    .TE_B(_00735_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08556_ (.A(north_double[7]),
    .TE_B(_00736_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08557_ (.A(north_double[6]),
    .TE_B(_00737_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08558_ (.A(north_double[5]),
    .TE_B(_00738_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08559_ (.A(north_double[4]),
    .TE_B(_00739_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08560_ (.A(south_single[3]),
    .TE_B(_00740_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08561_ (.A(south_single[2]),
    .TE_B(_00741_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08562_ (.A(south_single[1]),
    .TE_B(_00742_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08563_ (.A(south_single[0]),
    .TE_B(_00743_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08564_ (.A(shift_out_hard),
    .TE_B(_00744_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08565_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00745_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08566_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00746_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08567_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00747_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08568_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00748_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08569_ (.A(south_double[7]),
    .TE_B(_00749_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08570_ (.A(south_double[6]),
    .TE_B(_00750_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08571_ (.A(south_double[5]),
    .TE_B(_00751_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08572_ (.A(south_double[4]),
    .TE_B(_00752_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08573_ (.A(north_double[7]),
    .TE_B(_00753_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08574_ (.A(north_double[6]),
    .TE_B(_00754_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08575_ (.A(north_double[5]),
    .TE_B(_00755_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08576_ (.A(north_double[4]),
    .TE_B(_00756_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08577_ (.A(south_single[3]),
    .TE_B(_00757_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08578_ (.A(south_single[2]),
    .TE_B(_00758_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08579_ (.A(south_single[1]),
    .TE_B(_00759_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08580_ (.A(south_single[0]),
    .TE_B(_00760_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08581_ (.A(shift_out_hard),
    .TE_B(_00761_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08582_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00762_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08583_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00763_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08584_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00764_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08585_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00765_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08586_ (.A(south_double[7]),
    .TE_B(_00766_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08587_ (.A(south_double[6]),
    .TE_B(_00767_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08588_ (.A(south_double[5]),
    .TE_B(_00768_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08589_ (.A(south_double[4]),
    .TE_B(_00769_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08590_ (.A(north_double[7]),
    .TE_B(_00770_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08591_ (.A(north_double[6]),
    .TE_B(_00771_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08592_ (.A(north_double[5]),
    .TE_B(_00772_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08593_ (.A(north_double[4]),
    .TE_B(_00773_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08594_ (.A(south_single[3]),
    .TE_B(_00774_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08595_ (.A(south_single[2]),
    .TE_B(_00775_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08596_ (.A(south_single[1]),
    .TE_B(_00776_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08597_ (.A(south_single[0]),
    .TE_B(_00777_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08598_ (.A(shift_out_hard),
    .TE_B(_00778_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08599_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00779_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08600_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00780_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08601_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00781_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08602_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00782_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08603_ (.A(south_double[7]),
    .TE_B(_00783_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08604_ (.A(south_double[6]),
    .TE_B(_00784_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08605_ (.A(south_double[5]),
    .TE_B(_00785_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08606_ (.A(south_double[4]),
    .TE_B(_00786_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08607_ (.A(north_double[7]),
    .TE_B(_00787_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08608_ (.A(north_double[6]),
    .TE_B(_00788_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08609_ (.A(north_double[5]),
    .TE_B(_00789_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08610_ (.A(north_double[4]),
    .TE_B(_00790_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08611_ (.A(south_single[3]),
    .TE_B(_00791_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08612_ (.A(south_single[2]),
    .TE_B(_00792_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08613_ (.A(south_single[1]),
    .TE_B(_00793_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08614_ (.A(south_single[0]),
    .TE_B(_00794_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08615_ (.A(shift_out_hard),
    .TE_B(_00795_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08616_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00796_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08617_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00797_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08618_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00798_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08619_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00799_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08620_ (.A(south_double[7]),
    .TE_B(_00800_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08621_ (.A(south_double[6]),
    .TE_B(_00801_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08622_ (.A(south_double[5]),
    .TE_B(_00802_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08623_ (.A(south_double[4]),
    .TE_B(_00803_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08624_ (.A(north_double[7]),
    .TE_B(_00804_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08625_ (.A(north_double[6]),
    .TE_B(_00805_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08626_ (.A(north_double[5]),
    .TE_B(_00806_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08627_ (.A(north_double[4]),
    .TE_B(_00807_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08628_ (.A(south_single[3]),
    .TE_B(_00808_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08629_ (.A(south_single[2]),
    .TE_B(_00809_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08630_ (.A(south_single[1]),
    .TE_B(_00810_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08631_ (.A(south_single[0]),
    .TE_B(_00811_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08632_ (.A(shift_out_hard),
    .TE_B(_00611_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08633_ (.A(shift_out_hard),
    .TE_B(_00617_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _08634_ (.A(shift_out_hard),
    .TE_B(_00623_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _08635_ (.A(shift_out_hard),
    .TE_B(_00629_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _08636_ (.A(shift_out_hard),
    .TE_B(_00635_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08637_ (.A(shift_out_hard),
    .TE_B(_00641_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08638_ (.A(shift_out_hard),
    .TE_B(_00647_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08639_ (.A(shift_out_hard),
    .TE_B(_00653_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08640_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00612_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08641_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00618_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _08642_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00624_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _08643_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00630_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _08644_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00636_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08645_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00642_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08646_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00648_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08647_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00654_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08648_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00613_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08649_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00619_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _08650_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00625_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _08651_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00631_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _08652_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00637_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08653_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00643_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08654_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00649_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08655_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00655_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08656_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00614_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08657_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00620_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _08658_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00626_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _08659_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00632_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _08660_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00638_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08661_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00644_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08662_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00650_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08663_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00656_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08664_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00615_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _08665_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00621_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _08666_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00627_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _08667_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00633_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _08668_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00639_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08669_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00645_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08670_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00651_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08671_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00657_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08672_ (.A(cb_east_in[4]),
    .TE_B(_00812_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08673_ (.A(cb_east_in[3]),
    .TE_B(_00813_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08674_ (.A(cb_east_in[2]),
    .TE_B(_00814_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08675_ (.A(cb_east_in[1]),
    .TE_B(_00815_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08676_ (.A(cb_east_in[0]),
    .TE_B(_00816_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08677_ (.A(south_double[7]),
    .TE_B(_00817_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08678_ (.A(south_double[6]),
    .TE_B(_00818_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08679_ (.A(south_double[5]),
    .TE_B(_00819_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08680_ (.A(south_double[4]),
    .TE_B(_00820_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08681_ (.A(north_double[7]),
    .TE_B(_00821_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08682_ (.A(north_double[6]),
    .TE_B(_00822_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08683_ (.A(north_double[5]),
    .TE_B(_00823_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08684_ (.A(north_double[4]),
    .TE_B(_00824_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08685_ (.A(south_single[3]),
    .TE_B(_00825_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08686_ (.A(south_single[2]),
    .TE_B(_00826_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08687_ (.A(south_single[1]),
    .TE_B(_00827_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08688_ (.A(south_single[0]),
    .TE_B(_00828_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08689_ (.A(cb_east_in[4]),
    .TE_B(_00829_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08690_ (.A(cb_east_in[3]),
    .TE_B(_00830_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08691_ (.A(cb_east_in[2]),
    .TE_B(_00831_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08692_ (.A(cb_east_in[1]),
    .TE_B(_00832_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08693_ (.A(cb_east_in[0]),
    .TE_B(_00833_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08694_ (.A(south_double[7]),
    .TE_B(_00834_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08695_ (.A(south_double[6]),
    .TE_B(_00835_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08696_ (.A(south_double[5]),
    .TE_B(_00836_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08697_ (.A(south_double[4]),
    .TE_B(_00837_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08698_ (.A(north_double[7]),
    .TE_B(_00838_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08699_ (.A(north_double[6]),
    .TE_B(_00839_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08700_ (.A(north_double[5]),
    .TE_B(_00840_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08701_ (.A(north_double[4]),
    .TE_B(_00841_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08702_ (.A(south_single[3]),
    .TE_B(_00842_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08703_ (.A(south_single[2]),
    .TE_B(_00843_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08704_ (.A(south_single[1]),
    .TE_B(_00844_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08705_ (.A(south_single[0]),
    .TE_B(_00845_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08706_ (.A(cb_east_in[4]),
    .TE_B(_00846_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08707_ (.A(cb_east_in[3]),
    .TE_B(_00847_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08708_ (.A(cb_east_in[2]),
    .TE_B(_00848_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08709_ (.A(cb_east_in[1]),
    .TE_B(_00849_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08710_ (.A(cb_east_in[0]),
    .TE_B(_00850_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08711_ (.A(south_double[7]),
    .TE_B(_00851_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08712_ (.A(south_double[6]),
    .TE_B(_00852_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08713_ (.A(south_double[5]),
    .TE_B(_00853_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08714_ (.A(south_double[4]),
    .TE_B(_00854_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08715_ (.A(north_double[7]),
    .TE_B(_00855_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08716_ (.A(north_double[6]),
    .TE_B(_00856_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08717_ (.A(north_double[5]),
    .TE_B(_00857_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08718_ (.A(north_double[4]),
    .TE_B(_00858_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08719_ (.A(south_single[3]),
    .TE_B(_00859_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08720_ (.A(south_single[2]),
    .TE_B(_00860_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08721_ (.A(south_single[1]),
    .TE_B(_00861_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08722_ (.A(south_single[0]),
    .TE_B(_00862_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08723_ (.A(cb_east_in[4]),
    .TE_B(_00863_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08724_ (.A(cb_east_in[3]),
    .TE_B(_00864_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08725_ (.A(cb_east_in[2]),
    .TE_B(_00865_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08726_ (.A(cb_east_in[1]),
    .TE_B(_00866_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08727_ (.A(cb_east_in[0]),
    .TE_B(_00867_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08728_ (.A(south_double[7]),
    .TE_B(_00868_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08729_ (.A(south_double[6]),
    .TE_B(_00869_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08730_ (.A(south_double[5]),
    .TE_B(_00870_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08731_ (.A(south_double[4]),
    .TE_B(_00871_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08732_ (.A(north_double[7]),
    .TE_B(_00872_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08733_ (.A(north_double[6]),
    .TE_B(_00873_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08734_ (.A(north_double[5]),
    .TE_B(_00874_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08735_ (.A(north_double[4]),
    .TE_B(_00875_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08736_ (.A(south_single[3]),
    .TE_B(_00876_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08737_ (.A(south_single[2]),
    .TE_B(_00877_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08738_ (.A(south_single[1]),
    .TE_B(_00878_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08739_ (.A(south_single[0]),
    .TE_B(_00879_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08740_ (.A(cb_east_in[4]),
    .TE_B(_00880_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08741_ (.A(cb_east_in[3]),
    .TE_B(_00881_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08742_ (.A(cb_east_in[2]),
    .TE_B(_00882_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08743_ (.A(cb_east_in[1]),
    .TE_B(_00883_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08744_ (.A(cb_east_in[0]),
    .TE_B(_00884_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08745_ (.A(south_double[7]),
    .TE_B(_00885_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08746_ (.A(south_double[6]),
    .TE_B(_00886_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08747_ (.A(south_double[5]),
    .TE_B(_00887_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08748_ (.A(south_double[4]),
    .TE_B(_00888_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08749_ (.A(north_double[7]),
    .TE_B(_00889_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08750_ (.A(north_double[6]),
    .TE_B(_00890_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08751_ (.A(north_double[5]),
    .TE_B(_00891_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08752_ (.A(north_double[4]),
    .TE_B(_00892_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08753_ (.A(south_single[3]),
    .TE_B(_00893_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08754_ (.A(south_single[2]),
    .TE_B(_00894_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08755_ (.A(south_single[1]),
    .TE_B(_00895_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08756_ (.A(south_single[0]),
    .TE_B(_00896_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08757_ (.A(cb_east_in[4]),
    .TE_B(_00897_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08758_ (.A(cb_east_in[3]),
    .TE_B(_00898_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08759_ (.A(cb_east_in[2]),
    .TE_B(_00899_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08760_ (.A(cb_east_in[1]),
    .TE_B(_00900_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08761_ (.A(cb_east_in[0]),
    .TE_B(_00901_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08762_ (.A(south_double[7]),
    .TE_B(_00902_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08763_ (.A(south_double[6]),
    .TE_B(_00903_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08764_ (.A(south_double[5]),
    .TE_B(_00904_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08765_ (.A(south_double[4]),
    .TE_B(_00905_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08766_ (.A(north_double[7]),
    .TE_B(_00906_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08767_ (.A(north_double[6]),
    .TE_B(_00907_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08768_ (.A(north_double[5]),
    .TE_B(_00908_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08769_ (.A(north_double[4]),
    .TE_B(_00909_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08770_ (.A(south_single[3]),
    .TE_B(_00910_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08771_ (.A(south_single[2]),
    .TE_B(_00911_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08772_ (.A(south_single[1]),
    .TE_B(_00912_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08773_ (.A(south_single[0]),
    .TE_B(_00913_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08774_ (.A(cb_east_in[4]),
    .TE_B(_00914_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08775_ (.A(cb_east_in[3]),
    .TE_B(_00915_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08776_ (.A(cb_east_in[2]),
    .TE_B(_00916_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08777_ (.A(cb_east_in[1]),
    .TE_B(_00917_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08778_ (.A(cb_east_in[0]),
    .TE_B(_00918_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08779_ (.A(south_double[7]),
    .TE_B(_00919_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08780_ (.A(south_double[6]),
    .TE_B(_00920_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08781_ (.A(south_double[5]),
    .TE_B(_00921_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08782_ (.A(south_double[4]),
    .TE_B(_00922_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08783_ (.A(north_double[7]),
    .TE_B(_00923_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08784_ (.A(north_double[6]),
    .TE_B(_00924_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08785_ (.A(north_double[5]),
    .TE_B(_00925_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08786_ (.A(north_double[4]),
    .TE_B(_00926_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08787_ (.A(south_single[3]),
    .TE_B(_00927_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08788_ (.A(south_single[2]),
    .TE_B(_00928_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08789_ (.A(south_single[1]),
    .TE_B(_00929_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08790_ (.A(south_single[0]),
    .TE_B(_00930_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08791_ (.A(cb_east_in[4]),
    .TE_B(_00931_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08792_ (.A(cb_east_in[3]),
    .TE_B(_00932_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08793_ (.A(cb_east_in[2]),
    .TE_B(_00933_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08794_ (.A(cb_east_in[1]),
    .TE_B(_00934_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08795_ (.A(cb_east_in[0]),
    .TE_B(_00935_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08796_ (.A(south_double[7]),
    .TE_B(_00936_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08797_ (.A(south_double[6]),
    .TE_B(_00937_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08798_ (.A(south_double[5]),
    .TE_B(_00938_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08799_ (.A(south_double[4]),
    .TE_B(_00939_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08800_ (.A(north_double[7]),
    .TE_B(_00940_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08801_ (.A(north_double[6]),
    .TE_B(_00941_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08802_ (.A(north_double[5]),
    .TE_B(_00942_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08803_ (.A(north_double[4]),
    .TE_B(_00943_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08804_ (.A(south_single[3]),
    .TE_B(_00944_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08805_ (.A(south_single[2]),
    .TE_B(_00945_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08806_ (.A(south_single[1]),
    .TE_B(_00946_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08807_ (.A(south_single[0]),
    .TE_B(_00947_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08808_ (.A(cb_east_in[4]),
    .TE_B(_00948_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08809_ (.A(cb_east_in[3]),
    .TE_B(_00949_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08810_ (.A(cb_east_in[2]),
    .TE_B(_00950_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08811_ (.A(cb_east_in[1]),
    .TE_B(_00951_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08812_ (.A(cb_east_in[0]),
    .TE_B(_00952_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08813_ (.A(south_double[7]),
    .TE_B(_00953_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08814_ (.A(south_double[6]),
    .TE_B(_00954_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08815_ (.A(south_double[5]),
    .TE_B(_00955_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08816_ (.A(south_double[4]),
    .TE_B(_00956_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08817_ (.A(north_double[7]),
    .TE_B(_00957_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08818_ (.A(north_double[6]),
    .TE_B(_00958_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08819_ (.A(north_double[5]),
    .TE_B(_00959_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08820_ (.A(north_double[4]),
    .TE_B(_00960_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08821_ (.A(south_single[3]),
    .TE_B(_00961_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08822_ (.A(south_single[2]),
    .TE_B(_00962_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08823_ (.A(south_single[1]),
    .TE_B(_00963_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08824_ (.A(south_single[0]),
    .TE_B(_00964_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08825_ (.A(cb_east_in[4]),
    .TE_B(_00965_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08826_ (.A(cb_east_in[3]),
    .TE_B(_00966_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08827_ (.A(cb_east_in[2]),
    .TE_B(_00967_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08828_ (.A(cb_east_in[1]),
    .TE_B(_00968_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08829_ (.A(cb_east_in[0]),
    .TE_B(_00969_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08830_ (.A(south_double[7]),
    .TE_B(_00970_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08831_ (.A(south_double[6]),
    .TE_B(_00971_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08832_ (.A(south_double[5]),
    .TE_B(_00972_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08833_ (.A(south_double[4]),
    .TE_B(_00973_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08834_ (.A(north_double[7]),
    .TE_B(_00974_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08835_ (.A(north_double[6]),
    .TE_B(_00975_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08836_ (.A(north_double[5]),
    .TE_B(_00976_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08837_ (.A(north_double[4]),
    .TE_B(_00977_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08838_ (.A(south_single[3]),
    .TE_B(_00978_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08839_ (.A(south_single[2]),
    .TE_B(_00979_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08840_ (.A(south_single[1]),
    .TE_B(_00980_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08841_ (.A(south_single[0]),
    .TE_B(_00981_),
    .Z(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08842_ (.A(cb_north_in[4]),
    .TE_B(_00142_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _08843_ (.A(cb_north_in[4]),
    .TE_B(_00143_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _08844_ (.A(cb_north_in[4]),
    .TE_B(_00144_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _08845_ (.A(cb_north_in[4]),
    .TE_B(_00145_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _08846_ (.A(cb_north_in[4]),
    .TE_B(_00146_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08847_ (.A(cb_north_in[4]),
    .TE_B(_00147_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08848_ (.A(cb_north_in[4]),
    .TE_B(_00148_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08849_ (.A(cb_north_in[4]),
    .TE_B(_00149_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08850_ (.A(cb_north_in[3]),
    .TE_B(_00150_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _08851_ (.A(cb_north_in[3]),
    .TE_B(_00151_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _08852_ (.A(cb_north_in[3]),
    .TE_B(_00152_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _08853_ (.A(cb_north_in[3]),
    .TE_B(_00153_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _08854_ (.A(cb_north_in[3]),
    .TE_B(_00154_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08855_ (.A(cb_north_in[3]),
    .TE_B(_00155_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08856_ (.A(cb_north_in[3]),
    .TE_B(_00156_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08857_ (.A(cb_north_in[3]),
    .TE_B(_00157_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08858_ (.A(cb_north_in[2]),
    .TE_B(_00158_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _08859_ (.A(cb_north_in[2]),
    .TE_B(_00159_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _08860_ (.A(cb_north_in[2]),
    .TE_B(_00160_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _08861_ (.A(cb_north_in[2]),
    .TE_B(_00161_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _08862_ (.A(cb_north_in[2]),
    .TE_B(_00162_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08863_ (.A(cb_north_in[2]),
    .TE_B(_00163_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08864_ (.A(cb_north_in[2]),
    .TE_B(_00164_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08865_ (.A(cb_north_in[2]),
    .TE_B(_00165_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08866_ (.A(cb_north_in[1]),
    .TE_B(_00166_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _08867_ (.A(cb_north_in[1]),
    .TE_B(_00167_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _08868_ (.A(cb_north_in[1]),
    .TE_B(_00168_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _08869_ (.A(cb_north_in[1]),
    .TE_B(_00169_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _08870_ (.A(cb_north_in[1]),
    .TE_B(_00170_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08871_ (.A(cb_north_in[1]),
    .TE_B(_00171_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08872_ (.A(cb_north_in[1]),
    .TE_B(_00172_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08873_ (.A(cb_north_in[1]),
    .TE_B(_00173_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08874_ (.A(cb_north_in[0]),
    .TE_B(_00174_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _08875_ (.A(cb_north_in[0]),
    .TE_B(_00175_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _08876_ (.A(cb_north_in[0]),
    .TE_B(_00176_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _08877_ (.A(cb_north_in[0]),
    .TE_B(_00177_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _08878_ (.A(cb_north_in[0]),
    .TE_B(_00178_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _08879_ (.A(cb_north_in[0]),
    .TE_B(_00179_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _08880_ (.A(cb_north_in[0]),
    .TE_B(_00180_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _08881_ (.A(cb_north_in[0]),
    .TE_B(_00181_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _08882_ (.A(set_out_hard),
    .TE_B(_00182_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08883_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00183_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08884_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00184_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08885_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00185_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08886_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00186_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08887_ (.A(east_double[3]),
    .TE_B(_00187_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08888_ (.A(east_double[2]),
    .TE_B(_00188_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08889_ (.A(east_double[1]),
    .TE_B(_00189_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08890_ (.A(east_double[0]),
    .TE_B(_00190_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08891_ (.A(west_double[3]),
    .TE_B(_00196_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08892_ (.A(west_double[2]),
    .TE_B(_00202_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08893_ (.A(west_double[1]),
    .TE_B(_00208_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08894_ (.A(west_double[0]),
    .TE_B(_00214_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08895_ (.A(west_single[3]),
    .TE_B(_00220_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08896_ (.A(west_single[2]),
    .TE_B(_00226_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08897_ (.A(west_single[1]),
    .TE_B(_00232_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08898_ (.A(west_single[0]),
    .TE_B(_00238_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08899_ (.A(set_out_hard),
    .TE_B(_00239_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08900_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00240_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08901_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00241_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08902_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00242_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08903_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00243_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08904_ (.A(east_double[3]),
    .TE_B(_00244_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08905_ (.A(east_double[2]),
    .TE_B(_00245_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08906_ (.A(east_double[1]),
    .TE_B(_00246_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08907_ (.A(east_double[0]),
    .TE_B(_00247_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08908_ (.A(west_double[3]),
    .TE_B(_00248_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08909_ (.A(west_double[2]),
    .TE_B(_00249_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08910_ (.A(west_double[1]),
    .TE_B(_00250_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08911_ (.A(west_double[0]),
    .TE_B(_00251_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08912_ (.A(west_single[3]),
    .TE_B(_00252_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08913_ (.A(west_single[2]),
    .TE_B(_00253_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08914_ (.A(west_single[1]),
    .TE_B(_00254_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08915_ (.A(west_single[0]),
    .TE_B(_00255_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08916_ (.A(set_out_hard),
    .TE_B(_00256_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08917_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00257_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08918_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00258_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08919_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00259_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08920_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00260_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08921_ (.A(east_double[3]),
    .TE_B(_00261_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08922_ (.A(east_double[2]),
    .TE_B(_00262_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08923_ (.A(east_double[1]),
    .TE_B(_00263_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08924_ (.A(east_double[0]),
    .TE_B(_00264_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08925_ (.A(west_double[3]),
    .TE_B(_00265_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08926_ (.A(west_double[2]),
    .TE_B(_00266_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08927_ (.A(west_double[1]),
    .TE_B(_00267_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08928_ (.A(west_double[0]),
    .TE_B(_00268_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08929_ (.A(west_single[3]),
    .TE_B(_00269_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08930_ (.A(west_single[2]),
    .TE_B(_00270_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08931_ (.A(west_single[1]),
    .TE_B(_00271_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08932_ (.A(west_single[0]),
    .TE_B(_00272_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08933_ (.A(set_out_hard),
    .TE_B(_00273_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08934_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00274_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08935_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00275_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08936_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00276_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08937_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00277_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08938_ (.A(east_double[3]),
    .TE_B(_00278_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08939_ (.A(east_double[2]),
    .TE_B(_00279_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08940_ (.A(east_double[1]),
    .TE_B(_00280_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08941_ (.A(east_double[0]),
    .TE_B(_00281_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08942_ (.A(west_double[3]),
    .TE_B(_00282_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08943_ (.A(west_double[2]),
    .TE_B(_00283_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08944_ (.A(west_double[1]),
    .TE_B(_00284_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08945_ (.A(west_double[0]),
    .TE_B(_00285_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08946_ (.A(west_single[3]),
    .TE_B(_00286_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08947_ (.A(west_single[2]),
    .TE_B(_00287_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08948_ (.A(west_single[1]),
    .TE_B(_00288_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08949_ (.A(west_single[0]),
    .TE_B(_00289_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08950_ (.A(set_out_hard),
    .TE_B(_00290_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08951_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00291_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08952_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00292_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08953_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00293_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08954_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00294_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08955_ (.A(east_double[3]),
    .TE_B(_00295_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08956_ (.A(east_double[2]),
    .TE_B(_00296_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08957_ (.A(east_double[1]),
    .TE_B(_00297_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08958_ (.A(east_double[0]),
    .TE_B(_00298_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08959_ (.A(west_double[3]),
    .TE_B(_00299_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08960_ (.A(west_double[2]),
    .TE_B(_00300_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08961_ (.A(west_double[1]),
    .TE_B(_00301_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08962_ (.A(west_double[0]),
    .TE_B(_00302_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08963_ (.A(west_single[3]),
    .TE_B(_00303_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08964_ (.A(west_single[2]),
    .TE_B(_00304_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08965_ (.A(west_single[1]),
    .TE_B(_00305_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08966_ (.A(west_single[0]),
    .TE_B(_00306_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08967_ (.A(set_out_hard),
    .TE_B(_00307_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08968_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00308_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08969_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00309_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08970_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00310_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08971_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00311_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08972_ (.A(east_double[3]),
    .TE_B(_00312_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08973_ (.A(east_double[2]),
    .TE_B(_00313_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08974_ (.A(east_double[1]),
    .TE_B(_00314_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08975_ (.A(east_double[0]),
    .TE_B(_00315_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08976_ (.A(west_double[3]),
    .TE_B(_00316_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08977_ (.A(west_double[2]),
    .TE_B(_00317_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08978_ (.A(west_double[1]),
    .TE_B(_00318_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08979_ (.A(west_double[0]),
    .TE_B(_00319_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08980_ (.A(west_single[3]),
    .TE_B(_00320_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08981_ (.A(west_single[2]),
    .TE_B(_00321_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08982_ (.A(west_single[1]),
    .TE_B(_00322_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08983_ (.A(west_single[0]),
    .TE_B(_00323_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08984_ (.A(set_out_hard),
    .TE_B(_00324_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08985_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00325_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08986_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00326_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08987_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00327_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08988_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00328_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08989_ (.A(east_double[3]),
    .TE_B(_00329_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08990_ (.A(east_double[2]),
    .TE_B(_00330_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08991_ (.A(east_double[1]),
    .TE_B(_00331_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08992_ (.A(east_double[0]),
    .TE_B(_00332_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08993_ (.A(west_double[3]),
    .TE_B(_00333_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08994_ (.A(west_double[2]),
    .TE_B(_00334_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08995_ (.A(west_double[1]),
    .TE_B(_00335_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08996_ (.A(west_double[0]),
    .TE_B(_00336_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08997_ (.A(west_single[3]),
    .TE_B(_00337_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08998_ (.A(west_single[2]),
    .TE_B(_00338_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _08999_ (.A(west_single[1]),
    .TE_B(_00339_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09000_ (.A(west_single[0]),
    .TE_B(_00340_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09001_ (.A(set_out_hard),
    .TE_B(_00341_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09002_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00342_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09003_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00343_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09004_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00344_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09005_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00345_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09006_ (.A(east_double[3]),
    .TE_B(_00346_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09007_ (.A(east_double[2]),
    .TE_B(_00347_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09008_ (.A(east_double[1]),
    .TE_B(_00348_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09009_ (.A(east_double[0]),
    .TE_B(_00349_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09010_ (.A(west_double[3]),
    .TE_B(_00350_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09011_ (.A(west_double[2]),
    .TE_B(_00351_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09012_ (.A(west_double[1]),
    .TE_B(_00352_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09013_ (.A(west_double[0]),
    .TE_B(_00353_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09014_ (.A(west_single[3]),
    .TE_B(_00354_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09015_ (.A(west_single[2]),
    .TE_B(_00355_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09016_ (.A(west_single[1]),
    .TE_B(_00356_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09017_ (.A(west_single[0]),
    .TE_B(_00357_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09018_ (.A(set_out_hard),
    .TE_B(_00358_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09019_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00359_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09020_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00360_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09021_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00361_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09022_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00362_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09023_ (.A(east_double[3]),
    .TE_B(_00363_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09024_ (.A(east_double[2]),
    .TE_B(_00364_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09025_ (.A(east_double[1]),
    .TE_B(_00365_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09026_ (.A(east_double[0]),
    .TE_B(_00366_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09027_ (.A(west_double[3]),
    .TE_B(_00367_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09028_ (.A(west_double[2]),
    .TE_B(_00368_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09029_ (.A(west_double[1]),
    .TE_B(_00369_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09030_ (.A(west_double[0]),
    .TE_B(_00370_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09031_ (.A(west_single[3]),
    .TE_B(_00371_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09032_ (.A(west_single[2]),
    .TE_B(_00372_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09033_ (.A(west_single[1]),
    .TE_B(_00373_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09034_ (.A(west_single[0]),
    .TE_B(_00374_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09035_ (.A(set_out_hard),
    .TE_B(_00375_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09036_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00376_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09037_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00377_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09038_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00378_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09039_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00379_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09040_ (.A(east_double[3]),
    .TE_B(_00380_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09041_ (.A(east_double[2]),
    .TE_B(_00381_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09042_ (.A(east_double[1]),
    .TE_B(_00382_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09043_ (.A(east_double[0]),
    .TE_B(_00383_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09044_ (.A(west_double[3]),
    .TE_B(_00384_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09045_ (.A(west_double[2]),
    .TE_B(_00385_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09046_ (.A(west_double[1]),
    .TE_B(_00386_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09047_ (.A(west_double[0]),
    .TE_B(_00387_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09048_ (.A(west_single[3]),
    .TE_B(_00388_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09049_ (.A(west_single[2]),
    .TE_B(_00389_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09050_ (.A(west_single[1]),
    .TE_B(_00390_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09051_ (.A(west_single[0]),
    .TE_B(_00391_),
    .Z(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09052_ (.A(set_out_hard),
    .TE_B(_00191_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _09053_ (.A(set_out_hard),
    .TE_B(_00197_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _09054_ (.A(set_out_hard),
    .TE_B(_00203_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _09055_ (.A(set_out_hard),
    .TE_B(_00209_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _09056_ (.A(set_out_hard),
    .TE_B(_00215_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09057_ (.A(set_out_hard),
    .TE_B(_00221_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09058_ (.A(set_out_hard),
    .TE_B(_00227_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09059_ (.A(set_out_hard),
    .TE_B(_00233_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09060_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00192_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _09061_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00198_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _09062_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00204_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _09063_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00210_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _09064_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00216_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09065_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00222_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09066_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00228_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09067_ (.A(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00234_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09068_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00193_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _09069_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00199_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _09070_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00205_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _09071_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00211_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _09072_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00217_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09073_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00223_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09074_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00229_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09075_ (.A(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00235_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09076_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00194_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _09077_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00200_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _09078_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00206_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _09079_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00212_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _09080_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00218_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09081_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00224_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09082_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00230_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09083_ (.A(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00236_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09084_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00195_),
    .Z(west_double[3]));
 sky130_fd_sc_hd__ebufn_4 _09085_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00201_),
    .Z(west_double[2]));
 sky130_fd_sc_hd__ebufn_4 _09086_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00207_),
    .Z(west_double[1]));
 sky130_fd_sc_hd__ebufn_4 _09087_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00213_),
    .Z(west_double[0]));
 sky130_fd_sc_hd__ebufn_4 _09088_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00219_),
    .Z(west_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09089_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00225_),
    .Z(west_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09090_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00231_),
    .Z(west_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09091_ (.A(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00237_),
    .Z(west_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09092_ (.A(cb_north_in[4]),
    .TE_B(_00392_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09093_ (.A(cb_north_in[3]),
    .TE_B(_00393_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09094_ (.A(cb_north_in[2]),
    .TE_B(_00394_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09095_ (.A(cb_north_in[1]),
    .TE_B(_00395_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09096_ (.A(cb_north_in[0]),
    .TE_B(_00396_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09097_ (.A(east_double[3]),
    .TE_B(_00397_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09098_ (.A(east_double[2]),
    .TE_B(_00398_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09099_ (.A(east_double[1]),
    .TE_B(_00399_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09100_ (.A(east_double[0]),
    .TE_B(_00400_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09101_ (.A(west_double[3]),
    .TE_B(_00401_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09102_ (.A(west_double[2]),
    .TE_B(_00402_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09103_ (.A(west_double[1]),
    .TE_B(_00403_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09104_ (.A(west_double[0]),
    .TE_B(_00404_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09105_ (.A(west_single[3]),
    .TE_B(_00405_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09106_ (.A(west_single[2]),
    .TE_B(_00406_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09107_ (.A(west_single[1]),
    .TE_B(_00407_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09108_ (.A(west_single[0]),
    .TE_B(_00408_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09109_ (.A(cb_north_in[4]),
    .TE_B(_00409_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09110_ (.A(cb_north_in[3]),
    .TE_B(_00410_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09111_ (.A(cb_north_in[2]),
    .TE_B(_00411_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09112_ (.A(cb_north_in[1]),
    .TE_B(_00412_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09113_ (.A(cb_north_in[0]),
    .TE_B(_00413_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09114_ (.A(east_double[3]),
    .TE_B(_00414_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09115_ (.A(east_double[2]),
    .TE_B(_00415_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09116_ (.A(east_double[1]),
    .TE_B(_00416_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09117_ (.A(east_double[0]),
    .TE_B(_00417_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09118_ (.A(west_double[3]),
    .TE_B(_00418_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09119_ (.A(west_double[2]),
    .TE_B(_00419_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09120_ (.A(west_double[1]),
    .TE_B(_00420_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09121_ (.A(west_double[0]),
    .TE_B(_00421_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09122_ (.A(west_single[3]),
    .TE_B(_00422_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09123_ (.A(west_single[2]),
    .TE_B(_00423_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09124_ (.A(west_single[1]),
    .TE_B(_00424_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09125_ (.A(west_single[0]),
    .TE_B(_00425_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09126_ (.A(cb_north_in[4]),
    .TE_B(_00426_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09127_ (.A(cb_north_in[3]),
    .TE_B(_00427_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09128_ (.A(cb_north_in[2]),
    .TE_B(_00428_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09129_ (.A(cb_north_in[1]),
    .TE_B(_00429_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09130_ (.A(cb_north_in[0]),
    .TE_B(_00430_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09131_ (.A(east_double[3]),
    .TE_B(_00431_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09132_ (.A(east_double[2]),
    .TE_B(_00432_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09133_ (.A(east_double[1]),
    .TE_B(_00433_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09134_ (.A(east_double[0]),
    .TE_B(_00434_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09135_ (.A(west_double[3]),
    .TE_B(_00435_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09136_ (.A(west_double[2]),
    .TE_B(_00436_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09137_ (.A(west_double[1]),
    .TE_B(_00437_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09138_ (.A(west_double[0]),
    .TE_B(_00438_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09139_ (.A(west_single[3]),
    .TE_B(_00439_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09140_ (.A(west_single[2]),
    .TE_B(_00440_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09141_ (.A(west_single[1]),
    .TE_B(_00441_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09142_ (.A(west_single[0]),
    .TE_B(_00442_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09143_ (.A(cb_north_in[4]),
    .TE_B(_00443_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09144_ (.A(cb_north_in[3]),
    .TE_B(_00444_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09145_ (.A(cb_north_in[2]),
    .TE_B(_00445_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09146_ (.A(cb_north_in[1]),
    .TE_B(_00446_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09147_ (.A(cb_north_in[0]),
    .TE_B(_00447_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09148_ (.A(east_double[3]),
    .TE_B(_00448_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09149_ (.A(east_double[2]),
    .TE_B(_00449_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09150_ (.A(east_double[1]),
    .TE_B(_00450_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09151_ (.A(east_double[0]),
    .TE_B(_00451_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09152_ (.A(west_double[3]),
    .TE_B(_00452_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09153_ (.A(west_double[2]),
    .TE_B(_00453_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09154_ (.A(west_double[1]),
    .TE_B(_00454_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09155_ (.A(west_double[0]),
    .TE_B(_00455_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09156_ (.A(west_single[3]),
    .TE_B(_00456_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09157_ (.A(west_single[2]),
    .TE_B(_00457_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09158_ (.A(west_single[1]),
    .TE_B(_00458_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09159_ (.A(west_single[0]),
    .TE_B(_00459_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09160_ (.A(cb_north_in[4]),
    .TE_B(_00460_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09161_ (.A(cb_north_in[3]),
    .TE_B(_00461_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09162_ (.A(cb_north_in[2]),
    .TE_B(_00462_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09163_ (.A(cb_north_in[1]),
    .TE_B(_00463_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09164_ (.A(cb_north_in[0]),
    .TE_B(_00464_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09165_ (.A(east_double[3]),
    .TE_B(_00465_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09166_ (.A(east_double[2]),
    .TE_B(_00466_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09167_ (.A(east_double[1]),
    .TE_B(_00467_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09168_ (.A(east_double[0]),
    .TE_B(_00468_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09169_ (.A(west_double[3]),
    .TE_B(_00469_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09170_ (.A(west_double[2]),
    .TE_B(_00470_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09171_ (.A(west_double[1]),
    .TE_B(_00471_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09172_ (.A(west_double[0]),
    .TE_B(_00472_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09173_ (.A(west_single[3]),
    .TE_B(_00473_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09174_ (.A(west_single[2]),
    .TE_B(_00474_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09175_ (.A(west_single[1]),
    .TE_B(_00475_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09176_ (.A(west_single[0]),
    .TE_B(_00476_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09177_ (.A(cb_north_in[4]),
    .TE_B(_00477_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09178_ (.A(cb_north_in[3]),
    .TE_B(_00478_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09179_ (.A(cb_north_in[2]),
    .TE_B(_00479_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09180_ (.A(cb_north_in[1]),
    .TE_B(_00480_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09181_ (.A(cb_north_in[0]),
    .TE_B(_00481_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09182_ (.A(east_double[3]),
    .TE_B(_00482_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09183_ (.A(east_double[2]),
    .TE_B(_00483_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09184_ (.A(east_double[1]),
    .TE_B(_00484_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09185_ (.A(east_double[0]),
    .TE_B(_00485_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09186_ (.A(west_double[3]),
    .TE_B(_00486_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09187_ (.A(west_double[2]),
    .TE_B(_00487_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09188_ (.A(west_double[1]),
    .TE_B(_00488_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09189_ (.A(west_double[0]),
    .TE_B(_00489_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09190_ (.A(west_single[3]),
    .TE_B(_00490_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09191_ (.A(west_single[2]),
    .TE_B(_00491_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09192_ (.A(west_single[1]),
    .TE_B(_00492_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09193_ (.A(west_single[0]),
    .TE_B(_00493_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09194_ (.A(cb_north_in[4]),
    .TE_B(_00494_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09195_ (.A(cb_north_in[3]),
    .TE_B(_00495_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09196_ (.A(cb_north_in[2]),
    .TE_B(_00496_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09197_ (.A(cb_north_in[1]),
    .TE_B(_00497_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09198_ (.A(cb_north_in[0]),
    .TE_B(_00498_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09199_ (.A(east_double[3]),
    .TE_B(_00499_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09200_ (.A(east_double[2]),
    .TE_B(_00500_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09201_ (.A(east_double[1]),
    .TE_B(_00501_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09202_ (.A(east_double[0]),
    .TE_B(_00502_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09203_ (.A(west_double[3]),
    .TE_B(_00503_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09204_ (.A(west_double[2]),
    .TE_B(_00504_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09205_ (.A(west_double[1]),
    .TE_B(_00505_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09206_ (.A(west_double[0]),
    .TE_B(_00506_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09207_ (.A(west_single[3]),
    .TE_B(_00507_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09208_ (.A(west_single[2]),
    .TE_B(_00508_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09209_ (.A(west_single[1]),
    .TE_B(_00509_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09210_ (.A(west_single[0]),
    .TE_B(_00510_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09211_ (.A(cb_north_in[4]),
    .TE_B(_00511_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09212_ (.A(cb_north_in[3]),
    .TE_B(_00512_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09213_ (.A(cb_north_in[2]),
    .TE_B(_00513_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09214_ (.A(cb_north_in[1]),
    .TE_B(_00514_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09215_ (.A(cb_north_in[0]),
    .TE_B(_00515_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09216_ (.A(east_double[3]),
    .TE_B(_00516_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09217_ (.A(east_double[2]),
    .TE_B(_00517_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09218_ (.A(east_double[1]),
    .TE_B(_00518_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09219_ (.A(east_double[0]),
    .TE_B(_00519_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09220_ (.A(west_double[3]),
    .TE_B(_00520_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09221_ (.A(west_double[2]),
    .TE_B(_00521_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09222_ (.A(west_double[1]),
    .TE_B(_00522_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09223_ (.A(west_double[0]),
    .TE_B(_00523_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09224_ (.A(west_single[3]),
    .TE_B(_00524_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09225_ (.A(west_single[2]),
    .TE_B(_00525_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09226_ (.A(west_single[1]),
    .TE_B(_00526_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09227_ (.A(west_single[0]),
    .TE_B(_00527_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09228_ (.A(cb_north_in[4]),
    .TE_B(_00528_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09229_ (.A(cb_north_in[3]),
    .TE_B(_00529_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09230_ (.A(cb_north_in[2]),
    .TE_B(_00530_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09231_ (.A(cb_north_in[1]),
    .TE_B(_00531_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09232_ (.A(cb_north_in[0]),
    .TE_B(_00532_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09233_ (.A(east_double[3]),
    .TE_B(_00533_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09234_ (.A(east_double[2]),
    .TE_B(_00534_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09235_ (.A(east_double[1]),
    .TE_B(_00535_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09236_ (.A(east_double[0]),
    .TE_B(_00536_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09237_ (.A(west_double[3]),
    .TE_B(_00537_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09238_ (.A(west_double[2]),
    .TE_B(_00538_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09239_ (.A(west_double[1]),
    .TE_B(_00539_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09240_ (.A(west_double[0]),
    .TE_B(_00540_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09241_ (.A(west_single[3]),
    .TE_B(_00541_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09242_ (.A(west_single[2]),
    .TE_B(_00542_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09243_ (.A(west_single[1]),
    .TE_B(_00543_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09244_ (.A(west_single[0]),
    .TE_B(_00544_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09245_ (.A(cb_north_in[4]),
    .TE_B(_00545_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09246_ (.A(cb_north_in[3]),
    .TE_B(_00546_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09247_ (.A(cb_north_in[2]),
    .TE_B(_00547_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09248_ (.A(cb_north_in[1]),
    .TE_B(_00548_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09249_ (.A(cb_north_in[0]),
    .TE_B(_00549_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09250_ (.A(east_double[3]),
    .TE_B(_00550_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09251_ (.A(east_double[2]),
    .TE_B(_00551_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09252_ (.A(east_double[1]),
    .TE_B(_00552_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09253_ (.A(east_double[0]),
    .TE_B(_00553_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09254_ (.A(west_double[3]),
    .TE_B(_00554_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09255_ (.A(west_double[2]),
    .TE_B(_00555_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09256_ (.A(west_double[1]),
    .TE_B(_00556_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09257_ (.A(west_double[0]),
    .TE_B(_00557_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09258_ (.A(west_single[3]),
    .TE_B(_00558_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09259_ (.A(west_single[2]),
    .TE_B(_00559_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09260_ (.A(west_single[1]),
    .TE_B(_00560_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09261_ (.A(west_single[0]),
    .TE_B(_00561_),
    .Z(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09262_ (.A(cb_east_in[4]),
    .TE_B(_00562_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _09263_ (.A(cb_east_in[4]),
    .TE_B(_00563_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _09264_ (.A(cb_east_in[4]),
    .TE_B(_00564_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _09265_ (.A(cb_east_in[4]),
    .TE_B(_00565_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _09266_ (.A(cb_east_in[4]),
    .TE_B(_00566_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09267_ (.A(cb_east_in[4]),
    .TE_B(_00567_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09268_ (.A(cb_east_in[4]),
    .TE_B(_00568_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09269_ (.A(cb_east_in[4]),
    .TE_B(_00569_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09270_ (.A(cb_east_in[3]),
    .TE_B(_00570_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _09271_ (.A(cb_east_in[3]),
    .TE_B(_00571_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _09272_ (.A(cb_east_in[3]),
    .TE_B(_00572_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _09273_ (.A(cb_east_in[3]),
    .TE_B(_00573_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _09274_ (.A(cb_east_in[3]),
    .TE_B(_00574_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09275_ (.A(cb_east_in[3]),
    .TE_B(_00575_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09276_ (.A(cb_east_in[3]),
    .TE_B(_00576_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09277_ (.A(cb_east_in[3]),
    .TE_B(_00577_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09278_ (.A(cb_east_in[2]),
    .TE_B(_00578_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _09279_ (.A(cb_east_in[2]),
    .TE_B(_00579_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _09280_ (.A(cb_east_in[2]),
    .TE_B(_00580_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _09281_ (.A(cb_east_in[2]),
    .TE_B(_00581_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _09282_ (.A(cb_east_in[2]),
    .TE_B(_00582_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09283_ (.A(cb_east_in[2]),
    .TE_B(_00583_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09284_ (.A(cb_east_in[2]),
    .TE_B(_00584_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09285_ (.A(cb_east_in[2]),
    .TE_B(_00585_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09286_ (.A(cb_east_in[1]),
    .TE_B(_00586_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _09287_ (.A(cb_east_in[1]),
    .TE_B(_00587_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _09288_ (.A(cb_east_in[1]),
    .TE_B(_00588_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _09289_ (.A(cb_east_in[1]),
    .TE_B(_00589_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _09290_ (.A(cb_east_in[1]),
    .TE_B(_00590_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09291_ (.A(cb_east_in[1]),
    .TE_B(_00591_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09292_ (.A(cb_east_in[1]),
    .TE_B(_00592_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09293_ (.A(cb_east_in[1]),
    .TE_B(_00593_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09294_ (.A(cb_east_in[0]),
    .TE_B(_00594_),
    .Z(north_double[7]));
 sky130_fd_sc_hd__ebufn_4 _09295_ (.A(cb_east_in[0]),
    .TE_B(_00595_),
    .Z(north_double[6]));
 sky130_fd_sc_hd__ebufn_4 _09296_ (.A(cb_east_in[0]),
    .TE_B(_00596_),
    .Z(north_double[5]));
 sky130_fd_sc_hd__ebufn_4 _09297_ (.A(cb_east_in[0]),
    .TE_B(_00597_),
    .Z(north_double[4]));
 sky130_fd_sc_hd__ebufn_4 _09298_ (.A(cb_east_in[0]),
    .TE_B(_00598_),
    .Z(south_single[3]));
 sky130_fd_sc_hd__ebufn_4 _09299_ (.A(cb_east_in[0]),
    .TE_B(_00599_),
    .Z(south_single[2]));
 sky130_fd_sc_hd__ebufn_4 _09300_ (.A(cb_east_in[0]),
    .TE_B(_00600_),
    .Z(south_single[1]));
 sky130_fd_sc_hd__ebufn_4 _09301_ (.A(cb_east_in[0]),
    .TE_B(_00601_),
    .Z(south_single[0]));
 sky130_fd_sc_hd__ebufn_4 _09302_ (.A(shift_out_hard),
    .TE_B(_00602_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09303_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00603_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09304_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00604_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09305_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00605_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09306_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00606_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09307_ (.A(south_double[7]),
    .TE_B(_00607_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09308_ (.A(south_double[6]),
    .TE_B(_00608_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09309_ (.A(south_double[5]),
    .TE_B(_00609_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09310_ (.A(south_double[4]),
    .TE_B(_00610_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09311_ (.A(north_double[7]),
    .TE_B(_00616_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09312_ (.A(north_double[6]),
    .TE_B(_00622_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09313_ (.A(north_double[5]),
    .TE_B(_00628_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09314_ (.A(north_double[4]),
    .TE_B(_00634_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09315_ (.A(south_single[3]),
    .TE_B(_00640_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09316_ (.A(south_single[2]),
    .TE_B(_00646_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09317_ (.A(south_single[1]),
    .TE_B(_00652_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09318_ (.A(south_single[0]),
    .TE_B(_00658_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09319_ (.A(shift_out_hard),
    .TE_B(_00659_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09320_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00660_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09321_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00661_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09322_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00662_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09323_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00663_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09324_ (.A(south_double[7]),
    .TE_B(_00664_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09325_ (.A(south_double[6]),
    .TE_B(_00665_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09326_ (.A(south_double[5]),
    .TE_B(_00666_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09327_ (.A(south_double[4]),
    .TE_B(_00667_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09328_ (.A(north_double[7]),
    .TE_B(_00668_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09329_ (.A(north_double[6]),
    .TE_B(_00669_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09330_ (.A(north_double[5]),
    .TE_B(_00670_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09331_ (.A(north_double[4]),
    .TE_B(_00671_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09332_ (.A(south_single[3]),
    .TE_B(_00672_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09333_ (.A(south_single[2]),
    .TE_B(_00673_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09334_ (.A(south_single[1]),
    .TE_B(_00674_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09335_ (.A(south_single[0]),
    .TE_B(_00675_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09336_ (.A(shift_out_hard),
    .TE_B(_00676_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09337_ (.A(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .TE_B(_00677_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09338_ (.A(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .TE_B(_00678_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09339_ (.A(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ),
    .TE_B(_00679_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09340_ (.A(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.b ),
    .TE_B(_00680_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09341_ (.A(south_double[7]),
    .TE_B(_00681_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09342_ (.A(south_double[6]),
    .TE_B(_00682_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09343_ (.A(south_double[5]),
    .TE_B(_00683_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09344_ (.A(south_double[4]),
    .TE_B(_00684_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09345_ (.A(north_double[7]),
    .TE_B(_00685_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__ebufn_4 _09346_ (.A(north_double[6]),
    .TE_B(_00686_),
    .Z(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.a ));
 sky130_fd_sc_hd__dfxtp_4 _09347_ (.D(_02023_),
    .Q(_04315_),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09348_ (.D(_02024_),
    .Q(\slice.sliceluroni.muxes.config_state[0] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09349_ (.D(_02025_),
    .Q(\slice.sliceluroni.muxes.config_state[1] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09350_ (.D(_02026_),
    .Q(\slice.sliceluroni.use_cc ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09351_ (.D(_02027_),
    .Q(_04168_),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09352_ (.D(_02028_),
    .Q(_04217_),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09353_ (.D(_02029_),
    .Q(_04266_),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09354_ (.D(_02030_),
    .Q(clb_west_out[2]),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09355_ (.D(_02031_),
    .Q(clb_west_out[3]),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09356_ (.D(_02032_),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09357_ (.D(_02033_),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09358_ (.D(_02034_),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.b ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09359_ (.D(_02035_),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.b ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09360_ (.D(_02036_),
    .Q(clb_south_out[2]),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09361_ (.D(_02037_),
    .Q(clb_south_out[3]),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09362_ (.D(_02039_),
    .Q(\cb_east.inst.configuroni.comb_shifter.config_data[421] ),
    .CLK(clknet_7_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09363_ (.D(_02041_),
    .Q(shift_out_hard),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09364_ (.D(_02043_),
    .Q(\cb_east.inst.cb_conf_bus[1] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09365_ (.D(_02045_),
    .Q(\cb_east.inst.cb_conf_bus[2] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09366_ (.D(_02047_),
    .Q(\cb_east.inst.cb_conf_bus[3] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09367_ (.D(_02049_),
    .Q(\cb_east.inst.cb_conf_bus[4] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09368_ (.D(_02051_),
    .Q(\cb_east.inst.cb_conf_bus[5] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09369_ (.D(_02053_),
    .Q(\cb_east.inst.cb_conf_bus[6] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09370_ (.D(_02055_),
    .Q(\cb_east.inst.cb_conf_bus[7] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09371_ (.D(_02057_),
    .Q(\cb_east.inst.cb_conf_bus[8] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09372_ (.D(_02059_),
    .Q(\cb_east.inst.cb_conf_bus[9] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09373_ (.D(_02061_),
    .Q(\cb_east.inst.cb_conf_bus[10] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09374_ (.D(_02063_),
    .Q(\cb_east.inst.cb_conf_bus[11] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09375_ (.D(_02065_),
    .Q(\cb_east.inst.cb_conf_bus[12] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09376_ (.D(_02067_),
    .Q(\cb_east.inst.cb_conf_bus[13] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09377_ (.D(_02069_),
    .Q(\cb_east.inst.cb_conf_bus[14] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09378_ (.D(_02071_),
    .Q(\cb_east.inst.cb_conf_bus[15] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09379_ (.D(_02073_),
    .Q(\cb_east.inst.cb_conf_bus[16] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09380_ (.D(_02075_),
    .Q(\cb_east.inst.cb_conf_bus[17] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09381_ (.D(_02077_),
    .Q(\cb_east.inst.cb_conf_bus[18] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09382_ (.D(_02079_),
    .Q(\cb_east.inst.cb_conf_bus[19] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09383_ (.D(_02081_),
    .Q(\cb_east.inst.cb_conf_bus[20] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09384_ (.D(_02083_),
    .Q(\cb_east.inst.cb_conf_bus[21] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09385_ (.D(_02085_),
    .Q(\cb_east.inst.cb_conf_bus[22] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09386_ (.D(_02087_),
    .Q(\cb_east.inst.cb_conf_bus[23] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09387_ (.D(_02089_),
    .Q(\cb_east.inst.cb_conf_bus[24] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09388_ (.D(_02091_),
    .Q(\cb_east.inst.cb_conf_bus[25] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09389_ (.D(_02093_),
    .Q(\cb_east.inst.cb_conf_bus[26] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09390_ (.D(_02095_),
    .Q(\cb_east.inst.cb_conf_bus[27] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09391_ (.D(_02097_),
    .Q(\cb_east.inst.cb_conf_bus[28] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09392_ (.D(_02099_),
    .Q(\cb_east.inst.cb_conf_bus[29] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09393_ (.D(_02101_),
    .Q(\cb_east.inst.cb_conf_bus[30] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09394_ (.D(_02103_),
    .Q(\cb_east.inst.cb_conf_bus[31] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09395_ (.D(_02105_),
    .Q(\cb_east.inst.cb_conf_bus[32] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09396_ (.D(_02107_),
    .Q(\cb_east.inst.cb_conf_bus[33] ),
    .CLK(clknet_7_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09397_ (.D(_02109_),
    .Q(\cb_east.inst.cb_conf_bus[34] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09398_ (.D(_02111_),
    .Q(\cb_east.inst.cb_conf_bus[35] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09399_ (.D(_02113_),
    .Q(\cb_east.inst.cb_conf_bus[36] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09400_ (.D(_02115_),
    .Q(\cb_east.inst.cb_conf_bus[37] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09401_ (.D(_02117_),
    .Q(\cb_east.inst.cb_conf_bus[38] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09402_ (.D(_02119_),
    .Q(\cb_east.inst.cb_conf_bus[39] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09403_ (.D(_02121_),
    .Q(\cb_east.inst.cb_conf_bus[40] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09404_ (.D(_02123_),
    .Q(\cb_east.inst.cb_conf_bus[41] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09405_ (.D(_02125_),
    .Q(\cb_east.inst.cb_conf_bus[42] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09406_ (.D(_02127_),
    .Q(\cb_east.inst.cb_conf_bus[43] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09407_ (.D(_02129_),
    .Q(\cb_east.inst.cb_conf_bus[44] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09408_ (.D(_02131_),
    .Q(\cb_east.inst.cb_conf_bus[45] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09409_ (.D(_02133_),
    .Q(\cb_east.inst.cb_conf_bus[46] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09410_ (.D(_02135_),
    .Q(\cb_east.inst.cb_conf_bus[47] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09411_ (.D(_02137_),
    .Q(\cb_east.inst.cb_conf_bus[48] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09412_ (.D(_02139_),
    .Q(\cb_east.inst.cb_conf_bus[49] ),
    .CLK(clknet_7_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09413_ (.D(_02141_),
    .Q(\cb_east.inst.cb_conf_bus[50] ),
    .CLK(clknet_7_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09414_ (.D(_02143_),
    .Q(\cb_east.inst.cb_conf_bus[51] ),
    .CLK(clknet_7_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09415_ (.D(_02145_),
    .Q(\cb_east.inst.cb_conf_bus[52] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09416_ (.D(_02147_),
    .Q(\cb_east.inst.cb_conf_bus[53] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09417_ (.D(_02149_),
    .Q(\cb_east.inst.cb_conf_bus[54] ),
    .CLK(clknet_7_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09418_ (.D(_02151_),
    .Q(\cb_east.inst.cb_conf_bus[55] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09419_ (.D(_02153_),
    .Q(\cb_east.inst.cb_conf_bus[56] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09420_ (.D(_02155_),
    .Q(\cb_east.inst.cb_conf_bus[57] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09421_ (.D(_02157_),
    .Q(\cb_east.inst.cb_conf_bus[58] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09422_ (.D(_02159_),
    .Q(\cb_east.inst.cb_conf_bus[59] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09423_ (.D(_02161_),
    .Q(\cb_east.inst.cb_conf_bus[60] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09424_ (.D(_02163_),
    .Q(\cb_east.inst.cb_conf_bus[61] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09425_ (.D(_02165_),
    .Q(\cb_east.inst.cb_conf_bus[62] ),
    .CLK(clknet_7_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09426_ (.D(_02167_),
    .Q(\cb_east.inst.cb_conf_bus[63] ),
    .CLK(clknet_7_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09427_ (.D(_02169_),
    .Q(\cb_east.inst.cb_conf_bus[64] ),
    .CLK(clknet_7_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09428_ (.D(_02171_),
    .Q(\cb_east.inst.cb_conf_bus[65] ),
    .CLK(clknet_7_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09429_ (.D(_02173_),
    .Q(\cb_east.inst.cb_conf_bus[66] ),
    .CLK(clknet_7_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09430_ (.D(_02175_),
    .Q(\cb_east.inst.cb_conf_bus[67] ),
    .CLK(clknet_7_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09431_ (.D(_02177_),
    .Q(\cb_east.inst.cb_conf_bus[68] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09432_ (.D(_02179_),
    .Q(\cb_east.inst.cb_conf_bus[69] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09433_ (.D(_02181_),
    .Q(\cb_east.inst.cb_conf_bus[70] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09434_ (.D(_02183_),
    .Q(\cb_east.inst.cb_conf_bus[71] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09435_ (.D(_02185_),
    .Q(\cb_east.inst.cb_conf_bus[72] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09436_ (.D(_02187_),
    .Q(\cb_east.inst.cb_conf_bus[73] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09437_ (.D(_02189_),
    .Q(\cb_east.inst.cb_conf_bus[74] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09438_ (.D(_02191_),
    .Q(\cb_east.inst.cb_conf_bus[75] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09439_ (.D(_02193_),
    .Q(\cb_east.inst.cb_conf_bus[76] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09440_ (.D(_02195_),
    .Q(\cb_east.inst.cb_conf_bus[77] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09441_ (.D(_02197_),
    .Q(\cb_east.inst.cb_conf_bus[78] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09442_ (.D(_02199_),
    .Q(\cb_east.inst.cb_conf_bus[79] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09443_ (.D(_02201_),
    .Q(\cb_east.inst.cb_conf_bus[80] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09444_ (.D(_02203_),
    .Q(\cb_east.inst.cb_conf_bus[81] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09445_ (.D(_02205_),
    .Q(\cb_east.inst.cb_conf_bus[82] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09446_ (.D(_02207_),
    .Q(\cb_east.inst.cb_conf_bus[83] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09447_ (.D(_02209_),
    .Q(\cb_east.inst.cb_conf_bus[84] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09448_ (.D(_02211_),
    .Q(\cb_east.inst.cb_conf_bus[85] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09449_ (.D(_02213_),
    .Q(\cb_east.inst.cb_conf_bus[86] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09450_ (.D(_02215_),
    .Q(\cb_east.inst.cb_conf_bus[87] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09451_ (.D(_02217_),
    .Q(\cb_east.inst.cb_conf_bus[88] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09452_ (.D(_02219_),
    .Q(\cb_east.inst.cb_conf_bus[89] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09453_ (.D(_02221_),
    .Q(\cb_east.inst.cb_conf_bus[90] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09454_ (.D(_02223_),
    .Q(\cb_east.inst.cb_conf_bus[91] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09455_ (.D(_02225_),
    .Q(\cb_east.inst.cb_conf_bus[92] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09456_ (.D(_02227_),
    .Q(\cb_east.inst.cb_conf_bus[93] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09457_ (.D(_02229_),
    .Q(\cb_east.inst.cb_conf_bus[94] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09458_ (.D(_02231_),
    .Q(\cb_east.inst.cb_conf_bus[95] ),
    .CLK(clknet_7_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09459_ (.D(_02233_),
    .Q(\cb_east.inst.cb_conf_bus[96] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09460_ (.D(_02235_),
    .Q(\cb_east.inst.cb_conf_bus[97] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09461_ (.D(_02237_),
    .Q(\cb_east.inst.cb_conf_bus[98] ),
    .CLK(clknet_7_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09462_ (.D(_02239_),
    .Q(\cb_east.inst.cb_conf_bus[99] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09463_ (.D(_02241_),
    .Q(\cb_east.inst.cb_conf_bus[100] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09464_ (.D(_02243_),
    .Q(\cb_east.inst.cb_conf_bus[101] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09465_ (.D(_02245_),
    .Q(\cb_east.inst.cb_conf_bus[102] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09466_ (.D(_02247_),
    .Q(\cb_east.inst.cb_conf_bus[103] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09467_ (.D(_02249_),
    .Q(\cb_east.inst.cb_conf_bus[104] ),
    .CLK(clknet_7_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09468_ (.D(_02251_),
    .Q(\cb_east.inst.cb_conf_bus[105] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09469_ (.D(_02253_),
    .Q(\cb_east.inst.cb_conf_bus[106] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09470_ (.D(_02255_),
    .Q(\cb_east.inst.cb_conf_bus[107] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09471_ (.D(_02257_),
    .Q(\cb_east.inst.cb_conf_bus[108] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09472_ (.D(_02259_),
    .Q(\cb_east.inst.cb_conf_bus[109] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09473_ (.D(_02261_),
    .Q(\cb_east.inst.cb_conf_bus[110] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09474_ (.D(_02263_),
    .Q(\cb_east.inst.cb_conf_bus[111] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09475_ (.D(_02265_),
    .Q(\cb_east.inst.cb_conf_bus[112] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09476_ (.D(_02267_),
    .Q(\cb_east.inst.cb_conf_bus[113] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09477_ (.D(_02269_),
    .Q(\cb_east.inst.cb_conf_bus[114] ),
    .CLK(clknet_7_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09478_ (.D(_02271_),
    .Q(\cb_east.inst.cb_conf_bus[115] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09479_ (.D(_02273_),
    .Q(\cb_east.inst.cb_conf_bus[116] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09480_ (.D(_02275_),
    .Q(\cb_east.inst.cb_conf_bus[117] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09481_ (.D(_02277_),
    .Q(\cb_east.inst.cb_conf_bus[118] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09482_ (.D(_02279_),
    .Q(\cb_east.inst.cb_conf_bus[119] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09483_ (.D(_02281_),
    .Q(\cb_east.inst.cb_conf_bus[120] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09484_ (.D(_02283_),
    .Q(\cb_east.inst.cb_conf_bus[121] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09485_ (.D(_02285_),
    .Q(\cb_east.inst.cb_conf_bus[122] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09486_ (.D(_02287_),
    .Q(\cb_east.inst.cb_conf_bus[123] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09487_ (.D(_02289_),
    .Q(\cb_east.inst.cb_conf_bus[124] ),
    .CLK(clknet_7_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09488_ (.D(_02291_),
    .Q(\cb_east.inst.cb_conf_bus[125] ),
    .CLK(clknet_7_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09489_ (.D(_02293_),
    .Q(\cb_east.inst.cb_conf_bus[126] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09490_ (.D(_02295_),
    .Q(\cb_east.inst.cb_conf_bus[127] ),
    .CLK(clknet_7_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09491_ (.D(_02297_),
    .Q(\cb_east.inst.cb_conf_bus[128] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09492_ (.D(_02299_),
    .Q(\cb_east.inst.cb_conf_bus[129] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09493_ (.D(_02301_),
    .Q(\cb_east.inst.cb_conf_bus[130] ),
    .CLK(clknet_7_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09494_ (.D(_02303_),
    .Q(\cb_east.inst.cb_conf_bus[131] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09495_ (.D(_02305_),
    .Q(\cb_east.inst.cb_conf_bus[132] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09496_ (.D(_02307_),
    .Q(\cb_east.inst.cb_conf_bus[133] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09497_ (.D(_02309_),
    .Q(\cb_east.inst.cb_conf_bus[134] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09498_ (.D(_02311_),
    .Q(\cb_east.inst.cb_conf_bus[135] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09499_ (.D(_02313_),
    .Q(\cb_east.inst.cb_conf_bus[136] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09500_ (.D(_02315_),
    .Q(\cb_east.inst.cb_conf_bus[137] ),
    .CLK(clknet_7_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09501_ (.D(_02317_),
    .Q(\cb_east.inst.cb_conf_bus[138] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09502_ (.D(_02319_),
    .Q(\cb_east.inst.cb_conf_bus[139] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09503_ (.D(_02321_),
    .Q(\cb_east.inst.cb_conf_bus[140] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09504_ (.D(_02323_),
    .Q(\cb_east.inst.cb_conf_bus[141] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09505_ (.D(_02325_),
    .Q(\cb_east.inst.cb_conf_bus[142] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09506_ (.D(_02327_),
    .Q(\cb_east.inst.cb_conf_bus[143] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09507_ (.D(_02329_),
    .Q(\cb_east.inst.cb_conf_bus[144] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09508_ (.D(_02331_),
    .Q(\cb_east.inst.cb_conf_bus[145] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09509_ (.D(_02333_),
    .Q(\cb_east.inst.cb_conf_bus[146] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09510_ (.D(_02335_),
    .Q(\cb_east.inst.cb_conf_bus[147] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09511_ (.D(_02337_),
    .Q(\cb_east.inst.cb_conf_bus[148] ),
    .CLK(clknet_7_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09512_ (.D(_02339_),
    .Q(\cb_east.inst.cb_conf_bus[149] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09513_ (.D(_02341_),
    .Q(\cb_east.inst.cb_conf_bus[150] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09514_ (.D(_02343_),
    .Q(\cb_east.inst.cb_conf_bus[151] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09515_ (.D(_02345_),
    .Q(\cb_east.inst.cb_conf_bus[152] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09516_ (.D(_02347_),
    .Q(\cb_east.inst.cb_conf_bus[153] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09517_ (.D(_02349_),
    .Q(\cb_east.inst.cb_conf_bus[154] ),
    .CLK(clknet_7_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09518_ (.D(_02351_),
    .Q(\cb_east.inst.cb_conf_bus[155] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09519_ (.D(_02353_),
    .Q(\cb_east.inst.cb_conf_bus[156] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09520_ (.D(_02355_),
    .Q(\cb_east.inst.cb_conf_bus[157] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09521_ (.D(_02357_),
    .Q(\cb_east.inst.cb_conf_bus[158] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09522_ (.D(_02359_),
    .Q(\cb_east.inst.cb_conf_bus[159] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09523_ (.D(_02361_),
    .Q(\cb_east.inst.cb_conf_bus[160] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09524_ (.D(_02363_),
    .Q(\cb_east.inst.cb_conf_bus[161] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09525_ (.D(_02365_),
    .Q(\cb_east.inst.cb_conf_bus[162] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09526_ (.D(_02367_),
    .Q(\cb_east.inst.cb_conf_bus[163] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09527_ (.D(_02369_),
    .Q(\cb_east.inst.cb_conf_bus[164] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09528_ (.D(_02371_),
    .Q(\cb_east.inst.cb_conf_bus[165] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09529_ (.D(_02373_),
    .Q(\cb_east.inst.cb_conf_bus[166] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09530_ (.D(_02375_),
    .Q(\cb_east.inst.cb_conf_bus[167] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09531_ (.D(_02377_),
    .Q(\cb_east.inst.cb_conf_bus[168] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09532_ (.D(_02379_),
    .Q(\cb_east.inst.cb_conf_bus[169] ),
    .CLK(clknet_7_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09533_ (.D(_02381_),
    .Q(\cb_east.inst.cb_conf_bus[170] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09534_ (.D(_02383_),
    .Q(\cb_east.inst.cb_conf_bus[171] ),
    .CLK(clknet_7_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09535_ (.D(_02385_),
    .Q(\cb_east.inst.cb_conf_bus[172] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09536_ (.D(_02387_),
    .Q(\cb_east.inst.cb_conf_bus[173] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09537_ (.D(_02389_),
    .Q(\cb_east.inst.cb_conf_bus[174] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09538_ (.D(_02391_),
    .Q(\cb_east.inst.cb_conf_bus[175] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09539_ (.D(_02393_),
    .Q(\cb_east.inst.cb_conf_bus[176] ),
    .CLK(clknet_7_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09540_ (.D(_02395_),
    .Q(\cb_east.inst.cb_conf_bus[177] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09541_ (.D(_02397_),
    .Q(\cb_east.inst.cb_conf_bus[178] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09542_ (.D(_02399_),
    .Q(\cb_east.inst.cb_conf_bus[179] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09543_ (.D(_02401_),
    .Q(\cb_east.inst.cb_conf_bus[180] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09544_ (.D(_02403_),
    .Q(\cb_east.inst.cb_conf_bus[181] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09545_ (.D(_02405_),
    .Q(\cb_east.inst.cb_conf_bus[182] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09546_ (.D(_02407_),
    .Q(\cb_east.inst.cb_conf_bus[183] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09547_ (.D(_02409_),
    .Q(\cb_east.inst.cb_conf_bus[184] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09548_ (.D(_02411_),
    .Q(\cb_east.inst.cb_conf_bus[185] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09549_ (.D(_02413_),
    .Q(\cb_east.inst.cb_conf_bus[186] ),
    .CLK(clknet_7_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09550_ (.D(_02415_),
    .Q(\cb_east.inst.cb_conf_bus[187] ),
    .CLK(clknet_7_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09551_ (.D(_02417_),
    .Q(\cb_east.inst.cb_conf_bus[188] ),
    .CLK(clknet_7_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09552_ (.D(_02419_),
    .Q(\cb_east.inst.cb_conf_bus[189] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09553_ (.D(_02421_),
    .Q(\cb_east.inst.cb_conf_bus[190] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09554_ (.D(_02423_),
    .Q(\cb_east.inst.cb_conf_bus[191] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09555_ (.D(_02425_),
    .Q(\cb_east.inst.cb_conf_bus[192] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09556_ (.D(_02427_),
    .Q(\cb_east.inst.cb_conf_bus[193] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09557_ (.D(_02429_),
    .Q(\cb_east.inst.cb_conf_bus[194] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09558_ (.D(_02431_),
    .Q(\cb_east.inst.cb_conf_bus[195] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09559_ (.D(_02433_),
    .Q(\cb_east.inst.cb_conf_bus[196] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09560_ (.D(_02435_),
    .Q(\cb_east.inst.cb_conf_bus[197] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09561_ (.D(_02437_),
    .Q(\cb_east.inst.cb_conf_bus[198] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09562_ (.D(_02439_),
    .Q(\cb_east.inst.cb_conf_bus[199] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09563_ (.D(_02441_),
    .Q(\cb_east.inst.cb_conf_bus[200] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09564_ (.D(_02443_),
    .Q(\cb_east.inst.cb_conf_bus[201] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09565_ (.D(_02445_),
    .Q(\cb_east.inst.cb_conf_bus[202] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09566_ (.D(_02447_),
    .Q(\cb_east.inst.cb_conf_bus[203] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09567_ (.D(_02449_),
    .Q(\cb_east.inst.cb_conf_bus[204] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09568_ (.D(_02451_),
    .Q(\cb_east.inst.cb_conf_bus[205] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09569_ (.D(_02453_),
    .Q(\cb_east.inst.cb_conf_bus[206] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09570_ (.D(_02455_),
    .Q(\cb_east.inst.cb_conf_bus[207] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09571_ (.D(_02457_),
    .Q(\cb_east.inst.cb_conf_bus[208] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09572_ (.D(_02459_),
    .Q(\cb_east.inst.cb_conf_bus[209] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09573_ (.D(_02461_),
    .Q(\cb_east.inst.cb_conf_bus[210] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09574_ (.D(_02463_),
    .Q(\cb_east.inst.cb_conf_bus[211] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09575_ (.D(_02465_),
    .Q(\cb_east.inst.cb_conf_bus[212] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09576_ (.D(_02467_),
    .Q(\cb_east.inst.cb_conf_bus[213] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09577_ (.D(_02469_),
    .Q(\cb_east.inst.cb_conf_bus[214] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09578_ (.D(_02471_),
    .Q(\cb_east.inst.cb_conf_bus[215] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09579_ (.D(_02473_),
    .Q(\cb_east.inst.cb_conf_bus[216] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09580_ (.D(_02475_),
    .Q(\cb_east.inst.cb_conf_bus[217] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09581_ (.D(_02477_),
    .Q(\cb_east.inst.cb_conf_bus[218] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09582_ (.D(_02479_),
    .Q(\cb_east.inst.cb_conf_bus[219] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09583_ (.D(_02481_),
    .Q(\cb_east.inst.cb_conf_bus[220] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09584_ (.D(_02483_),
    .Q(\cb_east.inst.cb_conf_bus[221] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09585_ (.D(_02485_),
    .Q(\cb_east.inst.cb_conf_bus[222] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09586_ (.D(_02487_),
    .Q(\cb_east.inst.cb_conf_bus[223] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09587_ (.D(_02489_),
    .Q(\cb_east.inst.cb_conf_bus[224] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09588_ (.D(_02491_),
    .Q(\cb_east.inst.cb_conf_bus[225] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09589_ (.D(_02493_),
    .Q(\cb_east.inst.cb_conf_bus[226] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09590_ (.D(_02495_),
    .Q(\cb_east.inst.cb_conf_bus[227] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09591_ (.D(_02497_),
    .Q(\cb_east.inst.cb_conf_bus[228] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09592_ (.D(_02499_),
    .Q(\cb_east.inst.cb_conf_bus[229] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09593_ (.D(_02501_),
    .Q(\cb_east.inst.cb_conf_bus[230] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09594_ (.D(_02503_),
    .Q(\cb_east.inst.cb_conf_bus[231] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09595_ (.D(_02505_),
    .Q(\cb_east.inst.cb_conf_bus[232] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09596_ (.D(_02507_),
    .Q(\cb_east.inst.cb_conf_bus[233] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09597_ (.D(_02509_),
    .Q(\cb_east.inst.cb_conf_bus[234] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09598_ (.D(_02511_),
    .Q(\cb_east.inst.cb_conf_bus[235] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09599_ (.D(_02513_),
    .Q(\cb_east.inst.cb_conf_bus[236] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09600_ (.D(_02515_),
    .Q(\cb_east.inst.cb_conf_bus[237] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09601_ (.D(_02517_),
    .Q(\cb_east.inst.cb_conf_bus[238] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09602_ (.D(_02519_),
    .Q(\cb_east.inst.cb_conf_bus[239] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09603_ (.D(_02521_),
    .Q(\cb_east.inst.cb_conf_bus[240] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09604_ (.D(_02523_),
    .Q(\cb_east.inst.cb_conf_bus[241] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09605_ (.D(_02525_),
    .Q(\cb_east.inst.cb_conf_bus[242] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09606_ (.D(_02527_),
    .Q(\cb_east.inst.cb_conf_bus[243] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09607_ (.D(_02529_),
    .Q(\cb_east.inst.cb_conf_bus[244] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09608_ (.D(_02531_),
    .Q(\cb_east.inst.cb_conf_bus[245] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09609_ (.D(_02533_),
    .Q(\cb_east.inst.cb_conf_bus[246] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09610_ (.D(_02535_),
    .Q(\cb_east.inst.cb_conf_bus[247] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09611_ (.D(_02537_),
    .Q(\cb_east.inst.cb_conf_bus[248] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09612_ (.D(_02539_),
    .Q(\cb_east.inst.cb_conf_bus[249] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09613_ (.D(_02541_),
    .Q(\cb_east.inst.cb_conf_bus[250] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09614_ (.D(_02543_),
    .Q(\cb_east.inst.cb_conf_bus[251] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09615_ (.D(_02545_),
    .Q(\cb_east.inst.cb_conf_bus[252] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09616_ (.D(_02547_),
    .Q(\cb_east.inst.cb_conf_bus[253] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09617_ (.D(_02549_),
    .Q(\cb_east.inst.cb_conf_bus[254] ),
    .CLK(clknet_7_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09618_ (.D(_02551_),
    .Q(\cb_east.inst.cb_conf_bus[255] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09619_ (.D(_02553_),
    .Q(\cb_east.inst.cb_conf_bus[256] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09620_ (.D(_02555_),
    .Q(\cb_east.inst.cb_conf_bus[257] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09621_ (.D(_02557_),
    .Q(\cb_east.inst.cb_conf_bus[258] ),
    .CLK(clknet_7_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09622_ (.D(_02559_),
    .Q(\cb_east.inst.cb_conf_bus[259] ),
    .CLK(clknet_7_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09623_ (.D(_02561_),
    .Q(\cb_east.inst.cb_conf_bus[260] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09624_ (.D(_02563_),
    .Q(\cb_east.inst.cb_conf_bus[261] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09625_ (.D(_02565_),
    .Q(\cb_east.inst.cb_conf_bus[262] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09626_ (.D(_02567_),
    .Q(\cb_east.inst.cb_conf_bus[263] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09627_ (.D(_02569_),
    .Q(\cb_east.inst.cb_conf_bus[264] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09628_ (.D(_02571_),
    .Q(\cb_east.inst.cb_conf_bus[265] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09629_ (.D(_02573_),
    .Q(\cb_east.inst.cb_conf_bus[266] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09630_ (.D(_02575_),
    .Q(\cb_east.inst.cb_conf_bus[267] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09631_ (.D(_02577_),
    .Q(\cb_east.inst.cb_conf_bus[268] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09632_ (.D(_02579_),
    .Q(\cb_east.inst.cb_conf_bus[269] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09633_ (.D(_02581_),
    .Q(\cb_east.inst.cb_conf_bus[270] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09634_ (.D(_02583_),
    .Q(\cb_east.inst.cb_conf_bus[271] ),
    .CLK(clknet_7_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09635_ (.D(_02585_),
    .Q(\cb_east.inst.cb_conf_bus[272] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09636_ (.D(_02587_),
    .Q(\cb_east.inst.cb_conf_bus[273] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09637_ (.D(_02589_),
    .Q(\cb_east.inst.cb_conf_bus[274] ),
    .CLK(clknet_7_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09638_ (.D(_02591_),
    .Q(\cb_east.inst.cb_conf_bus[275] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09639_ (.D(_02593_),
    .Q(\cb_east.inst.cb_conf_bus[276] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09640_ (.D(_02595_),
    .Q(\cb_east.inst.cb_conf_bus[277] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09641_ (.D(_02597_),
    .Q(\cb_east.inst.cb_conf_bus[278] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09642_ (.D(_02599_),
    .Q(\cb_east.inst.cb_conf_bus[279] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09643_ (.D(_02601_),
    .Q(\cb_east.inst.cb_conf_bus[280] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09644_ (.D(_02603_),
    .Q(\cb_east.inst.cb_conf_bus[281] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09645_ (.D(_02605_),
    .Q(\cb_east.inst.cb_conf_bus[282] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09646_ (.D(_02607_),
    .Q(\cb_east.inst.cb_conf_bus[283] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09647_ (.D(_02609_),
    .Q(\cb_east.inst.cb_conf_bus[284] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09648_ (.D(_02611_),
    .Q(\cb_east.inst.cb_conf_bus[285] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09649_ (.D(_02613_),
    .Q(\cb_east.inst.cb_conf_bus[286] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09650_ (.D(_02615_),
    .Q(\cb_east.inst.cb_conf_bus[287] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09651_ (.D(_02617_),
    .Q(\cb_east.inst.cb_conf_bus[288] ),
    .CLK(clknet_7_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09652_ (.D(_02619_),
    .Q(\cb_east.inst.cb_conf_bus[289] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09653_ (.D(_02621_),
    .Q(\cb_east.inst.cb_conf_bus[290] ),
    .CLK(clknet_7_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09654_ (.D(_02623_),
    .Q(\cb_east.inst.cb_conf_bus[291] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09655_ (.D(_02625_),
    .Q(\cb_east.inst.cb_conf_bus[292] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09656_ (.D(_02627_),
    .Q(\cb_east.inst.cb_conf_bus[293] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09657_ (.D(_02629_),
    .Q(\cb_east.inst.cb_conf_bus[294] ),
    .CLK(clknet_7_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09658_ (.D(_02631_),
    .Q(\cb_east.inst.cb_conf_bus[295] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09659_ (.D(_02633_),
    .Q(\cb_east.inst.cb_conf_bus[296] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09660_ (.D(_02635_),
    .Q(\cb_east.inst.cb_conf_bus[297] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09661_ (.D(_02637_),
    .Q(\cb_east.inst.cb_conf_bus[298] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09662_ (.D(_02639_),
    .Q(\cb_east.inst.cb_conf_bus[299] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09663_ (.D(_02641_),
    .Q(\cb_east.inst.cb_conf_bus[300] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09664_ (.D(_02643_),
    .Q(\cb_east.inst.cb_conf_bus[301] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09665_ (.D(_02645_),
    .Q(\cb_east.inst.cb_conf_bus[302] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09666_ (.D(_02647_),
    .Q(\cb_east.inst.cb_conf_bus[303] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09667_ (.D(_02649_),
    .Q(\cb_east.inst.cb_conf_bus[304] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09668_ (.D(_02651_),
    .Q(\cb_east.inst.cb_conf_bus[305] ),
    .CLK(clknet_7_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09669_ (.D(_02653_),
    .Q(\cb_east.inst.cb_conf_bus[306] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09670_ (.D(_02655_),
    .Q(\cb_east.inst.cb_conf_bus[307] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09671_ (.D(_02657_),
    .Q(\cb_east.inst.cb_conf_bus[308] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09672_ (.D(_02659_),
    .Q(\cb_east.inst.cb_conf_bus[309] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09673_ (.D(_02661_),
    .Q(\cb_east.inst.cb_conf_bus[310] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09674_ (.D(_02663_),
    .Q(\cb_east.inst.cb_conf_bus[311] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09675_ (.D(_02665_),
    .Q(\cb_east.inst.cb_conf_bus[312] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09676_ (.D(_02667_),
    .Q(\cb_east.inst.cb_conf_bus[313] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09677_ (.D(_02669_),
    .Q(\cb_east.inst.cb_conf_bus[314] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09678_ (.D(_02671_),
    .Q(\cb_east.inst.cb_conf_bus[315] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09679_ (.D(_02673_),
    .Q(\cb_east.inst.cb_conf_bus[316] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09680_ (.D(_02675_),
    .Q(\cb_east.inst.cb_conf_bus[317] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09681_ (.D(_02677_),
    .Q(\cb_east.inst.cb_conf_bus[318] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09682_ (.D(_02679_),
    .Q(\cb_east.inst.cb_conf_bus[319] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09683_ (.D(_02681_),
    .Q(\cb_east.inst.cb_conf_bus[320] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09684_ (.D(_02683_),
    .Q(\cb_east.inst.cb_conf_bus[321] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09685_ (.D(_02685_),
    .Q(\cb_east.inst.cb_conf_bus[322] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09686_ (.D(_02687_),
    .Q(\cb_east.inst.cb_conf_bus[323] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09687_ (.D(_02689_),
    .Q(\cb_east.inst.cb_conf_bus[324] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09688_ (.D(_02691_),
    .Q(\cb_east.inst.cb_conf_bus[325] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09689_ (.D(_02693_),
    .Q(\cb_east.inst.cb_conf_bus[326] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09690_ (.D(_02695_),
    .Q(\cb_east.inst.cb_conf_bus[327] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09691_ (.D(_02697_),
    .Q(\cb_east.inst.cb_conf_bus[328] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09692_ (.D(_02699_),
    .Q(\cb_east.inst.cb_conf_bus[329] ),
    .CLK(clknet_7_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09693_ (.D(_02701_),
    .Q(\cb_east.inst.cb_conf_bus[330] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09694_ (.D(_02703_),
    .Q(\cb_east.inst.cb_conf_bus[331] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09695_ (.D(_02705_),
    .Q(\cb_east.inst.cb_conf_bus[332] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09696_ (.D(_02707_),
    .Q(\cb_east.inst.cb_conf_bus[333] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09697_ (.D(_02709_),
    .Q(\cb_east.inst.cb_conf_bus[334] ),
    .CLK(clknet_7_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09698_ (.D(_02711_),
    .Q(\cb_east.inst.cb_conf_bus[335] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09699_ (.D(_02713_),
    .Q(\cb_east.inst.cb_conf_bus[336] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09700_ (.D(_02715_),
    .Q(\cb_east.inst.cb_conf_bus[337] ),
    .CLK(clknet_7_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09701_ (.D(_02717_),
    .Q(\cb_east.inst.cb_conf_bus[338] ),
    .CLK(clknet_7_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09702_ (.D(_02719_),
    .Q(\cb_east.inst.cb_conf_bus[339] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09703_ (.D(_02721_),
    .Q(\cb_east.inst.cb_conf_bus[340] ),
    .CLK(clknet_7_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09704_ (.D(_02723_),
    .Q(\cb_east.inst.cb_conf_bus[341] ),
    .CLK(clknet_7_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09705_ (.D(_02725_),
    .Q(\cb_east.inst.cb_conf_bus[342] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09706_ (.D(_02727_),
    .Q(\cb_east.inst.cb_conf_bus[343] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09707_ (.D(_02729_),
    .Q(\cb_east.inst.cb_conf_bus[344] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09708_ (.D(_02731_),
    .Q(\cb_east.inst.cb_conf_bus[345] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09709_ (.D(_02733_),
    .Q(\cb_east.inst.cb_conf_bus[346] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09710_ (.D(_02735_),
    .Q(\cb_east.inst.cb_conf_bus[347] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09711_ (.D(_02737_),
    .Q(\cb_east.inst.cb_conf_bus[348] ),
    .CLK(clknet_7_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09712_ (.D(_02739_),
    .Q(\cb_east.inst.cb_conf_bus[349] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09713_ (.D(_02741_),
    .Q(\cb_east.inst.cb_conf_bus[350] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09714_ (.D(_02743_),
    .Q(\cb_east.inst.cb_conf_bus[351] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09715_ (.D(_02745_),
    .Q(\cb_east.inst.cb_conf_bus[352] ),
    .CLK(clknet_7_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09716_ (.D(_02747_),
    .Q(\cb_east.inst.cb_conf_bus[353] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09717_ (.D(_02749_),
    .Q(\cb_east.inst.cb_conf_bus[354] ),
    .CLK(clknet_7_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09718_ (.D(_02751_),
    .Q(\cb_east.inst.cb_conf_bus[355] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09719_ (.D(_02753_),
    .Q(\cb_east.inst.cb_conf_bus[356] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09720_ (.D(_02755_),
    .Q(\cb_east.inst.cb_conf_bus[357] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09721_ (.D(_02757_),
    .Q(\cb_east.inst.cb_conf_bus[358] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09722_ (.D(_02759_),
    .Q(\cb_east.inst.cb_conf_bus[359] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09723_ (.D(_02761_),
    .Q(\cb_east.inst.cb_conf_bus[360] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09724_ (.D(_02763_),
    .Q(\cb_east.inst.cb_conf_bus[361] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09725_ (.D(_02765_),
    .Q(\cb_east.inst.cb_conf_bus[362] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09726_ (.D(_02767_),
    .Q(\cb_east.inst.cb_conf_bus[363] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09727_ (.D(_02769_),
    .Q(\cb_east.inst.cb_conf_bus[364] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09728_ (.D(_02771_),
    .Q(\cb_east.inst.cb_conf_bus[365] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09729_ (.D(_02773_),
    .Q(\cb_east.inst.cb_conf_bus[366] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09730_ (.D(_02775_),
    .Q(\cb_east.inst.cb_conf_bus[367] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09731_ (.D(_02777_),
    .Q(\cb_east.inst.cb_conf_bus[368] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09732_ (.D(_02779_),
    .Q(\cb_east.inst.cb_conf_bus[369] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09733_ (.D(_02781_),
    .Q(\cb_east.inst.cb_conf_bus[370] ),
    .CLK(clknet_7_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09734_ (.D(_02783_),
    .Q(\cb_east.inst.cb_conf_bus[371] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09735_ (.D(_02785_),
    .Q(\cb_east.inst.cb_conf_bus[372] ),
    .CLK(clknet_7_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09736_ (.D(_02787_),
    .Q(\cb_east.inst.cb_conf_bus[373] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09737_ (.D(_02789_),
    .Q(\cb_east.inst.cb_conf_bus[374] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09738_ (.D(_02791_),
    .Q(\cb_east.inst.cb_conf_bus[375] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09739_ (.D(_02793_),
    .Q(\cb_east.inst.cb_conf_bus[376] ),
    .CLK(clknet_7_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09740_ (.D(_02795_),
    .Q(\cb_east.inst.cb_conf_bus[377] ),
    .CLK(clknet_7_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09741_ (.D(_02797_),
    .Q(\cb_east.inst.cb_conf_bus[378] ),
    .CLK(clknet_7_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09742_ (.D(_02799_),
    .Q(\cb_east.inst.cb_conf_bus[379] ),
    .CLK(clknet_7_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09743_ (.D(_02801_),
    .Q(\cb_east.inst.cb_conf_bus[380] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09744_ (.D(_02803_),
    .Q(\cb_east.inst.cb_conf_bus[381] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09745_ (.D(_02805_),
    .Q(\cb_east.inst.cb_conf_bus[382] ),
    .CLK(clknet_7_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09746_ (.D(_02807_),
    .Q(\cb_east.inst.cb_conf_bus[383] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09747_ (.D(_02809_),
    .Q(\cb_east.inst.cb_conf_bus[384] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09748_ (.D(_02811_),
    .Q(\cb_east.inst.cb_conf_bus[385] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09749_ (.D(_02813_),
    .Q(\cb_east.inst.cb_conf_bus[386] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09750_ (.D(_02815_),
    .Q(\cb_east.inst.cb_conf_bus[387] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09751_ (.D(_02817_),
    .Q(\cb_east.inst.cb_conf_bus[388] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09752_ (.D(_02819_),
    .Q(\cb_east.inst.cb_conf_bus[389] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09753_ (.D(_02821_),
    .Q(\cb_east.inst.cb_conf_bus[390] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09754_ (.D(_02823_),
    .Q(\cb_east.inst.cb_conf_bus[391] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09755_ (.D(_02825_),
    .Q(\cb_east.inst.cb_conf_bus[392] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09756_ (.D(_02827_),
    .Q(\cb_east.inst.cb_conf_bus[393] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09757_ (.D(_02829_),
    .Q(\cb_east.inst.cb_conf_bus[394] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09758_ (.D(_02831_),
    .Q(\cb_east.inst.cb_conf_bus[395] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09759_ (.D(_02833_),
    .Q(\cb_east.inst.cb_conf_bus[396] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09760_ (.D(_02835_),
    .Q(\cb_east.inst.cb_conf_bus[397] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09761_ (.D(_02837_),
    .Q(\cb_east.inst.cb_conf_bus[398] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09762_ (.D(_02839_),
    .Q(\cb_east.inst.cb_conf_bus[399] ),
    .CLK(clknet_7_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09763_ (.D(_02841_),
    .Q(\cb_east.inst.cb_conf_bus[400] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09764_ (.D(_02843_),
    .Q(\cb_east.inst.cb_conf_bus[401] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09765_ (.D(_02845_),
    .Q(\cb_east.inst.cb_conf_bus[402] ),
    .CLK(clknet_7_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09766_ (.D(_02847_),
    .Q(\cb_east.inst.cb_conf_bus[403] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09767_ (.D(_02849_),
    .Q(\cb_east.inst.cb_conf_bus[404] ),
    .CLK(clknet_7_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09768_ (.D(_02851_),
    .Q(\cb_east.inst.cb_conf_bus[405] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09769_ (.D(_02853_),
    .Q(\cb_east.inst.cb_conf_bus[406] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09770_ (.D(_02855_),
    .Q(\cb_east.inst.cb_conf_bus[407] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09771_ (.D(_02857_),
    .Q(\cb_east.inst.cb_conf_bus[408] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09772_ (.D(_02859_),
    .Q(\cb_east.inst.cb_conf_bus[409] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09773_ (.D(_02861_),
    .Q(\cb_east.inst.cb_conf_bus[410] ),
    .CLK(clknet_7_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09774_ (.D(_02863_),
    .Q(\cb_east.inst.cb_conf_bus[411] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09775_ (.D(_02865_),
    .Q(\cb_east.inst.cb_conf_bus[412] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09776_ (.D(_02867_),
    .Q(\cb_east.inst.cb_conf_bus[413] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09777_ (.D(_02869_),
    .Q(\cb_east.inst.cb_conf_bus[414] ),
    .CLK(clknet_7_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09778_ (.D(_02871_),
    .Q(\cb_east.inst.cb_conf_bus[415] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09779_ (.D(_02873_),
    .Q(\cb_east.inst.cb_conf_bus[416] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09780_ (.D(_02875_),
    .Q(\cb_east.inst.cb_conf_bus[417] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09781_ (.D(_02877_),
    .Q(\cb_east.inst.cb_conf_bus[418] ),
    .CLK(clknet_7_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09782_ (.D(_02879_),
    .Q(\cb_east.inst.cb_conf_bus[419] ),
    .CLK(clknet_7_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09783_ (.D(_02881_),
    .Q(\cb_east.inst.configuroni.comb_shifter.config_data[420] ),
    .CLK(clknet_7_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09784_ (.D(_02883_),
    .Q(\sb.configuroni.comb_shifter.config_data[48] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09785_ (.D(_02885_),
    .Q(\sb.configuroni.comb_config[47] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09786_ (.D(_02887_),
    .Q(\sb.configuroni.comb_config[46] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09787_ (.D(_02889_),
    .Q(\sb.configuroni.comb_config[45] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09788_ (.D(_02891_),
    .Q(\sb.configuroni.comb_config[44] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09789_ (.D(_02893_),
    .Q(\sb.configuroni.comb_config[43] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09790_ (.D(_02895_),
    .Q(\sb.configuroni.comb_config[42] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09791_ (.D(_02897_),
    .Q(\sb.configuroni.comb_config[41] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09792_ (.D(_02899_),
    .Q(\sb.configuroni.comb_config[40] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09793_ (.D(_02901_),
    .Q(\sb.configuroni.comb_config[39] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09794_ (.D(_02903_),
    .Q(\sb.configuroni.comb_config[38] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09795_ (.D(_02905_),
    .Q(\sb.configuroni.comb_config[37] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09796_ (.D(_02907_),
    .Q(\sb.configuroni.comb_config[36] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09797_ (.D(_02909_),
    .Q(\sb.configuroni.comb_config[35] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09798_ (.D(_02911_),
    .Q(\sb.configuroni.comb_config[34] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09799_ (.D(_02913_),
    .Q(\sb.configuroni.comb_config[33] ),
    .CLK(clknet_7_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09800_ (.D(_02915_),
    .Q(\sb.configuroni.comb_config[32] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09801_ (.D(_02917_),
    .Q(\sb.configuroni.comb_config[31] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09802_ (.D(_02919_),
    .Q(\sb.configuroni.comb_config[30] ),
    .CLK(clknet_7_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09803_ (.D(_02921_),
    .Q(\sb.configuroni.comb_config[29] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09804_ (.D(_02923_),
    .Q(\sb.configuroni.comb_config[28] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09805_ (.D(_02925_),
    .Q(\sb.configuroni.comb_config[27] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09806_ (.D(_02927_),
    .Q(\sb.configuroni.comb_config[26] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09807_ (.D(_02929_),
    .Q(\sb.configuroni.comb_config[25] ),
    .CLK(clknet_7_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09808_ (.D(_02931_),
    .Q(\sb.configuroni.comb_config[24] ),
    .CLK(clknet_7_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09809_ (.D(_02933_),
    .Q(\sb.configuroni.comb_config[23] ),
    .CLK(clknet_7_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09810_ (.D(_02935_),
    .Q(\sb.configuroni.comb_config[22] ),
    .CLK(clknet_7_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09811_ (.D(_02937_),
    .Q(\sb.configuroni.comb_config[21] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09812_ (.D(_02939_),
    .Q(\sb.configuroni.comb_config[20] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09813_ (.D(_02941_),
    .Q(\sb.configuroni.comb_config[19] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09814_ (.D(_02943_),
    .Q(\sb.configuroni.comb_config[18] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09815_ (.D(_02945_),
    .Q(\sb.configuroni.comb_config[17] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09816_ (.D(_02947_),
    .Q(\sb.configuroni.comb_config[16] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09817_ (.D(_02949_),
    .Q(\sb.configuroni.comb_config[15] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09818_ (.D(_02951_),
    .Q(\sb.configuroni.comb_config[14] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09819_ (.D(_02953_),
    .Q(\sb.configuroni.comb_config[13] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09820_ (.D(_02955_),
    .Q(\sb.configuroni.comb_config[12] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09821_ (.D(_02957_),
    .Q(\sb.configuroni.comb_config[11] ),
    .CLK(clknet_7_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09822_ (.D(_02959_),
    .Q(\sb.configuroni.comb_config[10] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09823_ (.D(_02961_),
    .Q(\sb.configuroni.comb_config[9] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09824_ (.D(_02963_),
    .Q(\sb.configuroni.comb_config[8] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09825_ (.D(_02965_),
    .Q(\sb.configuroni.comb_config[7] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09826_ (.D(_02967_),
    .Q(\sb.configuroni.comb_config[6] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09827_ (.D(_02969_),
    .Q(\sb.configuroni.comb_config[5] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09828_ (.D(_02971_),
    .Q(\sb.configuroni.comb_config[4] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09829_ (.D(_02973_),
    .Q(\sb.configuroni.comb_config[3] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09830_ (.D(_02975_),
    .Q(\sb.configuroni.comb_config[2] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09831_ (.D(_02977_),
    .Q(\sb.configuroni.comb_config[1] ),
    .CLK(clknet_7_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09832_ (.D(_02979_),
    .Q(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .CLK(clknet_7_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09833_ (.D(_02981_),
    .Q(\sb.configuroni.comb_shifter.config_data[49] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09834_ (.D(_02983_),
    .Q(\slice.configuroni.mem_ctrl ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09835_ (.D(_02985_),
    .Q(\slice.configuroni.input_mux ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09836_ (.D(_02987_),
    .Q(\slice.configuroni.comb_shifter.config_data[135] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09837_ (.D(_02989_),
    .Q(\slice.configuroni.comb_config[134] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09838_ (.D(_02991_),
    .Q(\slice.configuroni.comb_config[133] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09839_ (.D(_02993_),
    .Q(\slice.configuroni.comb_config[132] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09840_ (.D(_02995_),
    .Q(\slice.configuroni.comb_config[131] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09841_ (.D(_02997_),
    .Q(\slice.configuroni.comb_config[130] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09842_ (.D(_02999_),
    .Q(\slice.configuroni.comb_config[129] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09843_ (.D(_03001_),
    .Q(\slice.configuroni.comb_config[128] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09844_ (.D(_03003_),
    .Q(\slice.configuroni.comb_config[127] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09845_ (.D(_03005_),
    .Q(\slice.configuroni.comb_config[126] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09846_ (.D(_03007_),
    .Q(\slice.configuroni.comb_config[125] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09847_ (.D(_03009_),
    .Q(\slice.configuroni.comb_config[124] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09848_ (.D(_03011_),
    .Q(\slice.configuroni.comb_config[123] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09849_ (.D(_03013_),
    .Q(\slice.configuroni.comb_config[122] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09850_ (.D(_03015_),
    .Q(\slice.configuroni.comb_config[121] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09851_ (.D(_03017_),
    .Q(\slice.configuroni.comb_config[120] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09852_ (.D(_03019_),
    .Q(\slice.configuroni.comb_config[119] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09853_ (.D(_03021_),
    .Q(\slice.configuroni.comb_config[118] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09854_ (.D(_03023_),
    .Q(\slice.configuroni.comb_config[117] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09855_ (.D(_03025_),
    .Q(\slice.configuroni.comb_config[116] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09856_ (.D(_03027_),
    .Q(\slice.configuroni.comb_config[115] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09857_ (.D(_03029_),
    .Q(\slice.configuroni.comb_config[114] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09858_ (.D(_03031_),
    .Q(\slice.configuroni.comb_config[113] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09859_ (.D(_03033_),
    .Q(\slice.configuroni.comb_config[112] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09860_ (.D(_03035_),
    .Q(\slice.configuroni.comb_config[111] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09861_ (.D(_03037_),
    .Q(\slice.configuroni.comb_config[110] ),
    .CLK(clknet_7_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09862_ (.D(_03039_),
    .Q(\slice.configuroni.comb_config[109] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09863_ (.D(_03041_),
    .Q(\slice.configuroni.comb_config[108] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09864_ (.D(_03043_),
    .Q(\slice.configuroni.comb_config[107] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09865_ (.D(_03045_),
    .Q(\slice.configuroni.comb_config[106] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09866_ (.D(_03047_),
    .Q(\slice.configuroni.comb_config[105] ),
    .CLK(clknet_7_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09867_ (.D(_03049_),
    .Q(\slice.configuroni.comb_config[104] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09868_ (.D(_03051_),
    .Q(\slice.configuroni.comb_config[103] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09869_ (.D(_03053_),
    .Q(\slice.configuroni.comb_config[102] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09870_ (.D(_03055_),
    .Q(\slice.configuroni.comb_config[101] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09871_ (.D(_03057_),
    .Q(\slice.configuroni.comb_config[100] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09872_ (.D(_03059_),
    .Q(\slice.configuroni.comb_config[99] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09873_ (.D(_03061_),
    .Q(\slice.configuroni.comb_config[98] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09874_ (.D(_03063_),
    .Q(\slice.configuroni.comb_config[97] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09875_ (.D(_03065_),
    .Q(\slice.configuroni.comb_config[96] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09876_ (.D(_03067_),
    .Q(\slice.configuroni.comb_config[95] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09877_ (.D(_03069_),
    .Q(\slice.configuroni.comb_config[94] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09878_ (.D(_03071_),
    .Q(\slice.configuroni.comb_config[93] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09879_ (.D(_03073_),
    .Q(\slice.configuroni.comb_config[92] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09880_ (.D(_03075_),
    .Q(\slice.configuroni.comb_config[91] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09881_ (.D(_03077_),
    .Q(\slice.configuroni.comb_config[90] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09882_ (.D(_03079_),
    .Q(\slice.configuroni.comb_config[89] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09883_ (.D(_03081_),
    .Q(\slice.configuroni.comb_config[88] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09884_ (.D(_03083_),
    .Q(\slice.configuroni.comb_config[87] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09885_ (.D(_03085_),
    .Q(\slice.configuroni.comb_config[86] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09886_ (.D(_03087_),
    .Q(\slice.configuroni.comb_config[85] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09887_ (.D(_03089_),
    .Q(\slice.configuroni.comb_config[84] ),
    .CLK(clknet_7_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09888_ (.D(_03091_),
    .Q(\slice.configuroni.comb_config[83] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09889_ (.D(_03093_),
    .Q(\slice.configuroni.comb_config[82] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09890_ (.D(_03095_),
    .Q(\slice.configuroni.comb_config[81] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09891_ (.D(_03097_),
    .Q(\slice.configuroni.comb_config[80] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09892_ (.D(_03099_),
    .Q(\slice.configuroni.comb_config[79] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09893_ (.D(_03101_),
    .Q(\slice.configuroni.comb_config[78] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09894_ (.D(_03103_),
    .Q(\slice.configuroni.comb_config[77] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09895_ (.D(_03105_),
    .Q(\slice.configuroni.comb_config[76] ),
    .CLK(clknet_7_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09896_ (.D(_03107_),
    .Q(\slice.configuroni.comb_config[75] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09897_ (.D(_03109_),
    .Q(\slice.configuroni.comb_config[74] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09898_ (.D(_03111_),
    .Q(\slice.configuroni.comb_config[73] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09899_ (.D(_03113_),
    .Q(\slice.configuroni.comb_config[72] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09900_ (.D(_03115_),
    .Q(\slice.configuroni.comb_config[71] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09901_ (.D(_03117_),
    .Q(\slice.configuroni.comb_config[70] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09902_ (.D(_03119_),
    .Q(\slice.configuroni.comb_config[69] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09903_ (.D(_03121_),
    .Q(\slice.configuroni.comb_config[68] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09904_ (.D(_03123_),
    .Q(\slice.configuroni.comb_config[67] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09905_ (.D(_03125_),
    .Q(\slice.configuroni.comb_config[66] ),
    .CLK(clknet_7_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09906_ (.D(_03127_),
    .Q(\slice.configuroni.comb_config[65] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09907_ (.D(_03129_),
    .Q(\slice.configuroni.comb_config[64] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09908_ (.D(_03131_),
    .Q(\slice.configuroni.comb_config[63] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09909_ (.D(_03133_),
    .Q(\slice.configuroni.comb_config[62] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09910_ (.D(_03135_),
    .Q(\slice.configuroni.comb_config[61] ),
    .CLK(clknet_7_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09911_ (.D(_03137_),
    .Q(\slice.configuroni.comb_config[60] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09912_ (.D(_03139_),
    .Q(\slice.configuroni.comb_config[59] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09913_ (.D(_03141_),
    .Q(\slice.configuroni.comb_config[58] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09914_ (.D(_03143_),
    .Q(\slice.configuroni.comb_config[57] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09915_ (.D(_03145_),
    .Q(\slice.configuroni.comb_config[56] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09916_ (.D(_03147_),
    .Q(\slice.configuroni.comb_config[55] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09917_ (.D(_03149_),
    .Q(\slice.configuroni.comb_config[54] ),
    .CLK(clknet_7_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09918_ (.D(_03151_),
    .Q(\slice.configuroni.comb_config[53] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09919_ (.D(_03153_),
    .Q(\slice.configuroni.comb_config[52] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09920_ (.D(_03155_),
    .Q(\slice.configuroni.comb_config[51] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09921_ (.D(_03157_),
    .Q(\slice.configuroni.comb_config[50] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09922_ (.D(_03159_),
    .Q(\slice.configuroni.comb_config[49] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09923_ (.D(_03161_),
    .Q(\slice.configuroni.comb_config[48] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09924_ (.D(_03163_),
    .Q(\slice.configuroni.comb_config[47] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09925_ (.D(_03165_),
    .Q(\slice.configuroni.comb_config[46] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09926_ (.D(_03167_),
    .Q(\slice.configuroni.comb_config[45] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09927_ (.D(_03169_),
    .Q(\slice.configuroni.comb_config[44] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09928_ (.D(_03171_),
    .Q(\slice.configuroni.comb_config[43] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09929_ (.D(_03173_),
    .Q(\slice.configuroni.comb_config[42] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09930_ (.D(_03175_),
    .Q(\slice.configuroni.comb_config[41] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09931_ (.D(_03177_),
    .Q(\slice.configuroni.comb_config[40] ),
    .CLK(clknet_7_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09932_ (.D(_03179_),
    .Q(\slice.configuroni.comb_config[39] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09933_ (.D(_03181_),
    .Q(\slice.configuroni.comb_config[38] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09934_ (.D(_03183_),
    .Q(\slice.configuroni.comb_config[37] ),
    .CLK(clknet_7_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09935_ (.D(_03185_),
    .Q(\slice.configuroni.comb_config[36] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09936_ (.D(_03187_),
    .Q(\slice.configuroni.comb_config[35] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09937_ (.D(_03189_),
    .Q(\slice.configuroni.comb_config[34] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09938_ (.D(_03191_),
    .Q(\slice.configuroni.comb_config[33] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09939_ (.D(_03193_),
    .Q(\slice.configuroni.comb_config[32] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09940_ (.D(_03195_),
    .Q(\slice.configuroni.comb_config[31] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09941_ (.D(_03197_),
    .Q(\slice.configuroni.comb_config[30] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09942_ (.D(_03199_),
    .Q(\slice.configuroni.comb_config[29] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09943_ (.D(_03201_),
    .Q(\slice.configuroni.comb_config[28] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09944_ (.D(_03203_),
    .Q(\slice.configuroni.comb_config[27] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09945_ (.D(_03205_),
    .Q(\slice.configuroni.comb_config[26] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09946_ (.D(_03207_),
    .Q(\slice.configuroni.comb_config[25] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09947_ (.D(_03209_),
    .Q(\slice.configuroni.comb_config[24] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09948_ (.D(_03211_),
    .Q(\slice.configuroni.comb_config[23] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09949_ (.D(_03213_),
    .Q(\slice.configuroni.comb_config[22] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09950_ (.D(_03215_),
    .Q(\slice.configuroni.comb_config[21] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09951_ (.D(_03217_),
    .Q(\slice.configuroni.comb_config[20] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09952_ (.D(_03219_),
    .Q(\slice.configuroni.comb_config[19] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09953_ (.D(_03221_),
    .Q(\slice.configuroni.comb_config[18] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09954_ (.D(_03223_),
    .Q(\slice.configuroni.comb_config[17] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09955_ (.D(_03225_),
    .Q(\slice.configuroni.comb_config[16] ),
    .CLK(clknet_7_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09956_ (.D(_03227_),
    .Q(\slice.configuroni.comb_config[15] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09957_ (.D(_03229_),
    .Q(\slice.configuroni.comb_config[14] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09958_ (.D(_03231_),
    .Q(\slice.configuroni.comb_config[13] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09959_ (.D(_03233_),
    .Q(\slice.configuroni.comb_config[12] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09960_ (.D(_03235_),
    .Q(\slice.configuroni.comb_config[11] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09961_ (.D(_03237_),
    .Q(\slice.configuroni.comb_config[10] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09962_ (.D(_03239_),
    .Q(\slice.configuroni.comb_config[9] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09963_ (.D(_03241_),
    .Q(\slice.configuroni.comb_config[8] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09964_ (.D(_03243_),
    .Q(\slice.configuroni.comb_config[7] ),
    .CLK(clknet_7_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09965_ (.D(_03245_),
    .Q(\slice.configuroni.comb_config[6] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09966_ (.D(_03247_),
    .Q(\slice.configuroni.comb_config[5] ),
    .CLK(clknet_7_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09967_ (.D(_03249_),
    .Q(\slice.configuroni.comb_config[4] ),
    .CLK(clknet_7_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09968_ (.D(_03251_),
    .Q(\slice.configuroni.comb_config[3] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09969_ (.D(_03253_),
    .Q(\slice.configuroni.comb_config[2] ),
    .CLK(clknet_7_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09970_ (.D(_03255_),
    .Q(\slice.configuroni.comb_config[1] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09971_ (.D(_03257_),
    .Q(\slice.configuroni.comb_config[0] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09972_ (.D(_03259_),
    .Q(\slice.configuroni.comb_shifter.config_data[136] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09973_ (.D(_03261_),
    .Q(\slice.configuroni.mem_config[6] ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09974_ (.D(_03263_),
    .Q(\slice.configuroni.mem_config[5] ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09975_ (.D(_03265_),
    .Q(\slice.configuroni.mem_config[4] ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09976_ (.D(_03267_),
    .Q(\slice.configuroni.mem_config[3] ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09977_ (.D(_03269_),
    .Q(\slice.configuroni.mem_config[2] ),
    .CLK(clknet_7_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09978_ (.D(_03271_),
    .Q(\slice.configuroni.mem_config[1] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09979_ (.D(_03273_),
    .Q(\cb_north.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09980_ (.D(_03275_),
    .Q(\slice.configuroni.mem_config[7] ),
    .CLK(clknet_7_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09981_ (.D(_03277_),
    .Q(\cb_north.inst.configuroni.comb_shifter.config_data[421] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09982_ (.D(_03279_),
    .Q(\cb_north.inst.cb_conf_bus[0] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09983_ (.D(_03281_),
    .Q(\cb_north.inst.cb_conf_bus[1] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09984_ (.D(_03283_),
    .Q(\cb_north.inst.cb_conf_bus[2] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09985_ (.D(_03285_),
    .Q(\cb_north.inst.cb_conf_bus[3] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09986_ (.D(_03287_),
    .Q(\cb_north.inst.cb_conf_bus[4] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09987_ (.D(_03289_),
    .Q(\cb_north.inst.cb_conf_bus[5] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09988_ (.D(_03291_),
    .Q(\cb_north.inst.cb_conf_bus[6] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09989_ (.D(_03293_),
    .Q(\cb_north.inst.cb_conf_bus[7] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09990_ (.D(_03295_),
    .Q(\cb_north.inst.cb_conf_bus[8] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09991_ (.D(_03297_),
    .Q(\cb_north.inst.cb_conf_bus[9] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09992_ (.D(_03299_),
    .Q(\cb_north.inst.cb_conf_bus[10] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09993_ (.D(_03301_),
    .Q(\cb_north.inst.cb_conf_bus[11] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09994_ (.D(_03303_),
    .Q(\cb_north.inst.cb_conf_bus[12] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09995_ (.D(_03305_),
    .Q(\cb_north.inst.cb_conf_bus[13] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09996_ (.D(_03307_),
    .Q(\cb_north.inst.cb_conf_bus[14] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09997_ (.D(_03309_),
    .Q(\cb_north.inst.cb_conf_bus[15] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09998_ (.D(_03311_),
    .Q(\cb_north.inst.cb_conf_bus[16] ),
    .CLK(clknet_7_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _09999_ (.D(_03313_),
    .Q(\cb_north.inst.cb_conf_bus[17] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10000_ (.D(_03315_),
    .Q(\cb_north.inst.cb_conf_bus[18] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10001_ (.D(_03317_),
    .Q(\cb_north.inst.cb_conf_bus[19] ),
    .CLK(clknet_7_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10002_ (.D(_03319_),
    .Q(\cb_north.inst.cb_conf_bus[20] ),
    .CLK(clknet_7_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10003_ (.D(_03321_),
    .Q(\cb_north.inst.cb_conf_bus[21] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10004_ (.D(_03323_),
    .Q(\cb_north.inst.cb_conf_bus[22] ),
    .CLK(clknet_7_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10005_ (.D(_03325_),
    .Q(\cb_north.inst.cb_conf_bus[23] ),
    .CLK(clknet_7_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10006_ (.D(_03327_),
    .Q(\cb_north.inst.cb_conf_bus[24] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10007_ (.D(_03329_),
    .Q(\cb_north.inst.cb_conf_bus[25] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10008_ (.D(_03331_),
    .Q(\cb_north.inst.cb_conf_bus[26] ),
    .CLK(clknet_7_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10009_ (.D(_03333_),
    .Q(\cb_north.inst.cb_conf_bus[27] ),
    .CLK(clknet_7_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10010_ (.D(_03335_),
    .Q(\cb_north.inst.cb_conf_bus[28] ),
    .CLK(clknet_7_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10011_ (.D(_03337_),
    .Q(\cb_north.inst.cb_conf_bus[29] ),
    .CLK(clknet_7_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10012_ (.D(_03339_),
    .Q(\cb_north.inst.cb_conf_bus[30] ),
    .CLK(clknet_7_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10013_ (.D(_03341_),
    .Q(\cb_north.inst.cb_conf_bus[31] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10014_ (.D(_03343_),
    .Q(\cb_north.inst.cb_conf_bus[32] ),
    .CLK(clknet_7_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10015_ (.D(_03345_),
    .Q(\cb_north.inst.cb_conf_bus[33] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10016_ (.D(_03347_),
    .Q(\cb_north.inst.cb_conf_bus[34] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10017_ (.D(_03349_),
    .Q(\cb_north.inst.cb_conf_bus[35] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10018_ (.D(_03351_),
    .Q(\cb_north.inst.cb_conf_bus[36] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10019_ (.D(_03353_),
    .Q(\cb_north.inst.cb_conf_bus[37] ),
    .CLK(clknet_7_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10020_ (.D(_03355_),
    .Q(\cb_north.inst.cb_conf_bus[38] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10021_ (.D(_03357_),
    .Q(\cb_north.inst.cb_conf_bus[39] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10022_ (.D(_03359_),
    .Q(\cb_north.inst.cb_conf_bus[40] ),
    .CLK(clknet_7_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10023_ (.D(_03361_),
    .Q(\cb_north.inst.cb_conf_bus[41] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10024_ (.D(_03363_),
    .Q(\cb_north.inst.cb_conf_bus[42] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10025_ (.D(_03365_),
    .Q(\cb_north.inst.cb_conf_bus[43] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10026_ (.D(_03367_),
    .Q(\cb_north.inst.cb_conf_bus[44] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10027_ (.D(_03369_),
    .Q(\cb_north.inst.cb_conf_bus[45] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10028_ (.D(_03371_),
    .Q(\cb_north.inst.cb_conf_bus[46] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10029_ (.D(_03373_),
    .Q(\cb_north.inst.cb_conf_bus[47] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10030_ (.D(_03375_),
    .Q(\cb_north.inst.cb_conf_bus[48] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10031_ (.D(_03377_),
    .Q(\cb_north.inst.cb_conf_bus[49] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10032_ (.D(_03379_),
    .Q(\cb_north.inst.cb_conf_bus[50] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10033_ (.D(_03381_),
    .Q(\cb_north.inst.cb_conf_bus[51] ),
    .CLK(clknet_7_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10034_ (.D(_03383_),
    .Q(\cb_north.inst.cb_conf_bus[52] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10035_ (.D(_03385_),
    .Q(\cb_north.inst.cb_conf_bus[53] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10036_ (.D(_03387_),
    .Q(\cb_north.inst.cb_conf_bus[54] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10037_ (.D(_03389_),
    .Q(\cb_north.inst.cb_conf_bus[55] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10038_ (.D(_03391_),
    .Q(\cb_north.inst.cb_conf_bus[56] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10039_ (.D(_03393_),
    .Q(\cb_north.inst.cb_conf_bus[57] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10040_ (.D(_03395_),
    .Q(\cb_north.inst.cb_conf_bus[58] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10041_ (.D(_03397_),
    .Q(\cb_north.inst.cb_conf_bus[59] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10042_ (.D(_03399_),
    .Q(\cb_north.inst.cb_conf_bus[60] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10043_ (.D(_03401_),
    .Q(\cb_north.inst.cb_conf_bus[61] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10044_ (.D(_03403_),
    .Q(\cb_north.inst.cb_conf_bus[62] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10045_ (.D(_03405_),
    .Q(\cb_north.inst.cb_conf_bus[63] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10046_ (.D(_03407_),
    .Q(\cb_north.inst.cb_conf_bus[64] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10047_ (.D(_03409_),
    .Q(\cb_north.inst.cb_conf_bus[65] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10048_ (.D(_03411_),
    .Q(\cb_north.inst.cb_conf_bus[66] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10049_ (.D(_03413_),
    .Q(\cb_north.inst.cb_conf_bus[67] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10050_ (.D(_03415_),
    .Q(\cb_north.inst.cb_conf_bus[68] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10051_ (.D(_03417_),
    .Q(\cb_north.inst.cb_conf_bus[69] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10052_ (.D(_03419_),
    .Q(\cb_north.inst.cb_conf_bus[70] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10053_ (.D(_03421_),
    .Q(\cb_north.inst.cb_conf_bus[71] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10054_ (.D(_03423_),
    .Q(\cb_north.inst.cb_conf_bus[72] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10055_ (.D(_03425_),
    .Q(\cb_north.inst.cb_conf_bus[73] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10056_ (.D(_03427_),
    .Q(\cb_north.inst.cb_conf_bus[74] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10057_ (.D(_03429_),
    .Q(\cb_north.inst.cb_conf_bus[75] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10058_ (.D(_03431_),
    .Q(\cb_north.inst.cb_conf_bus[76] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10059_ (.D(_03433_),
    .Q(\cb_north.inst.cb_conf_bus[77] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10060_ (.D(_03435_),
    .Q(\cb_north.inst.cb_conf_bus[78] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10061_ (.D(_03437_),
    .Q(\cb_north.inst.cb_conf_bus[79] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10062_ (.D(_03439_),
    .Q(\cb_north.inst.cb_conf_bus[80] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10063_ (.D(_03441_),
    .Q(\cb_north.inst.cb_conf_bus[81] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10064_ (.D(_03443_),
    .Q(\cb_north.inst.cb_conf_bus[82] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10065_ (.D(_03445_),
    .Q(\cb_north.inst.cb_conf_bus[83] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10066_ (.D(_03447_),
    .Q(\cb_north.inst.cb_conf_bus[84] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10067_ (.D(_03449_),
    .Q(\cb_north.inst.cb_conf_bus[85] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10068_ (.D(_03451_),
    .Q(\cb_north.inst.cb_conf_bus[86] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10069_ (.D(_03453_),
    .Q(\cb_north.inst.cb_conf_bus[87] ),
    .CLK(clknet_7_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10070_ (.D(_03455_),
    .Q(\cb_north.inst.cb_conf_bus[88] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10071_ (.D(_03457_),
    .Q(\cb_north.inst.cb_conf_bus[89] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10072_ (.D(_03459_),
    .Q(\cb_north.inst.cb_conf_bus[90] ),
    .CLK(clknet_7_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10073_ (.D(_03461_),
    .Q(\cb_north.inst.cb_conf_bus[91] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10074_ (.D(_03463_),
    .Q(\cb_north.inst.cb_conf_bus[92] ),
    .CLK(clknet_7_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10075_ (.D(_03465_),
    .Q(\cb_north.inst.cb_conf_bus[93] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10076_ (.D(_03467_),
    .Q(\cb_north.inst.cb_conf_bus[94] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10077_ (.D(_03469_),
    .Q(\cb_north.inst.cb_conf_bus[95] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10078_ (.D(_03471_),
    .Q(\cb_north.inst.cb_conf_bus[96] ),
    .CLK(clknet_7_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10079_ (.D(_03473_),
    .Q(\cb_north.inst.cb_conf_bus[97] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10080_ (.D(_03475_),
    .Q(\cb_north.inst.cb_conf_bus[98] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10081_ (.D(_03477_),
    .Q(\cb_north.inst.cb_conf_bus[99] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10082_ (.D(_03479_),
    .Q(\cb_north.inst.cb_conf_bus[100] ),
    .CLK(clknet_7_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10083_ (.D(_03481_),
    .Q(\cb_north.inst.cb_conf_bus[101] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10084_ (.D(_03483_),
    .Q(\cb_north.inst.cb_conf_bus[102] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10085_ (.D(_03485_),
    .Q(\cb_north.inst.cb_conf_bus[103] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10086_ (.D(_03487_),
    .Q(\cb_north.inst.cb_conf_bus[104] ),
    .CLK(clknet_7_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10087_ (.D(_03489_),
    .Q(\cb_north.inst.cb_conf_bus[105] ),
    .CLK(clknet_7_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10088_ (.D(_03491_),
    .Q(\cb_north.inst.cb_conf_bus[106] ),
    .CLK(clknet_7_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10089_ (.D(_03493_),
    .Q(\cb_north.inst.cb_conf_bus[107] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10090_ (.D(_03495_),
    .Q(\cb_north.inst.cb_conf_bus[108] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10091_ (.D(_03497_),
    .Q(\cb_north.inst.cb_conf_bus[109] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10092_ (.D(_03499_),
    .Q(\cb_north.inst.cb_conf_bus[110] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10093_ (.D(_03501_),
    .Q(\cb_north.inst.cb_conf_bus[111] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10094_ (.D(_03503_),
    .Q(\cb_north.inst.cb_conf_bus[112] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10095_ (.D(_03505_),
    .Q(\cb_north.inst.cb_conf_bus[113] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10096_ (.D(_03507_),
    .Q(\cb_north.inst.cb_conf_bus[114] ),
    .CLK(clknet_7_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10097_ (.D(_03509_),
    .Q(\cb_north.inst.cb_conf_bus[115] ),
    .CLK(clknet_7_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10098_ (.D(_03511_),
    .Q(\cb_north.inst.cb_conf_bus[116] ),
    .CLK(clknet_7_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10099_ (.D(_03513_),
    .Q(\cb_north.inst.cb_conf_bus[117] ),
    .CLK(clknet_7_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10100_ (.D(_03515_),
    .Q(\cb_north.inst.cb_conf_bus[118] ),
    .CLK(clknet_7_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10101_ (.D(_03517_),
    .Q(\cb_north.inst.cb_conf_bus[119] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10102_ (.D(_03519_),
    .Q(\cb_north.inst.cb_conf_bus[120] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10103_ (.D(_03521_),
    .Q(\cb_north.inst.cb_conf_bus[121] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10104_ (.D(_03523_),
    .Q(\cb_north.inst.cb_conf_bus[122] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10105_ (.D(_03525_),
    .Q(\cb_north.inst.cb_conf_bus[123] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10106_ (.D(_03527_),
    .Q(\cb_north.inst.cb_conf_bus[124] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10107_ (.D(_03529_),
    .Q(\cb_north.inst.cb_conf_bus[125] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10108_ (.D(_03531_),
    .Q(\cb_north.inst.cb_conf_bus[126] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10109_ (.D(_03533_),
    .Q(\cb_north.inst.cb_conf_bus[127] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10110_ (.D(_03535_),
    .Q(\cb_north.inst.cb_conf_bus[128] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10111_ (.D(_03537_),
    .Q(\cb_north.inst.cb_conf_bus[129] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10112_ (.D(_03539_),
    .Q(\cb_north.inst.cb_conf_bus[130] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10113_ (.D(_03541_),
    .Q(\cb_north.inst.cb_conf_bus[131] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10114_ (.D(_03543_),
    .Q(\cb_north.inst.cb_conf_bus[132] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10115_ (.D(_03545_),
    .Q(\cb_north.inst.cb_conf_bus[133] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10116_ (.D(_03547_),
    .Q(\cb_north.inst.cb_conf_bus[134] ),
    .CLK(clknet_7_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10117_ (.D(_03549_),
    .Q(\cb_north.inst.cb_conf_bus[135] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10118_ (.D(_03551_),
    .Q(\cb_north.inst.cb_conf_bus[136] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10119_ (.D(_03553_),
    .Q(\cb_north.inst.cb_conf_bus[137] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10120_ (.D(_03555_),
    .Q(\cb_north.inst.cb_conf_bus[138] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10121_ (.D(_03557_),
    .Q(\cb_north.inst.cb_conf_bus[139] ),
    .CLK(clknet_7_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10122_ (.D(_03559_),
    .Q(\cb_north.inst.cb_conf_bus[140] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10123_ (.D(_03561_),
    .Q(\cb_north.inst.cb_conf_bus[141] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10124_ (.D(_03563_),
    .Q(\cb_north.inst.cb_conf_bus[142] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10125_ (.D(_03565_),
    .Q(\cb_north.inst.cb_conf_bus[143] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10126_ (.D(_03567_),
    .Q(\cb_north.inst.cb_conf_bus[144] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10127_ (.D(_03569_),
    .Q(\cb_north.inst.cb_conf_bus[145] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10128_ (.D(_03571_),
    .Q(\cb_north.inst.cb_conf_bus[146] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10129_ (.D(_03573_),
    .Q(\cb_north.inst.cb_conf_bus[147] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10130_ (.D(_03575_),
    .Q(\cb_north.inst.cb_conf_bus[148] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10131_ (.D(_03577_),
    .Q(\cb_north.inst.cb_conf_bus[149] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10132_ (.D(_03579_),
    .Q(\cb_north.inst.cb_conf_bus[150] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10133_ (.D(_03581_),
    .Q(\cb_north.inst.cb_conf_bus[151] ),
    .CLK(clknet_7_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10134_ (.D(_03583_),
    .Q(\cb_north.inst.cb_conf_bus[152] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10135_ (.D(_03585_),
    .Q(\cb_north.inst.cb_conf_bus[153] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10136_ (.D(_03587_),
    .Q(\cb_north.inst.cb_conf_bus[154] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10137_ (.D(_03589_),
    .Q(\cb_north.inst.cb_conf_bus[155] ),
    .CLK(clknet_7_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10138_ (.D(_03591_),
    .Q(\cb_north.inst.cb_conf_bus[156] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10139_ (.D(_03593_),
    .Q(\cb_north.inst.cb_conf_bus[157] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10140_ (.D(_03595_),
    .Q(\cb_north.inst.cb_conf_bus[158] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10141_ (.D(_03597_),
    .Q(\cb_north.inst.cb_conf_bus[159] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10142_ (.D(_03599_),
    .Q(\cb_north.inst.cb_conf_bus[160] ),
    .CLK(clknet_7_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10143_ (.D(_03601_),
    .Q(\cb_north.inst.cb_conf_bus[161] ),
    .CLK(clknet_7_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10144_ (.D(_03603_),
    .Q(\cb_north.inst.cb_conf_bus[162] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10145_ (.D(_03605_),
    .Q(\cb_north.inst.cb_conf_bus[163] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10146_ (.D(_03607_),
    .Q(\cb_north.inst.cb_conf_bus[164] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10147_ (.D(_03609_),
    .Q(\cb_north.inst.cb_conf_bus[165] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10148_ (.D(_03611_),
    .Q(\cb_north.inst.cb_conf_bus[166] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10149_ (.D(_03613_),
    .Q(\cb_north.inst.cb_conf_bus[167] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10150_ (.D(_03615_),
    .Q(\cb_north.inst.cb_conf_bus[168] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10151_ (.D(_03617_),
    .Q(\cb_north.inst.cb_conf_bus[169] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10152_ (.D(_03619_),
    .Q(\cb_north.inst.cb_conf_bus[170] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10153_ (.D(_03621_),
    .Q(\cb_north.inst.cb_conf_bus[171] ),
    .CLK(clknet_7_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10154_ (.D(_03623_),
    .Q(\cb_north.inst.cb_conf_bus[172] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10155_ (.D(_03625_),
    .Q(\cb_north.inst.cb_conf_bus[173] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10156_ (.D(_03627_),
    .Q(\cb_north.inst.cb_conf_bus[174] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10157_ (.D(_03629_),
    .Q(\cb_north.inst.cb_conf_bus[175] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10158_ (.D(_03631_),
    .Q(\cb_north.inst.cb_conf_bus[176] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10159_ (.D(_03633_),
    .Q(\cb_north.inst.cb_conf_bus[177] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10160_ (.D(_03635_),
    .Q(\cb_north.inst.cb_conf_bus[178] ),
    .CLK(clknet_7_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10161_ (.D(_03637_),
    .Q(\cb_north.inst.cb_conf_bus[179] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10162_ (.D(_03639_),
    .Q(\cb_north.inst.cb_conf_bus[180] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10163_ (.D(_03641_),
    .Q(\cb_north.inst.cb_conf_bus[181] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10164_ (.D(_03643_),
    .Q(\cb_north.inst.cb_conf_bus[182] ),
    .CLK(clknet_7_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10165_ (.D(_03645_),
    .Q(\cb_north.inst.cb_conf_bus[183] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10166_ (.D(_03647_),
    .Q(\cb_north.inst.cb_conf_bus[184] ),
    .CLK(clknet_7_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10167_ (.D(_03649_),
    .Q(\cb_north.inst.cb_conf_bus[185] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10168_ (.D(_03651_),
    .Q(\cb_north.inst.cb_conf_bus[186] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10169_ (.D(_03653_),
    .Q(\cb_north.inst.cb_conf_bus[187] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10170_ (.D(_03655_),
    .Q(\cb_north.inst.cb_conf_bus[188] ),
    .CLK(clknet_7_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10171_ (.D(_03657_),
    .Q(\cb_north.inst.cb_conf_bus[189] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10172_ (.D(_03659_),
    .Q(\cb_north.inst.cb_conf_bus[190] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10173_ (.D(_03661_),
    .Q(\cb_north.inst.cb_conf_bus[191] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10174_ (.D(_03663_),
    .Q(\cb_north.inst.cb_conf_bus[192] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10175_ (.D(_03665_),
    .Q(\cb_north.inst.cb_conf_bus[193] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10176_ (.D(_03667_),
    .Q(\cb_north.inst.cb_conf_bus[194] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10177_ (.D(_03669_),
    .Q(\cb_north.inst.cb_conf_bus[195] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10178_ (.D(_03671_),
    .Q(\cb_north.inst.cb_conf_bus[196] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10179_ (.D(_03673_),
    .Q(\cb_north.inst.cb_conf_bus[197] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10180_ (.D(_03675_),
    .Q(\cb_north.inst.cb_conf_bus[198] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10181_ (.D(_03677_),
    .Q(\cb_north.inst.cb_conf_bus[199] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10182_ (.D(_03679_),
    .Q(\cb_north.inst.cb_conf_bus[200] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10183_ (.D(_03681_),
    .Q(\cb_north.inst.cb_conf_bus[201] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10184_ (.D(_03683_),
    .Q(\cb_north.inst.cb_conf_bus[202] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10185_ (.D(_03685_),
    .Q(\cb_north.inst.cb_conf_bus[203] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10186_ (.D(_03687_),
    .Q(\cb_north.inst.cb_conf_bus[204] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10187_ (.D(_03689_),
    .Q(\cb_north.inst.cb_conf_bus[205] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10188_ (.D(_03691_),
    .Q(\cb_north.inst.cb_conf_bus[206] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10189_ (.D(_03693_),
    .Q(\cb_north.inst.cb_conf_bus[207] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10190_ (.D(_03695_),
    .Q(\cb_north.inst.cb_conf_bus[208] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10191_ (.D(_03697_),
    .Q(\cb_north.inst.cb_conf_bus[209] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10192_ (.D(_03699_),
    .Q(\cb_north.inst.cb_conf_bus[210] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10193_ (.D(_03701_),
    .Q(\cb_north.inst.cb_conf_bus[211] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10194_ (.D(_03703_),
    .Q(\cb_north.inst.cb_conf_bus[212] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10195_ (.D(_03705_),
    .Q(\cb_north.inst.cb_conf_bus[213] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10196_ (.D(_03707_),
    .Q(\cb_north.inst.cb_conf_bus[214] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10197_ (.D(_03709_),
    .Q(\cb_north.inst.cb_conf_bus[215] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10198_ (.D(_03711_),
    .Q(\cb_north.inst.cb_conf_bus[216] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10199_ (.D(_03713_),
    .Q(\cb_north.inst.cb_conf_bus[217] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10200_ (.D(_03715_),
    .Q(\cb_north.inst.cb_conf_bus[218] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10201_ (.D(_03717_),
    .Q(\cb_north.inst.cb_conf_bus[219] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10202_ (.D(_03719_),
    .Q(\cb_north.inst.cb_conf_bus[220] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10203_ (.D(_03721_),
    .Q(\cb_north.inst.cb_conf_bus[221] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10204_ (.D(_03723_),
    .Q(\cb_north.inst.cb_conf_bus[222] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10205_ (.D(_03725_),
    .Q(\cb_north.inst.cb_conf_bus[223] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10206_ (.D(_03727_),
    .Q(\cb_north.inst.cb_conf_bus[224] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10207_ (.D(_03729_),
    .Q(\cb_north.inst.cb_conf_bus[225] ),
    .CLK(clknet_7_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10208_ (.D(_03731_),
    .Q(\cb_north.inst.cb_conf_bus[226] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10209_ (.D(_03733_),
    .Q(\cb_north.inst.cb_conf_bus[227] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10210_ (.D(_03735_),
    .Q(\cb_north.inst.cb_conf_bus[228] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10211_ (.D(_03737_),
    .Q(\cb_north.inst.cb_conf_bus[229] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10212_ (.D(_03739_),
    .Q(\cb_north.inst.cb_conf_bus[230] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10213_ (.D(_03741_),
    .Q(\cb_north.inst.cb_conf_bus[231] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10214_ (.D(_03743_),
    .Q(\cb_north.inst.cb_conf_bus[232] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10215_ (.D(_03745_),
    .Q(\cb_north.inst.cb_conf_bus[233] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10216_ (.D(_03747_),
    .Q(\cb_north.inst.cb_conf_bus[234] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10217_ (.D(_03749_),
    .Q(\cb_north.inst.cb_conf_bus[235] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10218_ (.D(_03751_),
    .Q(\cb_north.inst.cb_conf_bus[236] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10219_ (.D(_03753_),
    .Q(\cb_north.inst.cb_conf_bus[237] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10220_ (.D(_03755_),
    .Q(\cb_north.inst.cb_conf_bus[238] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10221_ (.D(_03757_),
    .Q(\cb_north.inst.cb_conf_bus[239] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10222_ (.D(_03759_),
    .Q(\cb_north.inst.cb_conf_bus[240] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10223_ (.D(_03761_),
    .Q(\cb_north.inst.cb_conf_bus[241] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10224_ (.D(_03763_),
    .Q(\cb_north.inst.cb_conf_bus[242] ),
    .CLK(clknet_7_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10225_ (.D(_03765_),
    .Q(\cb_north.inst.cb_conf_bus[243] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10226_ (.D(_03767_),
    .Q(\cb_north.inst.cb_conf_bus[244] ),
    .CLK(clknet_7_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10227_ (.D(_03769_),
    .Q(\cb_north.inst.cb_conf_bus[245] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10228_ (.D(_03771_),
    .Q(\cb_north.inst.cb_conf_bus[246] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10229_ (.D(_03773_),
    .Q(\cb_north.inst.cb_conf_bus[247] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10230_ (.D(_03775_),
    .Q(\cb_north.inst.cb_conf_bus[248] ),
    .CLK(clknet_7_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10231_ (.D(_03777_),
    .Q(\cb_north.inst.cb_conf_bus[249] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10232_ (.D(_03779_),
    .Q(\cb_north.inst.cb_conf_bus[250] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10233_ (.D(_03781_),
    .Q(\cb_north.inst.cb_conf_bus[251] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10234_ (.D(_03783_),
    .Q(\cb_north.inst.cb_conf_bus[252] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10235_ (.D(_03785_),
    .Q(\cb_north.inst.cb_conf_bus[253] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10236_ (.D(_03787_),
    .Q(\cb_north.inst.cb_conf_bus[254] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10237_ (.D(_03789_),
    .Q(\cb_north.inst.cb_conf_bus[255] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10238_ (.D(_03791_),
    .Q(\cb_north.inst.cb_conf_bus[256] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10239_ (.D(_03793_),
    .Q(\cb_north.inst.cb_conf_bus[257] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10240_ (.D(_03795_),
    .Q(\cb_north.inst.cb_conf_bus[258] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10241_ (.D(_03797_),
    .Q(\cb_north.inst.cb_conf_bus[259] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10242_ (.D(_03799_),
    .Q(\cb_north.inst.cb_conf_bus[260] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10243_ (.D(_03801_),
    .Q(\cb_north.inst.cb_conf_bus[261] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10244_ (.D(_03803_),
    .Q(\cb_north.inst.cb_conf_bus[262] ),
    .CLK(clknet_7_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10245_ (.D(_03805_),
    .Q(\cb_north.inst.cb_conf_bus[263] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10246_ (.D(_03807_),
    .Q(\cb_north.inst.cb_conf_bus[264] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10247_ (.D(_03809_),
    .Q(\cb_north.inst.cb_conf_bus[265] ),
    .CLK(clknet_7_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10248_ (.D(_03811_),
    .Q(\cb_north.inst.cb_conf_bus[266] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10249_ (.D(_03813_),
    .Q(\cb_north.inst.cb_conf_bus[267] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10250_ (.D(_03815_),
    .Q(\cb_north.inst.cb_conf_bus[268] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10251_ (.D(_03817_),
    .Q(\cb_north.inst.cb_conf_bus[269] ),
    .CLK(clknet_7_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10252_ (.D(_03819_),
    .Q(\cb_north.inst.cb_conf_bus[270] ),
    .CLK(clknet_7_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10253_ (.D(_03821_),
    .Q(\cb_north.inst.cb_conf_bus[271] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10254_ (.D(_03823_),
    .Q(\cb_north.inst.cb_conf_bus[272] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10255_ (.D(_03825_),
    .Q(\cb_north.inst.cb_conf_bus[273] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10256_ (.D(_03827_),
    .Q(\cb_north.inst.cb_conf_bus[274] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10257_ (.D(_03829_),
    .Q(\cb_north.inst.cb_conf_bus[275] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10258_ (.D(_03831_),
    .Q(\cb_north.inst.cb_conf_bus[276] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10259_ (.D(_03833_),
    .Q(\cb_north.inst.cb_conf_bus[277] ),
    .CLK(clknet_7_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10260_ (.D(_03835_),
    .Q(\cb_north.inst.cb_conf_bus[278] ),
    .CLK(clknet_7_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10261_ (.D(_03837_),
    .Q(\cb_north.inst.cb_conf_bus[279] ),
    .CLK(clknet_7_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10262_ (.D(_03839_),
    .Q(\cb_north.inst.cb_conf_bus[280] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10263_ (.D(_03841_),
    .Q(\cb_north.inst.cb_conf_bus[281] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10264_ (.D(_03843_),
    .Q(\cb_north.inst.cb_conf_bus[282] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10265_ (.D(_03845_),
    .Q(\cb_north.inst.cb_conf_bus[283] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10266_ (.D(_03847_),
    .Q(\cb_north.inst.cb_conf_bus[284] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10267_ (.D(_03849_),
    .Q(\cb_north.inst.cb_conf_bus[285] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10268_ (.D(_03851_),
    .Q(\cb_north.inst.cb_conf_bus[286] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10269_ (.D(_03853_),
    .Q(\cb_north.inst.cb_conf_bus[287] ),
    .CLK(clknet_7_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10270_ (.D(_03855_),
    .Q(\cb_north.inst.cb_conf_bus[288] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10271_ (.D(_03857_),
    .Q(\cb_north.inst.cb_conf_bus[289] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10272_ (.D(_03859_),
    .Q(\cb_north.inst.cb_conf_bus[290] ),
    .CLK(clknet_7_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10273_ (.D(_03861_),
    .Q(\cb_north.inst.cb_conf_bus[291] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10274_ (.D(_03863_),
    .Q(\cb_north.inst.cb_conf_bus[292] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10275_ (.D(_03865_),
    .Q(\cb_north.inst.cb_conf_bus[293] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10276_ (.D(_03867_),
    .Q(\cb_north.inst.cb_conf_bus[294] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10277_ (.D(_03869_),
    .Q(\cb_north.inst.cb_conf_bus[295] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10278_ (.D(_03871_),
    .Q(\cb_north.inst.cb_conf_bus[296] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10279_ (.D(_03873_),
    .Q(\cb_north.inst.cb_conf_bus[297] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10280_ (.D(_03875_),
    .Q(\cb_north.inst.cb_conf_bus[298] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10281_ (.D(_03877_),
    .Q(\cb_north.inst.cb_conf_bus[299] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10282_ (.D(_03879_),
    .Q(\cb_north.inst.cb_conf_bus[300] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10283_ (.D(_03881_),
    .Q(\cb_north.inst.cb_conf_bus[301] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10284_ (.D(_03883_),
    .Q(\cb_north.inst.cb_conf_bus[302] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10285_ (.D(_03885_),
    .Q(\cb_north.inst.cb_conf_bus[303] ),
    .CLK(clknet_7_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10286_ (.D(_03887_),
    .Q(\cb_north.inst.cb_conf_bus[304] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10287_ (.D(_03889_),
    .Q(\cb_north.inst.cb_conf_bus[305] ),
    .CLK(clknet_7_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10288_ (.D(_03891_),
    .Q(\cb_north.inst.cb_conf_bus[306] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10289_ (.D(_03893_),
    .Q(\cb_north.inst.cb_conf_bus[307] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10290_ (.D(_03895_),
    .Q(\cb_north.inst.cb_conf_bus[308] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10291_ (.D(_03897_),
    .Q(\cb_north.inst.cb_conf_bus[309] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10292_ (.D(_03899_),
    .Q(\cb_north.inst.cb_conf_bus[310] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10293_ (.D(_03901_),
    .Q(\cb_north.inst.cb_conf_bus[311] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10294_ (.D(_03903_),
    .Q(\cb_north.inst.cb_conf_bus[312] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10295_ (.D(_03905_),
    .Q(\cb_north.inst.cb_conf_bus[313] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10296_ (.D(_03907_),
    .Q(\cb_north.inst.cb_conf_bus[314] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10297_ (.D(_03909_),
    .Q(\cb_north.inst.cb_conf_bus[315] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10298_ (.D(_03911_),
    .Q(\cb_north.inst.cb_conf_bus[316] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10299_ (.D(_03913_),
    .Q(\cb_north.inst.cb_conf_bus[317] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10300_ (.D(_03915_),
    .Q(\cb_north.inst.cb_conf_bus[318] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10301_ (.D(_03917_),
    .Q(\cb_north.inst.cb_conf_bus[319] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10302_ (.D(_03919_),
    .Q(\cb_north.inst.cb_conf_bus[320] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10303_ (.D(_03921_),
    .Q(\cb_north.inst.cb_conf_bus[321] ),
    .CLK(clknet_7_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10304_ (.D(_03923_),
    .Q(\cb_north.inst.cb_conf_bus[322] ),
    .CLK(clknet_7_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10305_ (.D(_03925_),
    .Q(\cb_north.inst.cb_conf_bus[323] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10306_ (.D(_03927_),
    .Q(\cb_north.inst.cb_conf_bus[324] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10307_ (.D(_03929_),
    .Q(\cb_north.inst.cb_conf_bus[325] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10308_ (.D(_03931_),
    .Q(\cb_north.inst.cb_conf_bus[326] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10309_ (.D(_03933_),
    .Q(\cb_north.inst.cb_conf_bus[327] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10310_ (.D(_03935_),
    .Q(\cb_north.inst.cb_conf_bus[328] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10311_ (.D(_03937_),
    .Q(\cb_north.inst.cb_conf_bus[329] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10312_ (.D(_03939_),
    .Q(\cb_north.inst.cb_conf_bus[330] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10313_ (.D(_03941_),
    .Q(\cb_north.inst.cb_conf_bus[331] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10314_ (.D(_03943_),
    .Q(\cb_north.inst.cb_conf_bus[332] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10315_ (.D(_03945_),
    .Q(\cb_north.inst.cb_conf_bus[333] ),
    .CLK(clknet_7_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10316_ (.D(_03947_),
    .Q(\cb_north.inst.cb_conf_bus[334] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10317_ (.D(_03949_),
    .Q(\cb_north.inst.cb_conf_bus[335] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10318_ (.D(_03951_),
    .Q(\cb_north.inst.cb_conf_bus[336] ),
    .CLK(clknet_7_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10319_ (.D(_03953_),
    .Q(\cb_north.inst.cb_conf_bus[337] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10320_ (.D(_03955_),
    .Q(\cb_north.inst.cb_conf_bus[338] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10321_ (.D(_03957_),
    .Q(\cb_north.inst.cb_conf_bus[339] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10322_ (.D(_03959_),
    .Q(\cb_north.inst.cb_conf_bus[340] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10323_ (.D(_03961_),
    .Q(\cb_north.inst.cb_conf_bus[341] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10324_ (.D(_03963_),
    .Q(\cb_north.inst.cb_conf_bus[342] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10325_ (.D(_03965_),
    .Q(\cb_north.inst.cb_conf_bus[343] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10326_ (.D(_03967_),
    .Q(\cb_north.inst.cb_conf_bus[344] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10327_ (.D(_03969_),
    .Q(\cb_north.inst.cb_conf_bus[345] ),
    .CLK(clknet_7_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10328_ (.D(_03971_),
    .Q(\cb_north.inst.cb_conf_bus[346] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10329_ (.D(_03973_),
    .Q(\cb_north.inst.cb_conf_bus[347] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10330_ (.D(_03975_),
    .Q(\cb_north.inst.cb_conf_bus[348] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10331_ (.D(_03977_),
    .Q(\cb_north.inst.cb_conf_bus[349] ),
    .CLK(clknet_7_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10332_ (.D(_03979_),
    .Q(\cb_north.inst.cb_conf_bus[350] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10333_ (.D(_03981_),
    .Q(\cb_north.inst.cb_conf_bus[351] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10334_ (.D(_03983_),
    .Q(\cb_north.inst.cb_conf_bus[352] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10335_ (.D(_03985_),
    .Q(\cb_north.inst.cb_conf_bus[353] ),
    .CLK(clknet_7_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10336_ (.D(_03987_),
    .Q(\cb_north.inst.cb_conf_bus[354] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10337_ (.D(_03989_),
    .Q(\cb_north.inst.cb_conf_bus[355] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10338_ (.D(_03991_),
    .Q(\cb_north.inst.cb_conf_bus[356] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10339_ (.D(_03993_),
    .Q(\cb_north.inst.cb_conf_bus[357] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10340_ (.D(_03995_),
    .Q(\cb_north.inst.cb_conf_bus[358] ),
    .CLK(clknet_7_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10341_ (.D(_03997_),
    .Q(\cb_north.inst.cb_conf_bus[359] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10342_ (.D(_03999_),
    .Q(\cb_north.inst.cb_conf_bus[360] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10343_ (.D(_04001_),
    .Q(\cb_north.inst.cb_conf_bus[361] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10344_ (.D(_04003_),
    .Q(\cb_north.inst.cb_conf_bus[362] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10345_ (.D(_04005_),
    .Q(\cb_north.inst.cb_conf_bus[363] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10346_ (.D(_04007_),
    .Q(\cb_north.inst.cb_conf_bus[364] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10347_ (.D(_04009_),
    .Q(\cb_north.inst.cb_conf_bus[365] ),
    .CLK(clknet_7_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10348_ (.D(_04011_),
    .Q(\cb_north.inst.cb_conf_bus[366] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10349_ (.D(_04013_),
    .Q(\cb_north.inst.cb_conf_bus[367] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10350_ (.D(_04015_),
    .Q(\cb_north.inst.cb_conf_bus[368] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10351_ (.D(_04017_),
    .Q(\cb_north.inst.cb_conf_bus[369] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10352_ (.D(_04019_),
    .Q(\cb_north.inst.cb_conf_bus[370] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10353_ (.D(_04021_),
    .Q(\cb_north.inst.cb_conf_bus[371] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10354_ (.D(_04023_),
    .Q(\cb_north.inst.cb_conf_bus[372] ),
    .CLK(clknet_7_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10355_ (.D(_04025_),
    .Q(\cb_north.inst.cb_conf_bus[373] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10356_ (.D(_04027_),
    .Q(\cb_north.inst.cb_conf_bus[374] ),
    .CLK(clknet_7_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10357_ (.D(_04029_),
    .Q(\cb_north.inst.cb_conf_bus[375] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10358_ (.D(_04031_),
    .Q(\cb_north.inst.cb_conf_bus[376] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10359_ (.D(_04033_),
    .Q(\cb_north.inst.cb_conf_bus[377] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10360_ (.D(_04035_),
    .Q(\cb_north.inst.cb_conf_bus[378] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10361_ (.D(_04037_),
    .Q(\cb_north.inst.cb_conf_bus[379] ),
    .CLK(clknet_7_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10362_ (.D(_04039_),
    .Q(\cb_north.inst.cb_conf_bus[380] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10363_ (.D(_04041_),
    .Q(\cb_north.inst.cb_conf_bus[381] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10364_ (.D(_04043_),
    .Q(\cb_north.inst.cb_conf_bus[382] ),
    .CLK(clknet_7_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10365_ (.D(_04045_),
    .Q(\cb_north.inst.cb_conf_bus[383] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10366_ (.D(_04047_),
    .Q(\cb_north.inst.cb_conf_bus[384] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10367_ (.D(_04049_),
    .Q(\cb_north.inst.cb_conf_bus[385] ),
    .CLK(clknet_7_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10368_ (.D(_04051_),
    .Q(\cb_north.inst.cb_conf_bus[386] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10369_ (.D(_04053_),
    .Q(\cb_north.inst.cb_conf_bus[387] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10370_ (.D(_04055_),
    .Q(\cb_north.inst.cb_conf_bus[388] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10371_ (.D(_04057_),
    .Q(\cb_north.inst.cb_conf_bus[389] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10372_ (.D(_04059_),
    .Q(\cb_north.inst.cb_conf_bus[390] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10373_ (.D(_04061_),
    .Q(\cb_north.inst.cb_conf_bus[391] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10374_ (.D(_04063_),
    .Q(\cb_north.inst.cb_conf_bus[392] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10375_ (.D(_04065_),
    .Q(\cb_north.inst.cb_conf_bus[393] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10376_ (.D(_04067_),
    .Q(\cb_north.inst.cb_conf_bus[394] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10377_ (.D(_04069_),
    .Q(\cb_north.inst.cb_conf_bus[395] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10378_ (.D(_04071_),
    .Q(\cb_north.inst.cb_conf_bus[396] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10379_ (.D(_04073_),
    .Q(\cb_north.inst.cb_conf_bus[397] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10380_ (.D(_04075_),
    .Q(\cb_north.inst.cb_conf_bus[398] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10381_ (.D(_04077_),
    .Q(\cb_north.inst.cb_conf_bus[399] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10382_ (.D(_04079_),
    .Q(\cb_north.inst.cb_conf_bus[400] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10383_ (.D(_04081_),
    .Q(\cb_north.inst.cb_conf_bus[401] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10384_ (.D(_04083_),
    .Q(\cb_north.inst.cb_conf_bus[402] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10385_ (.D(_04085_),
    .Q(\cb_north.inst.cb_conf_bus[403] ),
    .CLK(clknet_7_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10386_ (.D(_04087_),
    .Q(\cb_north.inst.cb_conf_bus[404] ),
    .CLK(clknet_7_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10387_ (.D(_04089_),
    .Q(\cb_north.inst.cb_conf_bus[405] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10388_ (.D(_04091_),
    .Q(\cb_north.inst.cb_conf_bus[406] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10389_ (.D(_04093_),
    .Q(\cb_north.inst.cb_conf_bus[407] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10390_ (.D(_04095_),
    .Q(\cb_north.inst.cb_conf_bus[408] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10391_ (.D(_04097_),
    .Q(\cb_north.inst.cb_conf_bus[409] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10392_ (.D(_04099_),
    .Q(\cb_north.inst.cb_conf_bus[410] ),
    .CLK(clknet_7_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10393_ (.D(_04101_),
    .Q(\cb_north.inst.cb_conf_bus[411] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10394_ (.D(_04103_),
    .Q(\cb_north.inst.cb_conf_bus[412] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10395_ (.D(_04105_),
    .Q(\cb_north.inst.cb_conf_bus[413] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10396_ (.D(_04107_),
    .Q(\cb_north.inst.cb_conf_bus[414] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10397_ (.D(_04109_),
    .Q(\cb_north.inst.cb_conf_bus[415] ),
    .CLK(clknet_7_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10398_ (.D(_04111_),
    .Q(\cb_north.inst.cb_conf_bus[416] ),
    .CLK(clknet_7_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10399_ (.D(_04113_),
    .Q(\cb_north.inst.cb_conf_bus[417] ),
    .CLK(clknet_7_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10400_ (.D(_04115_),
    .Q(\cb_north.inst.cb_conf_bus[418] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10401_ (.D(_04117_),
    .Q(\cb_north.inst.cb_conf_bus[419] ),
    .CLK(clknet_7_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _10402_ (.D(_04119_),
    .Q(\cb_north.inst.configuroni.comb_shifter.config_data[420] ),
    .CLK(clknet_7_73_0_clk));
 sky130_fd_sc_hd__dlxtp_1 _10403_ (.D(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_in ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10404_ (.D(\sb.configuroni.comb_config[1] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10405_ (.D(\sb.configuroni.comb_config[2] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10406_ (.D(\sb.configuroni.comb_config[3] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10407_ (.D(\sb.configuroni.comb_config[4] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10408_ (.D(\sb.configuroni.comb_config[5] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10409_ (.D(\sb.configuroni.comb_config[6] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10410_ (.D(\sb.configuroni.comb_config[7] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10411_ (.D(\sb.configuroni.comb_config[8] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.n1e1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10412_ (.D(\sb.configuroni.comb_config[9] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.e0s1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10413_ (.D(\sb.configuroni.comb_config[10] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.s0w0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10414_ (.D(\sb.configuroni.comb_config[11] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[0].elem.w1n0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10415_ (.D(\sb.configuroni.comb_config[12] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10416_ (.D(\sb.configuroni.comb_config[13] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10417_ (.D(\sb.configuroni.comb_config[14] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10418_ (.D(\sb.configuroni.comb_config[15] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10419_ (.D(\sb.configuroni.comb_config[16] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10420_ (.D(\sb.configuroni.comb_config[17] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10421_ (.D(\sb.configuroni.comb_config[18] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10422_ (.D(\sb.configuroni.comb_config[19] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10423_ (.D(\sb.configuroni.comb_config[20] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.n1e1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10424_ (.D(\sb.configuroni.comb_config[21] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.e0s1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10425_ (.D(\sb.configuroni.comb_config[22] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.s0w0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10426_ (.D(\sb.configuroni.comb_config[23] ),
    .Q(\sb.switcharoni.susb.switch_box_element_two[1].elem.w1n0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10427_ (.D(\sb.configuroni.comb_config[24] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10428_ (.D(\sb.configuroni.comb_config[25] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10429_ (.D(\sb.configuroni.comb_config[26] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10430_ (.D(\sb.configuroni.comb_config[27] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10431_ (.D(\sb.configuroni.comb_config[28] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10432_ (.D(\sb.configuroni.comb_config[29] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10433_ (.D(\sb.configuroni.comb_config[30] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10434_ (.D(\sb.configuroni.comb_config[31] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10435_ (.D(\sb.configuroni.comb_config[32] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n1e1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10436_ (.D(\sb.configuroni.comb_config[33] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e0s1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10437_ (.D(\sb.configuroni.comb_config[34] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s0w0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10438_ (.D(\sb.configuroni.comb_config[35] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w1n0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10439_ (.D(\sb.configuroni.comb_config[36] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10440_ (.D(\sb.configuroni.comb_config[37] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10441_ (.D(\sb.configuroni.comb_config[38] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10442_ (.D(\sb.configuroni.comb_config[39] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10443_ (.D(\sb.configuroni.comb_config[40] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0s0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10444_ (.D(\sb.configuroni.comb_config[41] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1w1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10445_ (.D(\sb.configuroni.comb_config[42] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1n1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10446_ (.D(\sb.configuroni.comb_config[43] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0e0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10447_ (.D(\sb.configuroni.comb_config[44] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n1e1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10448_ (.D(\sb.configuroni.comb_config[45] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e0s1.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10449_ (.D(\sb.configuroni.comb_config[46] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s0w0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10450_ (.D(\sb.configuroni.comb_config[47] ),
    .Q(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w1n0.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10451_ (.D(\slice.configuroni.comb_config[0] ),
    .Q(_04152_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10452_ (.D(\slice.configuroni.comb_config[1] ),
    .Q(_04159_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10453_ (.D(\slice.configuroni.comb_config[2] ),
    .Q(_04160_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10454_ (.D(\slice.configuroni.comb_config[3] ),
    .Q(_04161_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10455_ (.D(\slice.configuroni.comb_config[4] ),
    .Q(_04162_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10456_ (.D(\slice.configuroni.comb_config[5] ),
    .Q(_04163_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10457_ (.D(\slice.configuroni.comb_config[6] ),
    .Q(_04164_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10458_ (.D(\slice.configuroni.comb_config[7] ),
    .Q(_04165_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10459_ (.D(\slice.configuroni.comb_config[8] ),
    .Q(_04166_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10460_ (.D(\slice.configuroni.comb_config[9] ),
    .Q(_04167_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10461_ (.D(\slice.configuroni.comb_config[10] ),
    .Q(_04153_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10462_ (.D(\slice.configuroni.comb_config[11] ),
    .Q(_04154_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10463_ (.D(\slice.configuroni.comb_config[12] ),
    .Q(_04155_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10464_ (.D(\slice.configuroni.comb_config[13] ),
    .Q(_04156_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10465_ (.D(\slice.configuroni.comb_config[14] ),
    .Q(_04157_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10466_ (.D(\slice.configuroni.comb_config[15] ),
    .Q(_04158_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10467_ (.D(\slice.configuroni.comb_config[16] ),
    .Q(_04128_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10468_ (.D(\slice.configuroni.comb_config[17] ),
    .Q(_04135_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10469_ (.D(\slice.configuroni.comb_config[18] ),
    .Q(_04136_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10470_ (.D(\slice.configuroni.comb_config[19] ),
    .Q(_04137_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10471_ (.D(\slice.configuroni.comb_config[20] ),
    .Q(_04138_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10472_ (.D(\slice.configuroni.comb_config[21] ),
    .Q(_04139_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10473_ (.D(\slice.configuroni.comb_config[22] ),
    .Q(_04140_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10474_ (.D(\slice.configuroni.comb_config[23] ),
    .Q(_04141_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10475_ (.D(\slice.configuroni.comb_config[24] ),
    .Q(_04142_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10476_ (.D(\slice.configuroni.comb_config[25] ),
    .Q(_04143_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10477_ (.D(\slice.configuroni.comb_config[26] ),
    .Q(_04129_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10478_ (.D(\slice.configuroni.comb_config[27] ),
    .Q(_04130_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10479_ (.D(\slice.configuroni.comb_config[28] ),
    .Q(_04131_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10480_ (.D(\slice.configuroni.comb_config[29] ),
    .Q(_04132_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10481_ (.D(\slice.configuroni.comb_config[30] ),
    .Q(_04133_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10482_ (.D(\slice.configuroni.comb_config[31] ),
    .Q(_04134_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10483_ (.D(\slice.configuroni.comb_config[33] ),
    .Q(_04201_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10484_ (.D(\slice.configuroni.comb_config[34] ),
    .Q(_04208_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10485_ (.D(\slice.configuroni.comb_config[35] ),
    .Q(_04209_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10486_ (.D(\slice.configuroni.comb_config[36] ),
    .Q(_04210_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10487_ (.D(\slice.configuroni.comb_config[37] ),
    .Q(_04211_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10488_ (.D(\slice.configuroni.comb_config[38] ),
    .Q(_04212_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10489_ (.D(\slice.configuroni.comb_config[39] ),
    .Q(_04213_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10490_ (.D(\slice.configuroni.comb_config[40] ),
    .Q(_04214_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10491_ (.D(\slice.configuroni.comb_config[41] ),
    .Q(_04215_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10492_ (.D(\slice.configuroni.comb_config[42] ),
    .Q(_04216_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10493_ (.D(\slice.configuroni.comb_config[43] ),
    .Q(_04202_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10494_ (.D(\slice.configuroni.comb_config[44] ),
    .Q(_04203_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10495_ (.D(\slice.configuroni.comb_config[45] ),
    .Q(_04204_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10496_ (.D(\slice.configuroni.comb_config[46] ),
    .Q(_04205_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10497_ (.D(\slice.configuroni.comb_config[47] ),
    .Q(_04206_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10498_ (.D(\slice.configuroni.comb_config[48] ),
    .Q(_04207_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10499_ (.D(\slice.configuroni.comb_config[49] ),
    .Q(_04177_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10500_ (.D(\slice.configuroni.comb_config[50] ),
    .Q(_04184_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10501_ (.D(\slice.configuroni.comb_config[51] ),
    .Q(_04185_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10502_ (.D(\slice.configuroni.comb_config[52] ),
    .Q(_04186_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10503_ (.D(\slice.configuroni.comb_config[53] ),
    .Q(_04187_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10504_ (.D(\slice.configuroni.comb_config[54] ),
    .Q(_04188_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10505_ (.D(\slice.configuroni.comb_config[55] ),
    .Q(_04189_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10506_ (.D(\slice.configuroni.comb_config[56] ),
    .Q(_04190_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10507_ (.D(\slice.configuroni.comb_config[57] ),
    .Q(_04191_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10508_ (.D(\slice.configuroni.comb_config[58] ),
    .Q(_04192_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10509_ (.D(\slice.configuroni.comb_config[59] ),
    .Q(_04178_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10510_ (.D(\slice.configuroni.comb_config[60] ),
    .Q(_04179_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10511_ (.D(\slice.configuroni.comb_config[61] ),
    .Q(_04180_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10512_ (.D(\slice.configuroni.comb_config[62] ),
    .Q(_04181_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10513_ (.D(\slice.configuroni.comb_config[63] ),
    .Q(_04182_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10514_ (.D(\slice.configuroni.comb_config[64] ),
    .Q(_04183_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10515_ (.D(\slice.configuroni.comb_config[66] ),
    .Q(_04250_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10516_ (.D(\slice.configuroni.comb_config[67] ),
    .Q(_04257_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10517_ (.D(\slice.configuroni.comb_config[68] ),
    .Q(_04258_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10518_ (.D(\slice.configuroni.comb_config[69] ),
    .Q(_04259_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10519_ (.D(\slice.configuroni.comb_config[70] ),
    .Q(_04260_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10520_ (.D(\slice.configuroni.comb_config[71] ),
    .Q(_04261_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10521_ (.D(\slice.configuroni.comb_config[72] ),
    .Q(_04262_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10522_ (.D(\slice.configuroni.comb_config[73] ),
    .Q(_04263_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10523_ (.D(\slice.configuroni.comb_config[74] ),
    .Q(_04264_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10524_ (.D(\slice.configuroni.comb_config[75] ),
    .Q(_04265_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10525_ (.D(\slice.configuroni.comb_config[76] ),
    .Q(_04251_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10526_ (.D(\slice.configuroni.comb_config[77] ),
    .Q(_04252_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10527_ (.D(\slice.configuroni.comb_config[78] ),
    .Q(_04253_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10528_ (.D(\slice.configuroni.comb_config[79] ),
    .Q(_04254_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10529_ (.D(\slice.configuroni.comb_config[80] ),
    .Q(_04255_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10530_ (.D(\slice.configuroni.comb_config[81] ),
    .Q(_04256_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10531_ (.D(\slice.configuroni.comb_config[82] ),
    .Q(_04226_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10532_ (.D(\slice.configuroni.comb_config[83] ),
    .Q(_04233_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10533_ (.D(\slice.configuroni.comb_config[84] ),
    .Q(_04234_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10534_ (.D(\slice.configuroni.comb_config[85] ),
    .Q(_04235_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10535_ (.D(\slice.configuroni.comb_config[86] ),
    .Q(_04236_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10536_ (.D(\slice.configuroni.comb_config[87] ),
    .Q(_04237_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10537_ (.D(\slice.configuroni.comb_config[88] ),
    .Q(_04238_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10538_ (.D(\slice.configuroni.comb_config[89] ),
    .Q(_04239_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10539_ (.D(\slice.configuroni.comb_config[90] ),
    .Q(_04240_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10540_ (.D(\slice.configuroni.comb_config[91] ),
    .Q(_04241_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10541_ (.D(\slice.configuroni.comb_config[92] ),
    .Q(_04227_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10542_ (.D(\slice.configuroni.comb_config[93] ),
    .Q(_04228_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10543_ (.D(\slice.configuroni.comb_config[94] ),
    .Q(_04229_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10544_ (.D(\slice.configuroni.comb_config[95] ),
    .Q(_04230_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10545_ (.D(\slice.configuroni.comb_config[96] ),
    .Q(_04231_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10546_ (.D(\slice.configuroni.comb_config[97] ),
    .Q(_04232_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10547_ (.D(\slice.configuroni.comb_config[99] ),
    .Q(_04299_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10548_ (.D(\slice.configuroni.comb_config[100] ),
    .Q(_04306_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10549_ (.D(\slice.configuroni.comb_config[101] ),
    .Q(_04307_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10550_ (.D(\slice.configuroni.comb_config[102] ),
    .Q(_04308_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10551_ (.D(\slice.configuroni.comb_config[103] ),
    .Q(_04309_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10552_ (.D(\slice.configuroni.comb_config[104] ),
    .Q(_04310_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10553_ (.D(\slice.configuroni.comb_config[105] ),
    .Q(_04311_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10554_ (.D(\slice.configuroni.comb_config[106] ),
    .Q(_04312_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10555_ (.D(\slice.configuroni.comb_config[107] ),
    .Q(_04313_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10556_ (.D(\slice.configuroni.comb_config[108] ),
    .Q(_04314_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10557_ (.D(\slice.configuroni.comb_config[109] ),
    .Q(_04300_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10558_ (.D(\slice.configuroni.comb_config[110] ),
    .Q(_04301_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10559_ (.D(\slice.configuroni.comb_config[111] ),
    .Q(_04302_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10560_ (.D(\slice.configuroni.comb_config[112] ),
    .Q(_04303_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10561_ (.D(\slice.configuroni.comb_config[113] ),
    .Q(_04304_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10562_ (.D(\slice.configuroni.comb_config[114] ),
    .Q(_04305_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10563_ (.D(\slice.configuroni.comb_config[115] ),
    .Q(_04275_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10564_ (.D(\slice.configuroni.comb_config[116] ),
    .Q(_04282_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10565_ (.D(\slice.configuroni.comb_config[117] ),
    .Q(_04283_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10566_ (.D(\slice.configuroni.comb_config[118] ),
    .Q(_04284_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10567_ (.D(\slice.configuroni.comb_config[119] ),
    .Q(_04285_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10568_ (.D(\slice.configuroni.comb_config[120] ),
    .Q(_04286_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10569_ (.D(\slice.configuroni.comb_config[121] ),
    .Q(_04287_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10570_ (.D(\slice.configuroni.comb_config[122] ),
    .Q(_04288_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10571_ (.D(\slice.configuroni.comb_config[123] ),
    .Q(_04289_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10572_ (.D(\slice.configuroni.comb_config[124] ),
    .Q(_04290_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10573_ (.D(\slice.configuroni.comb_config[125] ),
    .Q(_04276_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10574_ (.D(\slice.configuroni.comb_config[126] ),
    .Q(_04277_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10575_ (.D(\slice.configuroni.comb_config[127] ),
    .Q(_04278_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10576_ (.D(\slice.configuroni.comb_config[128] ),
    .Q(_04279_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10577_ (.D(\slice.configuroni.comb_config[129] ),
    .Q(_04280_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10578_ (.D(\slice.configuroni.comb_config[130] ),
    .Q(_04281_),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10579_ (.D(\cb_north.inst.cb_conf_bus[0] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10580_ (.D(\cb_north.inst.cb_conf_bus[1] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10581_ (.D(\cb_north.inst.cb_conf_bus[2] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10582_ (.D(\cb_north.inst.cb_conf_bus[3] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10583_ (.D(\cb_north.inst.cb_conf_bus[4] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10584_ (.D(\cb_north.inst.cb_conf_bus[5] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10585_ (.D(\cb_north.inst.cb_conf_bus[6] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10586_ (.D(\cb_north.inst.cb_conf_bus[7] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10587_ (.D(\cb_north.inst.cb_conf_bus[8] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10588_ (.D(\cb_north.inst.cb_conf_bus[9] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10589_ (.D(\cb_north.inst.cb_conf_bus[10] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10590_ (.D(\cb_north.inst.cb_conf_bus[11] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10591_ (.D(\cb_north.inst.cb_conf_bus[12] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10592_ (.D(\cb_north.inst.cb_conf_bus[13] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10593_ (.D(\cb_north.inst.cb_conf_bus[14] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10594_ (.D(\cb_north.inst.cb_conf_bus[15] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10595_ (.D(\cb_north.inst.cb_conf_bus[16] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[0].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10596_ (.D(\cb_north.inst.cb_conf_bus[17] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10597_ (.D(\cb_north.inst.cb_conf_bus[18] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10598_ (.D(\cb_north.inst.cb_conf_bus[19] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10599_ (.D(\cb_north.inst.cb_conf_bus[20] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10600_ (.D(\cb_north.inst.cb_conf_bus[21] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10601_ (.D(\cb_north.inst.cb_conf_bus[22] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10602_ (.D(\cb_north.inst.cb_conf_bus[23] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10603_ (.D(\cb_north.inst.cb_conf_bus[24] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10604_ (.D(\cb_north.inst.cb_conf_bus[25] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10605_ (.D(\cb_north.inst.cb_conf_bus[26] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10606_ (.D(\cb_north.inst.cb_conf_bus[27] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10607_ (.D(\cb_north.inst.cb_conf_bus[28] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10608_ (.D(\cb_north.inst.cb_conf_bus[29] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10609_ (.D(\cb_north.inst.cb_conf_bus[30] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10610_ (.D(\cb_north.inst.cb_conf_bus[31] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10611_ (.D(\cb_north.inst.cb_conf_bus[32] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10612_ (.D(\cb_north.inst.cb_conf_bus[33] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[1].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10613_ (.D(\cb_north.inst.cb_conf_bus[34] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10614_ (.D(\cb_north.inst.cb_conf_bus[35] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10615_ (.D(\cb_north.inst.cb_conf_bus[36] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10616_ (.D(\cb_north.inst.cb_conf_bus[37] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10617_ (.D(\cb_north.inst.cb_conf_bus[38] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10618_ (.D(\cb_north.inst.cb_conf_bus[39] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10619_ (.D(\cb_north.inst.cb_conf_bus[40] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10620_ (.D(\cb_north.inst.cb_conf_bus[41] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10621_ (.D(\cb_north.inst.cb_conf_bus[42] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10622_ (.D(\cb_north.inst.cb_conf_bus[43] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10623_ (.D(\cb_north.inst.cb_conf_bus[44] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10624_ (.D(\cb_north.inst.cb_conf_bus[45] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10625_ (.D(\cb_north.inst.cb_conf_bus[46] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10626_ (.D(\cb_north.inst.cb_conf_bus[47] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10627_ (.D(\cb_north.inst.cb_conf_bus[48] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10628_ (.D(\cb_north.inst.cb_conf_bus[49] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10629_ (.D(\cb_north.inst.cb_conf_bus[50] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[2].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10630_ (.D(\cb_north.inst.cb_conf_bus[51] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10631_ (.D(\cb_north.inst.cb_conf_bus[52] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10632_ (.D(\cb_north.inst.cb_conf_bus[53] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10633_ (.D(\cb_north.inst.cb_conf_bus[54] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10634_ (.D(\cb_north.inst.cb_conf_bus[55] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10635_ (.D(\cb_north.inst.cb_conf_bus[56] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10636_ (.D(\cb_north.inst.cb_conf_bus[57] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10637_ (.D(\cb_north.inst.cb_conf_bus[58] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10638_ (.D(\cb_north.inst.cb_conf_bus[59] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10639_ (.D(\cb_north.inst.cb_conf_bus[60] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10640_ (.D(\cb_north.inst.cb_conf_bus[61] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10641_ (.D(\cb_north.inst.cb_conf_bus[62] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10642_ (.D(\cb_north.inst.cb_conf_bus[63] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10643_ (.D(\cb_north.inst.cb_conf_bus[64] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10644_ (.D(\cb_north.inst.cb_conf_bus[65] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10645_ (.D(\cb_north.inst.cb_conf_bus[66] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10646_ (.D(\cb_north.inst.cb_conf_bus[67] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[3].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10647_ (.D(\cb_north.inst.cb_conf_bus[68] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10648_ (.D(\cb_north.inst.cb_conf_bus[69] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10649_ (.D(\cb_north.inst.cb_conf_bus[70] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10650_ (.D(\cb_north.inst.cb_conf_bus[71] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10651_ (.D(\cb_north.inst.cb_conf_bus[72] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10652_ (.D(\cb_north.inst.cb_conf_bus[73] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10653_ (.D(\cb_north.inst.cb_conf_bus[74] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10654_ (.D(\cb_north.inst.cb_conf_bus[75] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10655_ (.D(\cb_north.inst.cb_conf_bus[76] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10656_ (.D(\cb_north.inst.cb_conf_bus[77] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10657_ (.D(\cb_north.inst.cb_conf_bus[78] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10658_ (.D(\cb_north.inst.cb_conf_bus[79] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10659_ (.D(\cb_north.inst.cb_conf_bus[80] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10660_ (.D(\cb_north.inst.cb_conf_bus[81] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10661_ (.D(\cb_north.inst.cb_conf_bus[82] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10662_ (.D(\cb_north.inst.cb_conf_bus[83] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10663_ (.D(\cb_north.inst.cb_conf_bus[84] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[4].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10664_ (.D(\cb_north.inst.cb_conf_bus[85] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10665_ (.D(\cb_north.inst.cb_conf_bus[86] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10666_ (.D(\cb_north.inst.cb_conf_bus[87] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10667_ (.D(\cb_north.inst.cb_conf_bus[88] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10668_ (.D(\cb_north.inst.cb_conf_bus[89] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10669_ (.D(\cb_north.inst.cb_conf_bus[90] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10670_ (.D(\cb_north.inst.cb_conf_bus[91] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10671_ (.D(\cb_north.inst.cb_conf_bus[92] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10672_ (.D(\cb_north.inst.cb_conf_bus[93] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10673_ (.D(\cb_north.inst.cb_conf_bus[94] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10674_ (.D(\cb_north.inst.cb_conf_bus[95] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10675_ (.D(\cb_north.inst.cb_conf_bus[96] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10676_ (.D(\cb_north.inst.cb_conf_bus[97] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10677_ (.D(\cb_north.inst.cb_conf_bus[98] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10678_ (.D(\cb_north.inst.cb_conf_bus[99] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10679_ (.D(\cb_north.inst.cb_conf_bus[100] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10680_ (.D(\cb_north.inst.cb_conf_bus[101] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[5].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10681_ (.D(\cb_north.inst.cb_conf_bus[102] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10682_ (.D(\cb_north.inst.cb_conf_bus[103] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10683_ (.D(\cb_north.inst.cb_conf_bus[104] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10684_ (.D(\cb_north.inst.cb_conf_bus[105] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10685_ (.D(\cb_north.inst.cb_conf_bus[106] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10686_ (.D(\cb_north.inst.cb_conf_bus[107] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10687_ (.D(\cb_north.inst.cb_conf_bus[108] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10688_ (.D(\cb_north.inst.cb_conf_bus[109] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10689_ (.D(\cb_north.inst.cb_conf_bus[110] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10690_ (.D(\cb_north.inst.cb_conf_bus[111] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10691_ (.D(\cb_north.inst.cb_conf_bus[112] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10692_ (.D(\cb_north.inst.cb_conf_bus[113] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10693_ (.D(\cb_north.inst.cb_conf_bus[114] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10694_ (.D(\cb_north.inst.cb_conf_bus[115] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10695_ (.D(\cb_north.inst.cb_conf_bus[116] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10696_ (.D(\cb_north.inst.cb_conf_bus[117] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10697_ (.D(\cb_north.inst.cb_conf_bus[118] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[6].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10698_ (.D(\cb_north.inst.cb_conf_bus[119] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10699_ (.D(\cb_north.inst.cb_conf_bus[120] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10700_ (.D(\cb_north.inst.cb_conf_bus[121] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10701_ (.D(\cb_north.inst.cb_conf_bus[122] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10702_ (.D(\cb_north.inst.cb_conf_bus[123] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10703_ (.D(\cb_north.inst.cb_conf_bus[124] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10704_ (.D(\cb_north.inst.cb_conf_bus[125] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10705_ (.D(\cb_north.inst.cb_conf_bus[126] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10706_ (.D(\cb_north.inst.cb_conf_bus[127] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10707_ (.D(\cb_north.inst.cb_conf_bus[128] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10708_ (.D(\cb_north.inst.cb_conf_bus[129] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10709_ (.D(\cb_north.inst.cb_conf_bus[130] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10710_ (.D(\cb_north.inst.cb_conf_bus[131] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10711_ (.D(\cb_north.inst.cb_conf_bus[132] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10712_ (.D(\cb_north.inst.cb_conf_bus[133] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10713_ (.D(\cb_north.inst.cb_conf_bus[134] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10714_ (.D(\cb_north.inst.cb_conf_bus[135] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[7].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10715_ (.D(\cb_north.inst.cb_conf_bus[136] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10716_ (.D(\cb_north.inst.cb_conf_bus[137] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10717_ (.D(\cb_north.inst.cb_conf_bus[138] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10718_ (.D(\cb_north.inst.cb_conf_bus[139] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10719_ (.D(\cb_north.inst.cb_conf_bus[140] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10720_ (.D(\cb_north.inst.cb_conf_bus[141] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10721_ (.D(\cb_north.inst.cb_conf_bus[142] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10722_ (.D(\cb_north.inst.cb_conf_bus[143] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10723_ (.D(\cb_north.inst.cb_conf_bus[144] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10724_ (.D(\cb_north.inst.cb_conf_bus[145] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10725_ (.D(\cb_north.inst.cb_conf_bus[146] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10726_ (.D(\cb_north.inst.cb_conf_bus[147] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10727_ (.D(\cb_north.inst.cb_conf_bus[148] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10728_ (.D(\cb_north.inst.cb_conf_bus[149] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10729_ (.D(\cb_north.inst.cb_conf_bus[150] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10730_ (.D(\cb_north.inst.cb_conf_bus[151] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10731_ (.D(\cb_north.inst.cb_conf_bus[152] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[8].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10732_ (.D(\cb_north.inst.cb_conf_bus[153] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10733_ (.D(\cb_north.inst.cb_conf_bus[154] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10734_ (.D(\cb_north.inst.cb_conf_bus[155] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10735_ (.D(\cb_north.inst.cb_conf_bus[156] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10736_ (.D(\cb_north.inst.cb_conf_bus[157] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10737_ (.D(\cb_north.inst.cb_conf_bus[158] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10738_ (.D(\cb_north.inst.cb_conf_bus[159] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10739_ (.D(\cb_north.inst.cb_conf_bus[160] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10740_ (.D(\cb_north.inst.cb_conf_bus[161] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10741_ (.D(\cb_north.inst.cb_conf_bus[162] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10742_ (.D(\cb_north.inst.cb_conf_bus[163] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10743_ (.D(\cb_north.inst.cb_conf_bus[164] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10744_ (.D(\cb_north.inst.cb_conf_bus[165] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10745_ (.D(\cb_north.inst.cb_conf_bus[166] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10746_ (.D(\cb_north.inst.cb_conf_bus[167] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10747_ (.D(\cb_north.inst.cb_conf_bus[168] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10748_ (.D(\cb_north.inst.cb_conf_bus[169] ),
    .Q(\cb_north.inst.connectaroni.clb0_inputs[9].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10749_ (.D(\cb_north.inst.cb_conf_bus[170] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10750_ (.D(\cb_north.inst.cb_conf_bus[171] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10751_ (.D(\cb_north.inst.cb_conf_bus[172] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10752_ (.D(\cb_north.inst.cb_conf_bus[173] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10753_ (.D(\cb_north.inst.cb_conf_bus[174] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10754_ (.D(\cb_north.inst.cb_conf_bus[175] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10755_ (.D(\cb_north.inst.cb_conf_bus[176] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10756_ (.D(\cb_north.inst.cb_conf_bus[177] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10757_ (.D(\cb_north.inst.cb_conf_bus[178] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10758_ (.D(\cb_north.inst.cb_conf_bus[179] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10759_ (.D(\cb_north.inst.cb_conf_bus[180] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10760_ (.D(\cb_north.inst.cb_conf_bus[181] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10761_ (.D(\cb_north.inst.cb_conf_bus[182] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10762_ (.D(\cb_north.inst.cb_conf_bus[183] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10763_ (.D(\cb_north.inst.cb_conf_bus[184] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10764_ (.D(\cb_north.inst.cb_conf_bus[185] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10765_ (.D(\cb_north.inst.cb_conf_bus[186] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10766_ (.D(\cb_north.inst.cb_conf_bus[187] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10767_ (.D(\cb_north.inst.cb_conf_bus[188] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10768_ (.D(\cb_north.inst.cb_conf_bus[189] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10769_ (.D(\cb_north.inst.cb_conf_bus[190] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10770_ (.D(\cb_north.inst.cb_conf_bus[191] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10771_ (.D(\cb_north.inst.cb_conf_bus[192] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10772_ (.D(\cb_north.inst.cb_conf_bus[193] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10773_ (.D(\cb_north.inst.cb_conf_bus[194] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10774_ (.D(\cb_north.inst.cb_conf_bus[195] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10775_ (.D(\cb_north.inst.cb_conf_bus[196] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10776_ (.D(\cb_north.inst.cb_conf_bus[197] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10777_ (.D(\cb_north.inst.cb_conf_bus[198] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10778_ (.D(\cb_north.inst.cb_conf_bus[199] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10779_ (.D(\cb_north.inst.cb_conf_bus[200] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10780_ (.D(\cb_north.inst.cb_conf_bus[201] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10781_ (.D(\cb_north.inst.cb_conf_bus[202] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10782_ (.D(\cb_north.inst.cb_conf_bus[203] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10783_ (.D(\cb_north.inst.cb_conf_bus[204] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10784_ (.D(\cb_north.inst.cb_conf_bus[205] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10785_ (.D(\cb_north.inst.cb_conf_bus[206] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10786_ (.D(\cb_north.inst.cb_conf_bus[207] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10787_ (.D(\cb_north.inst.cb_conf_bus[208] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10788_ (.D(\cb_north.inst.cb_conf_bus[209] ),
    .Q(\cb_north.inst.connectaroni.clb0_outputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10789_ (.D(\cb_north.inst.cb_conf_bus[210] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10790_ (.D(\cb_north.inst.cb_conf_bus[211] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10791_ (.D(\cb_north.inst.cb_conf_bus[212] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10792_ (.D(\cb_north.inst.cb_conf_bus[213] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10793_ (.D(\cb_north.inst.cb_conf_bus[214] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10794_ (.D(\cb_north.inst.cb_conf_bus[215] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10795_ (.D(\cb_north.inst.cb_conf_bus[216] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10796_ (.D(\cb_north.inst.cb_conf_bus[217] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10797_ (.D(\cb_north.inst.cb_conf_bus[218] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10798_ (.D(\cb_north.inst.cb_conf_bus[219] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10799_ (.D(\cb_north.inst.cb_conf_bus[220] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10800_ (.D(\cb_north.inst.cb_conf_bus[221] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10801_ (.D(\cb_north.inst.cb_conf_bus[222] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10802_ (.D(\cb_north.inst.cb_conf_bus[223] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10803_ (.D(\cb_north.inst.cb_conf_bus[224] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10804_ (.D(\cb_north.inst.cb_conf_bus[225] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10805_ (.D(\cb_north.inst.cb_conf_bus[226] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[0].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10806_ (.D(\cb_north.inst.cb_conf_bus[227] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10807_ (.D(\cb_north.inst.cb_conf_bus[228] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10808_ (.D(\cb_north.inst.cb_conf_bus[229] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10809_ (.D(\cb_north.inst.cb_conf_bus[230] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10810_ (.D(\cb_north.inst.cb_conf_bus[231] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10811_ (.D(\cb_north.inst.cb_conf_bus[232] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10812_ (.D(\cb_north.inst.cb_conf_bus[233] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10813_ (.D(\cb_north.inst.cb_conf_bus[234] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10814_ (.D(\cb_north.inst.cb_conf_bus[235] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10815_ (.D(\cb_north.inst.cb_conf_bus[236] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10816_ (.D(\cb_north.inst.cb_conf_bus[237] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10817_ (.D(\cb_north.inst.cb_conf_bus[238] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10818_ (.D(\cb_north.inst.cb_conf_bus[239] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10819_ (.D(\cb_north.inst.cb_conf_bus[240] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10820_ (.D(\cb_north.inst.cb_conf_bus[241] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10821_ (.D(\cb_north.inst.cb_conf_bus[242] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10822_ (.D(\cb_north.inst.cb_conf_bus[243] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[1].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10823_ (.D(\cb_north.inst.cb_conf_bus[244] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10824_ (.D(\cb_north.inst.cb_conf_bus[245] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10825_ (.D(\cb_north.inst.cb_conf_bus[246] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10826_ (.D(\cb_north.inst.cb_conf_bus[247] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10827_ (.D(\cb_north.inst.cb_conf_bus[248] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10828_ (.D(\cb_north.inst.cb_conf_bus[249] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10829_ (.D(\cb_north.inst.cb_conf_bus[250] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10830_ (.D(\cb_north.inst.cb_conf_bus[251] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10831_ (.D(\cb_north.inst.cb_conf_bus[252] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10832_ (.D(\cb_north.inst.cb_conf_bus[253] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10833_ (.D(\cb_north.inst.cb_conf_bus[254] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10834_ (.D(\cb_north.inst.cb_conf_bus[255] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10835_ (.D(\cb_north.inst.cb_conf_bus[256] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10836_ (.D(\cb_north.inst.cb_conf_bus[257] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10837_ (.D(\cb_north.inst.cb_conf_bus[258] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10838_ (.D(\cb_north.inst.cb_conf_bus[259] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10839_ (.D(\cb_north.inst.cb_conf_bus[260] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[2].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10840_ (.D(\cb_north.inst.cb_conf_bus[261] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10841_ (.D(\cb_north.inst.cb_conf_bus[262] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10842_ (.D(\cb_north.inst.cb_conf_bus[263] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10843_ (.D(\cb_north.inst.cb_conf_bus[264] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10844_ (.D(\cb_north.inst.cb_conf_bus[265] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10845_ (.D(\cb_north.inst.cb_conf_bus[266] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10846_ (.D(\cb_north.inst.cb_conf_bus[267] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10847_ (.D(\cb_north.inst.cb_conf_bus[268] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10848_ (.D(\cb_north.inst.cb_conf_bus[269] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10849_ (.D(\cb_north.inst.cb_conf_bus[270] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10850_ (.D(\cb_north.inst.cb_conf_bus[271] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10851_ (.D(\cb_north.inst.cb_conf_bus[272] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10852_ (.D(\cb_north.inst.cb_conf_bus[273] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10853_ (.D(\cb_north.inst.cb_conf_bus[274] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10854_ (.D(\cb_north.inst.cb_conf_bus[275] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10855_ (.D(\cb_north.inst.cb_conf_bus[276] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10856_ (.D(\cb_north.inst.cb_conf_bus[277] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[3].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10857_ (.D(\cb_north.inst.cb_conf_bus[278] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10858_ (.D(\cb_north.inst.cb_conf_bus[279] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10859_ (.D(\cb_north.inst.cb_conf_bus[280] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10860_ (.D(\cb_north.inst.cb_conf_bus[281] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10861_ (.D(\cb_north.inst.cb_conf_bus[282] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10862_ (.D(\cb_north.inst.cb_conf_bus[283] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10863_ (.D(\cb_north.inst.cb_conf_bus[284] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10864_ (.D(\cb_north.inst.cb_conf_bus[285] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10865_ (.D(\cb_north.inst.cb_conf_bus[286] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10866_ (.D(\cb_north.inst.cb_conf_bus[287] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10867_ (.D(\cb_north.inst.cb_conf_bus[288] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10868_ (.D(\cb_north.inst.cb_conf_bus[289] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10869_ (.D(\cb_north.inst.cb_conf_bus[290] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10870_ (.D(\cb_north.inst.cb_conf_bus[291] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10871_ (.D(\cb_north.inst.cb_conf_bus[292] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10872_ (.D(\cb_north.inst.cb_conf_bus[293] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10873_ (.D(\cb_north.inst.cb_conf_bus[294] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[4].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10874_ (.D(\cb_north.inst.cb_conf_bus[295] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10875_ (.D(\cb_north.inst.cb_conf_bus[296] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10876_ (.D(\cb_north.inst.cb_conf_bus[297] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10877_ (.D(\cb_north.inst.cb_conf_bus[298] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10878_ (.D(\cb_north.inst.cb_conf_bus[299] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10879_ (.D(\cb_north.inst.cb_conf_bus[300] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10880_ (.D(\cb_north.inst.cb_conf_bus[301] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10881_ (.D(\cb_north.inst.cb_conf_bus[302] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10882_ (.D(\cb_north.inst.cb_conf_bus[303] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10883_ (.D(\cb_north.inst.cb_conf_bus[304] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10884_ (.D(\cb_north.inst.cb_conf_bus[305] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10885_ (.D(\cb_north.inst.cb_conf_bus[306] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10886_ (.D(\cb_north.inst.cb_conf_bus[307] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10887_ (.D(\cb_north.inst.cb_conf_bus[308] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10888_ (.D(\cb_north.inst.cb_conf_bus[309] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10889_ (.D(\cb_north.inst.cb_conf_bus[310] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10890_ (.D(\cb_north.inst.cb_conf_bus[311] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[5].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10891_ (.D(\cb_north.inst.cb_conf_bus[312] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10892_ (.D(\cb_north.inst.cb_conf_bus[313] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10893_ (.D(\cb_north.inst.cb_conf_bus[314] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10894_ (.D(\cb_north.inst.cb_conf_bus[315] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10895_ (.D(\cb_north.inst.cb_conf_bus[316] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10896_ (.D(\cb_north.inst.cb_conf_bus[317] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10897_ (.D(\cb_north.inst.cb_conf_bus[318] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10898_ (.D(\cb_north.inst.cb_conf_bus[319] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10899_ (.D(\cb_north.inst.cb_conf_bus[320] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10900_ (.D(\cb_north.inst.cb_conf_bus[321] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10901_ (.D(\cb_north.inst.cb_conf_bus[322] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10902_ (.D(\cb_north.inst.cb_conf_bus[323] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10903_ (.D(\cb_north.inst.cb_conf_bus[324] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10904_ (.D(\cb_north.inst.cb_conf_bus[325] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10905_ (.D(\cb_north.inst.cb_conf_bus[326] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10906_ (.D(\cb_north.inst.cb_conf_bus[327] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10907_ (.D(\cb_north.inst.cb_conf_bus[328] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[6].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10908_ (.D(\cb_north.inst.cb_conf_bus[329] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10909_ (.D(\cb_north.inst.cb_conf_bus[330] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10910_ (.D(\cb_north.inst.cb_conf_bus[331] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10911_ (.D(\cb_north.inst.cb_conf_bus[332] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10912_ (.D(\cb_north.inst.cb_conf_bus[333] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10913_ (.D(\cb_north.inst.cb_conf_bus[334] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10914_ (.D(\cb_north.inst.cb_conf_bus[335] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10915_ (.D(\cb_north.inst.cb_conf_bus[336] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10916_ (.D(\cb_north.inst.cb_conf_bus[337] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10917_ (.D(\cb_north.inst.cb_conf_bus[338] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10918_ (.D(\cb_north.inst.cb_conf_bus[339] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10919_ (.D(\cb_north.inst.cb_conf_bus[340] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10920_ (.D(\cb_north.inst.cb_conf_bus[341] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10921_ (.D(\cb_north.inst.cb_conf_bus[342] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10922_ (.D(\cb_north.inst.cb_conf_bus[343] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10923_ (.D(\cb_north.inst.cb_conf_bus[344] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10924_ (.D(\cb_north.inst.cb_conf_bus[345] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[7].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10925_ (.D(\cb_north.inst.cb_conf_bus[346] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10926_ (.D(\cb_north.inst.cb_conf_bus[347] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10927_ (.D(\cb_north.inst.cb_conf_bus[348] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10928_ (.D(\cb_north.inst.cb_conf_bus[349] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10929_ (.D(\cb_north.inst.cb_conf_bus[350] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10930_ (.D(\cb_north.inst.cb_conf_bus[351] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10931_ (.D(\cb_north.inst.cb_conf_bus[352] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10932_ (.D(\cb_north.inst.cb_conf_bus[353] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10933_ (.D(\cb_north.inst.cb_conf_bus[354] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10934_ (.D(\cb_north.inst.cb_conf_bus[355] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10935_ (.D(\cb_north.inst.cb_conf_bus[356] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10936_ (.D(\cb_north.inst.cb_conf_bus[357] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10937_ (.D(\cb_north.inst.cb_conf_bus[358] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10938_ (.D(\cb_north.inst.cb_conf_bus[359] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10939_ (.D(\cb_north.inst.cb_conf_bus[360] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10940_ (.D(\cb_north.inst.cb_conf_bus[361] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10941_ (.D(\cb_north.inst.cb_conf_bus[362] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[8].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10942_ (.D(\cb_north.inst.cb_conf_bus[363] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10943_ (.D(\cb_north.inst.cb_conf_bus[364] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10944_ (.D(\cb_north.inst.cb_conf_bus[365] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10945_ (.D(\cb_north.inst.cb_conf_bus[366] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10946_ (.D(\cb_north.inst.cb_conf_bus[367] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10947_ (.D(\cb_north.inst.cb_conf_bus[368] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10948_ (.D(\cb_north.inst.cb_conf_bus[369] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10949_ (.D(\cb_north.inst.cb_conf_bus[370] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10950_ (.D(\cb_north.inst.cb_conf_bus[371] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10951_ (.D(\cb_north.inst.cb_conf_bus[372] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10952_ (.D(\cb_north.inst.cb_conf_bus[373] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10953_ (.D(\cb_north.inst.cb_conf_bus[374] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10954_ (.D(\cb_north.inst.cb_conf_bus[375] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10955_ (.D(\cb_north.inst.cb_conf_bus[376] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10956_ (.D(\cb_north.inst.cb_conf_bus[377] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10957_ (.D(\cb_north.inst.cb_conf_bus[378] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10958_ (.D(\cb_north.inst.cb_conf_bus[379] ),
    .Q(\cb_north.inst.connectaroni.clb1_inputs[9].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10959_ (.D(\cb_north.inst.cb_conf_bus[380] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10960_ (.D(\cb_north.inst.cb_conf_bus[381] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10961_ (.D(\cb_north.inst.cb_conf_bus[382] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10962_ (.D(\cb_north.inst.cb_conf_bus[383] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10963_ (.D(\cb_north.inst.cb_conf_bus[384] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10964_ (.D(\cb_north.inst.cb_conf_bus[385] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10965_ (.D(\cb_north.inst.cb_conf_bus[386] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10966_ (.D(\cb_north.inst.cb_conf_bus[387] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10967_ (.D(\cb_north.inst.cb_conf_bus[388] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10968_ (.D(\cb_north.inst.cb_conf_bus[389] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10969_ (.D(\cb_north.inst.cb_conf_bus[390] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10970_ (.D(\cb_north.inst.cb_conf_bus[391] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10971_ (.D(\cb_north.inst.cb_conf_bus[392] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10972_ (.D(\cb_north.inst.cb_conf_bus[393] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10973_ (.D(\cb_north.inst.cb_conf_bus[394] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10974_ (.D(\cb_north.inst.cb_conf_bus[395] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10975_ (.D(\cb_north.inst.cb_conf_bus[396] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10976_ (.D(\cb_north.inst.cb_conf_bus[397] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10977_ (.D(\cb_north.inst.cb_conf_bus[398] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10978_ (.D(\cb_north.inst.cb_conf_bus[399] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10979_ (.D(\cb_north.inst.cb_conf_bus[400] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10980_ (.D(\cb_north.inst.cb_conf_bus[401] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10981_ (.D(\cb_north.inst.cb_conf_bus[402] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10982_ (.D(\cb_north.inst.cb_conf_bus[403] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10983_ (.D(\cb_north.inst.cb_conf_bus[404] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10984_ (.D(\cb_north.inst.cb_conf_bus[405] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10985_ (.D(\cb_north.inst.cb_conf_bus[406] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10986_ (.D(\cb_north.inst.cb_conf_bus[407] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10987_ (.D(\cb_north.inst.cb_conf_bus[408] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10988_ (.D(\cb_north.inst.cb_conf_bus[409] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10989_ (.D(\cb_north.inst.cb_conf_bus[410] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10990_ (.D(\cb_north.inst.cb_conf_bus[411] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10991_ (.D(\cb_north.inst.cb_conf_bus[412] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10992_ (.D(\cb_north.inst.cb_conf_bus[413] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10993_ (.D(\cb_north.inst.cb_conf_bus[414] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10994_ (.D(\cb_north.inst.cb_conf_bus[415] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10995_ (.D(\cb_north.inst.cb_conf_bus[416] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10996_ (.D(\cb_north.inst.cb_conf_bus[417] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10997_ (.D(\cb_north.inst.cb_conf_bus[418] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10998_ (.D(\cb_north.inst.cb_conf_bus[419] ),
    .Q(\cb_north.inst.connectaroni.clb1_outputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _10999_ (.D(shift_out_hard),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11000_ (.D(\cb_east.inst.cb_conf_bus[1] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11001_ (.D(\cb_east.inst.cb_conf_bus[2] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11002_ (.D(\cb_east.inst.cb_conf_bus[3] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11003_ (.D(\cb_east.inst.cb_conf_bus[4] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11004_ (.D(\cb_east.inst.cb_conf_bus[5] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11005_ (.D(\cb_east.inst.cb_conf_bus[6] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11006_ (.D(\cb_east.inst.cb_conf_bus[7] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11007_ (.D(\cb_east.inst.cb_conf_bus[8] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11008_ (.D(\cb_east.inst.cb_conf_bus[9] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11009_ (.D(\cb_east.inst.cb_conf_bus[10] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11010_ (.D(\cb_east.inst.cb_conf_bus[11] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11011_ (.D(\cb_east.inst.cb_conf_bus[12] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11012_ (.D(\cb_east.inst.cb_conf_bus[13] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11013_ (.D(\cb_east.inst.cb_conf_bus[14] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11014_ (.D(\cb_east.inst.cb_conf_bus[15] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11015_ (.D(\cb_east.inst.cb_conf_bus[16] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[0].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11016_ (.D(\cb_east.inst.cb_conf_bus[17] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11017_ (.D(\cb_east.inst.cb_conf_bus[18] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11018_ (.D(\cb_east.inst.cb_conf_bus[19] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11019_ (.D(\cb_east.inst.cb_conf_bus[20] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11020_ (.D(\cb_east.inst.cb_conf_bus[21] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11021_ (.D(\cb_east.inst.cb_conf_bus[22] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11022_ (.D(\cb_east.inst.cb_conf_bus[23] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11023_ (.D(\cb_east.inst.cb_conf_bus[24] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11024_ (.D(\cb_east.inst.cb_conf_bus[25] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11025_ (.D(\cb_east.inst.cb_conf_bus[26] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11026_ (.D(\cb_east.inst.cb_conf_bus[27] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11027_ (.D(\cb_east.inst.cb_conf_bus[28] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11028_ (.D(\cb_east.inst.cb_conf_bus[29] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11029_ (.D(\cb_east.inst.cb_conf_bus[30] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11030_ (.D(\cb_east.inst.cb_conf_bus[31] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11031_ (.D(\cb_east.inst.cb_conf_bus[32] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11032_ (.D(\cb_east.inst.cb_conf_bus[33] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[1].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11033_ (.D(\cb_east.inst.cb_conf_bus[34] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11034_ (.D(\cb_east.inst.cb_conf_bus[35] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11035_ (.D(\cb_east.inst.cb_conf_bus[36] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11036_ (.D(\cb_east.inst.cb_conf_bus[37] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11037_ (.D(\cb_east.inst.cb_conf_bus[38] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11038_ (.D(\cb_east.inst.cb_conf_bus[39] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11039_ (.D(\cb_east.inst.cb_conf_bus[40] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11040_ (.D(\cb_east.inst.cb_conf_bus[41] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11041_ (.D(\cb_east.inst.cb_conf_bus[42] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11042_ (.D(\cb_east.inst.cb_conf_bus[43] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11043_ (.D(\cb_east.inst.cb_conf_bus[44] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11044_ (.D(\cb_east.inst.cb_conf_bus[45] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11045_ (.D(\cb_east.inst.cb_conf_bus[46] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11046_ (.D(\cb_east.inst.cb_conf_bus[47] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11047_ (.D(\cb_east.inst.cb_conf_bus[48] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11048_ (.D(\cb_east.inst.cb_conf_bus[49] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11049_ (.D(\cb_east.inst.cb_conf_bus[50] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[2].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11050_ (.D(\cb_east.inst.cb_conf_bus[51] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11051_ (.D(\cb_east.inst.cb_conf_bus[52] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11052_ (.D(\cb_east.inst.cb_conf_bus[53] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11053_ (.D(\cb_east.inst.cb_conf_bus[54] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11054_ (.D(\cb_east.inst.cb_conf_bus[55] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11055_ (.D(\cb_east.inst.cb_conf_bus[56] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11056_ (.D(\cb_east.inst.cb_conf_bus[57] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11057_ (.D(\cb_east.inst.cb_conf_bus[58] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11058_ (.D(\cb_east.inst.cb_conf_bus[59] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11059_ (.D(\cb_east.inst.cb_conf_bus[60] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11060_ (.D(\cb_east.inst.cb_conf_bus[61] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11061_ (.D(\cb_east.inst.cb_conf_bus[62] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11062_ (.D(\cb_east.inst.cb_conf_bus[63] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11063_ (.D(\cb_east.inst.cb_conf_bus[64] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11064_ (.D(\cb_east.inst.cb_conf_bus[65] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11065_ (.D(\cb_east.inst.cb_conf_bus[66] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11066_ (.D(\cb_east.inst.cb_conf_bus[67] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[3].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11067_ (.D(\cb_east.inst.cb_conf_bus[68] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11068_ (.D(\cb_east.inst.cb_conf_bus[69] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11069_ (.D(\cb_east.inst.cb_conf_bus[70] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11070_ (.D(\cb_east.inst.cb_conf_bus[71] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11071_ (.D(\cb_east.inst.cb_conf_bus[72] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11072_ (.D(\cb_east.inst.cb_conf_bus[73] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11073_ (.D(\cb_east.inst.cb_conf_bus[74] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11074_ (.D(\cb_east.inst.cb_conf_bus[75] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11075_ (.D(\cb_east.inst.cb_conf_bus[76] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11076_ (.D(\cb_east.inst.cb_conf_bus[77] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11077_ (.D(\cb_east.inst.cb_conf_bus[78] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11078_ (.D(\cb_east.inst.cb_conf_bus[79] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11079_ (.D(\cb_east.inst.cb_conf_bus[80] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11080_ (.D(\cb_east.inst.cb_conf_bus[81] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11081_ (.D(\cb_east.inst.cb_conf_bus[82] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11082_ (.D(\cb_east.inst.cb_conf_bus[83] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11083_ (.D(\cb_east.inst.cb_conf_bus[84] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[4].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11084_ (.D(\cb_east.inst.cb_conf_bus[85] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11085_ (.D(\cb_east.inst.cb_conf_bus[86] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11086_ (.D(\cb_east.inst.cb_conf_bus[87] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11087_ (.D(\cb_east.inst.cb_conf_bus[88] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11088_ (.D(\cb_east.inst.cb_conf_bus[89] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11089_ (.D(\cb_east.inst.cb_conf_bus[90] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11090_ (.D(\cb_east.inst.cb_conf_bus[91] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11091_ (.D(\cb_east.inst.cb_conf_bus[92] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11092_ (.D(\cb_east.inst.cb_conf_bus[93] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11093_ (.D(\cb_east.inst.cb_conf_bus[94] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11094_ (.D(\cb_east.inst.cb_conf_bus[95] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11095_ (.D(\cb_east.inst.cb_conf_bus[96] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11096_ (.D(\cb_east.inst.cb_conf_bus[97] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11097_ (.D(\cb_east.inst.cb_conf_bus[98] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11098_ (.D(\cb_east.inst.cb_conf_bus[99] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11099_ (.D(\cb_east.inst.cb_conf_bus[100] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11100_ (.D(\cb_east.inst.cb_conf_bus[101] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[5].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11101_ (.D(\cb_east.inst.cb_conf_bus[102] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11102_ (.D(\cb_east.inst.cb_conf_bus[103] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11103_ (.D(\cb_east.inst.cb_conf_bus[104] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11104_ (.D(\cb_east.inst.cb_conf_bus[105] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11105_ (.D(\cb_east.inst.cb_conf_bus[106] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11106_ (.D(\cb_east.inst.cb_conf_bus[107] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11107_ (.D(\cb_east.inst.cb_conf_bus[108] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11108_ (.D(\cb_east.inst.cb_conf_bus[109] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11109_ (.D(\cb_east.inst.cb_conf_bus[110] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11110_ (.D(\cb_east.inst.cb_conf_bus[111] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11111_ (.D(\cb_east.inst.cb_conf_bus[112] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11112_ (.D(\cb_east.inst.cb_conf_bus[113] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11113_ (.D(\cb_east.inst.cb_conf_bus[114] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11114_ (.D(\cb_east.inst.cb_conf_bus[115] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11115_ (.D(\cb_east.inst.cb_conf_bus[116] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11116_ (.D(\cb_east.inst.cb_conf_bus[117] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11117_ (.D(\cb_east.inst.cb_conf_bus[118] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[6].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11118_ (.D(\cb_east.inst.cb_conf_bus[119] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11119_ (.D(\cb_east.inst.cb_conf_bus[120] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11120_ (.D(\cb_east.inst.cb_conf_bus[121] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11121_ (.D(\cb_east.inst.cb_conf_bus[122] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11122_ (.D(\cb_east.inst.cb_conf_bus[123] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11123_ (.D(\cb_east.inst.cb_conf_bus[124] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11124_ (.D(\cb_east.inst.cb_conf_bus[125] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11125_ (.D(\cb_east.inst.cb_conf_bus[126] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11126_ (.D(\cb_east.inst.cb_conf_bus[127] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11127_ (.D(\cb_east.inst.cb_conf_bus[128] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11128_ (.D(\cb_east.inst.cb_conf_bus[129] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11129_ (.D(\cb_east.inst.cb_conf_bus[130] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11130_ (.D(\cb_east.inst.cb_conf_bus[131] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11131_ (.D(\cb_east.inst.cb_conf_bus[132] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11132_ (.D(\cb_east.inst.cb_conf_bus[133] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11133_ (.D(\cb_east.inst.cb_conf_bus[134] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11134_ (.D(\cb_east.inst.cb_conf_bus[135] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[7].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11135_ (.D(\cb_east.inst.cb_conf_bus[136] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11136_ (.D(\cb_east.inst.cb_conf_bus[137] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11137_ (.D(\cb_east.inst.cb_conf_bus[138] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11138_ (.D(\cb_east.inst.cb_conf_bus[139] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11139_ (.D(\cb_east.inst.cb_conf_bus[140] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11140_ (.D(\cb_east.inst.cb_conf_bus[141] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11141_ (.D(\cb_east.inst.cb_conf_bus[142] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11142_ (.D(\cb_east.inst.cb_conf_bus[143] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11143_ (.D(\cb_east.inst.cb_conf_bus[144] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11144_ (.D(\cb_east.inst.cb_conf_bus[145] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11145_ (.D(\cb_east.inst.cb_conf_bus[146] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11146_ (.D(\cb_east.inst.cb_conf_bus[147] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11147_ (.D(\cb_east.inst.cb_conf_bus[148] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11148_ (.D(\cb_east.inst.cb_conf_bus[149] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11149_ (.D(\cb_east.inst.cb_conf_bus[150] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11150_ (.D(\cb_east.inst.cb_conf_bus[151] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11151_ (.D(\cb_east.inst.cb_conf_bus[152] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[8].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11152_ (.D(\cb_east.inst.cb_conf_bus[153] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11153_ (.D(\cb_east.inst.cb_conf_bus[154] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11154_ (.D(\cb_east.inst.cb_conf_bus[155] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11155_ (.D(\cb_east.inst.cb_conf_bus[156] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11156_ (.D(\cb_east.inst.cb_conf_bus[157] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11157_ (.D(\cb_east.inst.cb_conf_bus[158] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11158_ (.D(\cb_east.inst.cb_conf_bus[159] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11159_ (.D(\cb_east.inst.cb_conf_bus[160] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11160_ (.D(\cb_east.inst.cb_conf_bus[161] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11161_ (.D(\cb_east.inst.cb_conf_bus[162] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11162_ (.D(\cb_east.inst.cb_conf_bus[163] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11163_ (.D(\cb_east.inst.cb_conf_bus[164] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11164_ (.D(\cb_east.inst.cb_conf_bus[165] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11165_ (.D(\cb_east.inst.cb_conf_bus[166] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11166_ (.D(\cb_east.inst.cb_conf_bus[167] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11167_ (.D(\cb_east.inst.cb_conf_bus[168] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11168_ (.D(\cb_east.inst.cb_conf_bus[169] ),
    .Q(\cb_east.inst.connectaroni.clb0_inputs[9].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11169_ (.D(\cb_east.inst.cb_conf_bus[170] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11170_ (.D(\cb_east.inst.cb_conf_bus[171] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11171_ (.D(\cb_east.inst.cb_conf_bus[172] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11172_ (.D(\cb_east.inst.cb_conf_bus[173] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11173_ (.D(\cb_east.inst.cb_conf_bus[174] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11174_ (.D(\cb_east.inst.cb_conf_bus[175] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11175_ (.D(\cb_east.inst.cb_conf_bus[176] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11176_ (.D(\cb_east.inst.cb_conf_bus[177] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11177_ (.D(\cb_east.inst.cb_conf_bus[178] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11178_ (.D(\cb_east.inst.cb_conf_bus[179] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11179_ (.D(\cb_east.inst.cb_conf_bus[180] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11180_ (.D(\cb_east.inst.cb_conf_bus[181] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11181_ (.D(\cb_east.inst.cb_conf_bus[182] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11182_ (.D(\cb_east.inst.cb_conf_bus[183] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11183_ (.D(\cb_east.inst.cb_conf_bus[184] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11184_ (.D(\cb_east.inst.cb_conf_bus[185] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11185_ (.D(\cb_east.inst.cb_conf_bus[186] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11186_ (.D(\cb_east.inst.cb_conf_bus[187] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11187_ (.D(\cb_east.inst.cb_conf_bus[188] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11188_ (.D(\cb_east.inst.cb_conf_bus[189] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11189_ (.D(\cb_east.inst.cb_conf_bus[190] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11190_ (.D(\cb_east.inst.cb_conf_bus[191] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11191_ (.D(\cb_east.inst.cb_conf_bus[192] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11192_ (.D(\cb_east.inst.cb_conf_bus[193] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11193_ (.D(\cb_east.inst.cb_conf_bus[194] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11194_ (.D(\cb_east.inst.cb_conf_bus[195] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11195_ (.D(\cb_east.inst.cb_conf_bus[196] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11196_ (.D(\cb_east.inst.cb_conf_bus[197] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11197_ (.D(\cb_east.inst.cb_conf_bus[198] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11198_ (.D(\cb_east.inst.cb_conf_bus[199] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11199_ (.D(\cb_east.inst.cb_conf_bus[200] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11200_ (.D(\cb_east.inst.cb_conf_bus[201] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11201_ (.D(\cb_east.inst.cb_conf_bus[202] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11202_ (.D(\cb_east.inst.cb_conf_bus[203] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11203_ (.D(\cb_east.inst.cb_conf_bus[204] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11204_ (.D(\cb_east.inst.cb_conf_bus[205] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11205_ (.D(\cb_east.inst.cb_conf_bus[206] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11206_ (.D(\cb_east.inst.cb_conf_bus[207] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11207_ (.D(\cb_east.inst.cb_conf_bus[208] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11208_ (.D(\cb_east.inst.cb_conf_bus[209] ),
    .Q(\cb_east.inst.connectaroni.clb0_outputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11209_ (.D(\cb_east.inst.cb_conf_bus[210] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11210_ (.D(\cb_east.inst.cb_conf_bus[211] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11211_ (.D(\cb_east.inst.cb_conf_bus[212] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11212_ (.D(\cb_east.inst.cb_conf_bus[213] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11213_ (.D(\cb_east.inst.cb_conf_bus[214] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11214_ (.D(\cb_east.inst.cb_conf_bus[215] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11215_ (.D(\cb_east.inst.cb_conf_bus[216] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11216_ (.D(\cb_east.inst.cb_conf_bus[217] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11217_ (.D(\cb_east.inst.cb_conf_bus[218] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11218_ (.D(\cb_east.inst.cb_conf_bus[219] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11219_ (.D(\cb_east.inst.cb_conf_bus[220] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11220_ (.D(\cb_east.inst.cb_conf_bus[221] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11221_ (.D(\cb_east.inst.cb_conf_bus[222] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11222_ (.D(\cb_east.inst.cb_conf_bus[223] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11223_ (.D(\cb_east.inst.cb_conf_bus[224] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11224_ (.D(\cb_east.inst.cb_conf_bus[225] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11225_ (.D(\cb_east.inst.cb_conf_bus[226] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[0].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11226_ (.D(\cb_east.inst.cb_conf_bus[227] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11227_ (.D(\cb_east.inst.cb_conf_bus[228] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11228_ (.D(\cb_east.inst.cb_conf_bus[229] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11229_ (.D(\cb_east.inst.cb_conf_bus[230] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11230_ (.D(\cb_east.inst.cb_conf_bus[231] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11231_ (.D(\cb_east.inst.cb_conf_bus[232] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11232_ (.D(\cb_east.inst.cb_conf_bus[233] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11233_ (.D(\cb_east.inst.cb_conf_bus[234] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11234_ (.D(\cb_east.inst.cb_conf_bus[235] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11235_ (.D(\cb_east.inst.cb_conf_bus[236] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11236_ (.D(\cb_east.inst.cb_conf_bus[237] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11237_ (.D(\cb_east.inst.cb_conf_bus[238] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11238_ (.D(\cb_east.inst.cb_conf_bus[239] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11239_ (.D(\cb_east.inst.cb_conf_bus[240] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11240_ (.D(\cb_east.inst.cb_conf_bus[241] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11241_ (.D(\cb_east.inst.cb_conf_bus[242] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11242_ (.D(\cb_east.inst.cb_conf_bus[243] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[1].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11243_ (.D(\cb_east.inst.cb_conf_bus[244] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11244_ (.D(\cb_east.inst.cb_conf_bus[245] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11245_ (.D(\cb_east.inst.cb_conf_bus[246] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11246_ (.D(\cb_east.inst.cb_conf_bus[247] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11247_ (.D(\cb_east.inst.cb_conf_bus[248] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11248_ (.D(\cb_east.inst.cb_conf_bus[249] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11249_ (.D(\cb_east.inst.cb_conf_bus[250] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11250_ (.D(\cb_east.inst.cb_conf_bus[251] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11251_ (.D(\cb_east.inst.cb_conf_bus[252] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11252_ (.D(\cb_east.inst.cb_conf_bus[253] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11253_ (.D(\cb_east.inst.cb_conf_bus[254] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11254_ (.D(\cb_east.inst.cb_conf_bus[255] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11255_ (.D(\cb_east.inst.cb_conf_bus[256] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11256_ (.D(\cb_east.inst.cb_conf_bus[257] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11257_ (.D(\cb_east.inst.cb_conf_bus[258] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11258_ (.D(\cb_east.inst.cb_conf_bus[259] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11259_ (.D(\cb_east.inst.cb_conf_bus[260] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[2].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11260_ (.D(\cb_east.inst.cb_conf_bus[261] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11261_ (.D(\cb_east.inst.cb_conf_bus[262] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11262_ (.D(\cb_east.inst.cb_conf_bus[263] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11263_ (.D(\cb_east.inst.cb_conf_bus[264] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11264_ (.D(\cb_east.inst.cb_conf_bus[265] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11265_ (.D(\cb_east.inst.cb_conf_bus[266] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11266_ (.D(\cb_east.inst.cb_conf_bus[267] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11267_ (.D(\cb_east.inst.cb_conf_bus[268] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11268_ (.D(\cb_east.inst.cb_conf_bus[269] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11269_ (.D(\cb_east.inst.cb_conf_bus[270] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11270_ (.D(\cb_east.inst.cb_conf_bus[271] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11271_ (.D(\cb_east.inst.cb_conf_bus[272] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11272_ (.D(\cb_east.inst.cb_conf_bus[273] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11273_ (.D(\cb_east.inst.cb_conf_bus[274] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11274_ (.D(\cb_east.inst.cb_conf_bus[275] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11275_ (.D(\cb_east.inst.cb_conf_bus[276] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11276_ (.D(\cb_east.inst.cb_conf_bus[277] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[3].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11277_ (.D(\cb_east.inst.cb_conf_bus[278] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11278_ (.D(\cb_east.inst.cb_conf_bus[279] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11279_ (.D(\cb_east.inst.cb_conf_bus[280] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11280_ (.D(\cb_east.inst.cb_conf_bus[281] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11281_ (.D(\cb_east.inst.cb_conf_bus[282] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11282_ (.D(\cb_east.inst.cb_conf_bus[283] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11283_ (.D(\cb_east.inst.cb_conf_bus[284] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11284_ (.D(\cb_east.inst.cb_conf_bus[285] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11285_ (.D(\cb_east.inst.cb_conf_bus[286] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11286_ (.D(\cb_east.inst.cb_conf_bus[287] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11287_ (.D(\cb_east.inst.cb_conf_bus[288] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11288_ (.D(\cb_east.inst.cb_conf_bus[289] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11289_ (.D(\cb_east.inst.cb_conf_bus[290] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11290_ (.D(\cb_east.inst.cb_conf_bus[291] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11291_ (.D(\cb_east.inst.cb_conf_bus[292] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11292_ (.D(\cb_east.inst.cb_conf_bus[293] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11293_ (.D(\cb_east.inst.cb_conf_bus[294] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[4].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11294_ (.D(\cb_east.inst.cb_conf_bus[295] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11295_ (.D(\cb_east.inst.cb_conf_bus[296] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11296_ (.D(\cb_east.inst.cb_conf_bus[297] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11297_ (.D(\cb_east.inst.cb_conf_bus[298] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11298_ (.D(\cb_east.inst.cb_conf_bus[299] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11299_ (.D(\cb_east.inst.cb_conf_bus[300] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11300_ (.D(\cb_east.inst.cb_conf_bus[301] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11301_ (.D(\cb_east.inst.cb_conf_bus[302] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11302_ (.D(\cb_east.inst.cb_conf_bus[303] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11303_ (.D(\cb_east.inst.cb_conf_bus[304] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11304_ (.D(\cb_east.inst.cb_conf_bus[305] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11305_ (.D(\cb_east.inst.cb_conf_bus[306] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11306_ (.D(\cb_east.inst.cb_conf_bus[307] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11307_ (.D(\cb_east.inst.cb_conf_bus[308] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11308_ (.D(\cb_east.inst.cb_conf_bus[309] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11309_ (.D(\cb_east.inst.cb_conf_bus[310] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11310_ (.D(\cb_east.inst.cb_conf_bus[311] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[5].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11311_ (.D(\cb_east.inst.cb_conf_bus[312] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11312_ (.D(\cb_east.inst.cb_conf_bus[313] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11313_ (.D(\cb_east.inst.cb_conf_bus[314] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11314_ (.D(\cb_east.inst.cb_conf_bus[315] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11315_ (.D(\cb_east.inst.cb_conf_bus[316] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11316_ (.D(\cb_east.inst.cb_conf_bus[317] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11317_ (.D(\cb_east.inst.cb_conf_bus[318] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11318_ (.D(\cb_east.inst.cb_conf_bus[319] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11319_ (.D(\cb_east.inst.cb_conf_bus[320] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11320_ (.D(\cb_east.inst.cb_conf_bus[321] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11321_ (.D(\cb_east.inst.cb_conf_bus[322] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11322_ (.D(\cb_east.inst.cb_conf_bus[323] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11323_ (.D(\cb_east.inst.cb_conf_bus[324] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11324_ (.D(\cb_east.inst.cb_conf_bus[325] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11325_ (.D(\cb_east.inst.cb_conf_bus[326] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11326_ (.D(\cb_east.inst.cb_conf_bus[327] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11327_ (.D(\cb_east.inst.cb_conf_bus[328] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[6].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11328_ (.D(\cb_east.inst.cb_conf_bus[329] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11329_ (.D(\cb_east.inst.cb_conf_bus[330] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11330_ (.D(\cb_east.inst.cb_conf_bus[331] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11331_ (.D(\cb_east.inst.cb_conf_bus[332] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11332_ (.D(\cb_east.inst.cb_conf_bus[333] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11333_ (.D(\cb_east.inst.cb_conf_bus[334] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11334_ (.D(\cb_east.inst.cb_conf_bus[335] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11335_ (.D(\cb_east.inst.cb_conf_bus[336] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11336_ (.D(\cb_east.inst.cb_conf_bus[337] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11337_ (.D(\cb_east.inst.cb_conf_bus[338] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11338_ (.D(\cb_east.inst.cb_conf_bus[339] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11339_ (.D(\cb_east.inst.cb_conf_bus[340] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11340_ (.D(\cb_east.inst.cb_conf_bus[341] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11341_ (.D(\cb_east.inst.cb_conf_bus[342] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11342_ (.D(\cb_east.inst.cb_conf_bus[343] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11343_ (.D(\cb_east.inst.cb_conf_bus[344] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11344_ (.D(\cb_east.inst.cb_conf_bus[345] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[7].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11345_ (.D(\cb_east.inst.cb_conf_bus[346] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11346_ (.D(\cb_east.inst.cb_conf_bus[347] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11347_ (.D(\cb_east.inst.cb_conf_bus[348] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11348_ (.D(\cb_east.inst.cb_conf_bus[349] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11349_ (.D(\cb_east.inst.cb_conf_bus[350] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11350_ (.D(\cb_east.inst.cb_conf_bus[351] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11351_ (.D(\cb_east.inst.cb_conf_bus[352] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11352_ (.D(\cb_east.inst.cb_conf_bus[353] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11353_ (.D(\cb_east.inst.cb_conf_bus[354] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11354_ (.D(\cb_east.inst.cb_conf_bus[355] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11355_ (.D(\cb_east.inst.cb_conf_bus[356] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11356_ (.D(\cb_east.inst.cb_conf_bus[357] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11357_ (.D(\cb_east.inst.cb_conf_bus[358] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11358_ (.D(\cb_east.inst.cb_conf_bus[359] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11359_ (.D(\cb_east.inst.cb_conf_bus[360] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11360_ (.D(\cb_east.inst.cb_conf_bus[361] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11361_ (.D(\cb_east.inst.cb_conf_bus[362] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[8].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11362_ (.D(\cb_east.inst.cb_conf_bus[363] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11363_ (.D(\cb_east.inst.cb_conf_bus[364] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11364_ (.D(\cb_east.inst.cb_conf_bus[365] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11365_ (.D(\cb_east.inst.cb_conf_bus[366] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11366_ (.D(\cb_east.inst.cb_conf_bus[367] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11367_ (.D(\cb_east.inst.cb_conf_bus[368] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11368_ (.D(\cb_east.inst.cb_conf_bus[369] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11369_ (.D(\cb_east.inst.cb_conf_bus[370] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11370_ (.D(\cb_east.inst.cb_conf_bus[371] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11371_ (.D(\cb_east.inst.cb_conf_bus[372] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[5].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11372_ (.D(\cb_east.inst.cb_conf_bus[373] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[6].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11373_ (.D(\cb_east.inst.cb_conf_bus[374] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].doubles[7].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11374_ (.D(\cb_east.inst.cb_conf_bus[375] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].directs[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11375_ (.D(\cb_east.inst.cb_conf_bus[376] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].directs[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11376_ (.D(\cb_east.inst.cb_conf_bus[377] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].directs[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11377_ (.D(\cb_east.inst.cb_conf_bus[378] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].directs[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11378_ (.D(\cb_east.inst.cb_conf_bus[379] ),
    .Q(\cb_east.inst.connectaroni.clb1_inputs[9].directs[4].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11379_ (.D(\cb_east.inst.cb_conf_bus[380] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11380_ (.D(\cb_east.inst.cb_conf_bus[381] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11381_ (.D(\cb_east.inst.cb_conf_bus[382] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11382_ (.D(\cb_east.inst.cb_conf_bus[383] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11383_ (.D(\cb_east.inst.cb_conf_bus[384] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11384_ (.D(\cb_east.inst.cb_conf_bus[385] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11385_ (.D(\cb_east.inst.cb_conf_bus[386] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11386_ (.D(\cb_east.inst.cb_conf_bus[387] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[0].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11387_ (.D(\cb_east.inst.cb_conf_bus[388] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11388_ (.D(\cb_east.inst.cb_conf_bus[389] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11389_ (.D(\cb_east.inst.cb_conf_bus[390] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11390_ (.D(\cb_east.inst.cb_conf_bus[391] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11391_ (.D(\cb_east.inst.cb_conf_bus[392] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11392_ (.D(\cb_east.inst.cb_conf_bus[393] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11393_ (.D(\cb_east.inst.cb_conf_bus[394] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11394_ (.D(\cb_east.inst.cb_conf_bus[395] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[1].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11395_ (.D(\cb_east.inst.cb_conf_bus[396] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11396_ (.D(\cb_east.inst.cb_conf_bus[397] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11397_ (.D(\cb_east.inst.cb_conf_bus[398] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11398_ (.D(\cb_east.inst.cb_conf_bus[399] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11399_ (.D(\cb_east.inst.cb_conf_bus[400] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11400_ (.D(\cb_east.inst.cb_conf_bus[401] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11401_ (.D(\cb_east.inst.cb_conf_bus[402] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11402_ (.D(\cb_east.inst.cb_conf_bus[403] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[2].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11403_ (.D(\cb_east.inst.cb_conf_bus[404] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11404_ (.D(\cb_east.inst.cb_conf_bus[405] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11405_ (.D(\cb_east.inst.cb_conf_bus[406] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11406_ (.D(\cb_east.inst.cb_conf_bus[407] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11407_ (.D(\cb_east.inst.cb_conf_bus[408] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11408_ (.D(\cb_east.inst.cb_conf_bus[409] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11409_ (.D(\cb_east.inst.cb_conf_bus[410] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11410_ (.D(\cb_east.inst.cb_conf_bus[411] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[3].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11411_ (.D(\cb_east.inst.cb_conf_bus[412] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].singles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11412_ (.D(\cb_east.inst.cb_conf_bus[413] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].singles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11413_ (.D(\cb_east.inst.cb_conf_bus[414] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].singles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11414_ (.D(\cb_east.inst.cb_conf_bus[415] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].singles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11415_ (.D(\cb_east.inst.cb_conf_bus[416] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[0].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11416_ (.D(\cb_east.inst.cb_conf_bus[417] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[1].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11417_ (.D(\cb_east.inst.cb_conf_bus[418] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[2].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__dlxtp_1 _11418_ (.D(\cb_east.inst.cb_conf_bus[419] ),
    .Q(\cb_east.inst.connectaroni.clb1_outputs[4].doubles[3].s.c ),
    .GATE(set_out_hard));
 sky130_fd_sc_hd__mux4_1 _11419_ (.A0(_04128_),
    .A1(_04135_),
    .A2(_04136_),
    .A3(_04137_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04120_));
 transmission_gate_cell _11420_ (.Cnot(_00057_),
    .C(_04124_),
    .A(_04120_),
    .B(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11421_ (.A0(_04138_),
    .A1(_04139_),
    .A2(_04140_),
    .A3(_04141_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04121_));
 transmission_gate_cell _11422_ (.Cnot(_00058_),
    .C(_04125_),
    .A(_04121_),
    .B(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11423_ (.A0(_04142_),
    .A1(_04143_),
    .A2(_04129_),
    .A3(_04130_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04122_));
 transmission_gate_cell _11424_ (.Cnot(_00059_),
    .C(_04126_),
    .A(_04122_),
    .B(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11425_ (.A0(_04131_),
    .A1(_04132_),
    .A2(_04133_),
    .A3(_04134_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04123_));
 transmission_gate_cell _11426_ (.Cnot(_00060_),
    .C(_04127_),
    .A(_04123_),
    .B(\cb_east.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11427_ (.A0(_04152_),
    .A1(_04159_),
    .A2(_04160_),
    .A3(_04161_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04144_));
 transmission_gate_cell _11428_ (.Cnot(_00061_),
    .C(_04148_),
    .A(_04144_),
    .B(\slice.sliceluroni.cc.P[0] ));
 sky130_fd_sc_hd__mux4_1 _11429_ (.A0(_04162_),
    .A1(_04163_),
    .A2(_04164_),
    .A3(_04165_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04145_));
 transmission_gate_cell _11430_ (.Cnot(_00062_),
    .C(_04149_),
    .A(_04145_),
    .B(\slice.sliceluroni.cc.P[0] ));
 sky130_fd_sc_hd__mux4_1 _11431_ (.A0(_04166_),
    .A1(_04167_),
    .A2(_04153_),
    .A3(_04154_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04146_));
 transmission_gate_cell _11432_ (.Cnot(_00063_),
    .C(_04150_),
    .A(_04146_),
    .B(\slice.sliceluroni.cc.P[0] ));
 sky130_fd_sc_hd__mux4_1 _11433_ (.A0(_04155_),
    .A1(_04156_),
    .A2(_04157_),
    .A3(_04158_),
    .S0(\cb_east.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_east.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04147_));
 transmission_gate_cell _11434_ (.Cnot(_00064_),
    .C(_04151_),
    .A(_04147_),
    .B(\slice.sliceluroni.cc.P[0] ));
 sky130_fd_sc_hd__mux4_1 _11435_ (.A0(_04177_),
    .A1(_04184_),
    .A2(_04185_),
    .A3(_04186_),
    .S0(clb_south_in[4]),
    .S1(clb_south_in[5]),
    .X(_04169_));
 transmission_gate_cell _11436_ (.Cnot(_00065_),
    .C(_04173_),
    .A(_04169_),
    .B(clb_south_out[1]));
 sky130_fd_sc_hd__mux4_1 _11437_ (.A0(_04187_),
    .A1(_04188_),
    .A2(_04189_),
    .A3(_04190_),
    .S0(clb_south_in[4]),
    .S1(clb_south_in[5]),
    .X(_04170_));
 transmission_gate_cell _11438_ (.Cnot(_00066_),
    .C(_04174_),
    .A(_04170_),
    .B(clb_south_out[1]));
 sky130_fd_sc_hd__mux4_1 _11439_ (.A0(_04191_),
    .A1(_04192_),
    .A2(_04178_),
    .A3(_04179_),
    .S0(clb_south_in[4]),
    .S1(clb_south_in[5]),
    .X(_04171_));
 transmission_gate_cell _11440_ (.Cnot(_00067_),
    .C(_04175_),
    .A(_04171_),
    .B(clb_south_out[1]));
 sky130_fd_sc_hd__mux4_1 _11441_ (.A0(_04180_),
    .A1(_04181_),
    .A2(_04182_),
    .A3(_04183_),
    .S0(clb_south_in[4]),
    .S1(clb_south_in[5]),
    .X(_04172_));
 transmission_gate_cell _11442_ (.Cnot(_00068_),
    .C(_04176_),
    .A(_04172_),
    .B(clb_south_out[1]));
 sky130_fd_sc_hd__mux4_1 _11443_ (.A0(_04201_),
    .A1(_04208_),
    .A2(_04209_),
    .A3(_04210_),
    .S0(clb_south_in[0]),
    .S1(clb_south_in[1]),
    .X(_04193_));
 transmission_gate_cell _11444_ (.Cnot(_00069_),
    .C(_04197_),
    .A(_04193_),
    .B(\slice.sliceluroni.cc.P[1] ));
 sky130_fd_sc_hd__mux4_1 _11445_ (.A0(_04211_),
    .A1(_04212_),
    .A2(_04213_),
    .A3(_04214_),
    .S0(clb_south_in[0]),
    .S1(clb_south_in[1]),
    .X(_04194_));
 transmission_gate_cell _11446_ (.Cnot(_00070_),
    .C(_04198_),
    .A(_04194_),
    .B(\slice.sliceluroni.cc.P[1] ));
 sky130_fd_sc_hd__mux4_1 _11447_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04202_),
    .A3(_04203_),
    .S0(clb_south_in[0]),
    .S1(clb_south_in[1]),
    .X(_04195_));
 transmission_gate_cell _11448_ (.Cnot(_00071_),
    .C(_04199_),
    .A(_04195_),
    .B(\slice.sliceluroni.cc.P[1] ));
 sky130_fd_sc_hd__mux4_1 _11449_ (.A0(_04204_),
    .A1(_04205_),
    .A2(_04206_),
    .A3(_04207_),
    .S0(clb_south_in[0]),
    .S1(clb_south_in[1]),
    .X(_04196_));
 transmission_gate_cell _11450_ (.Cnot(_00072_),
    .C(_04200_),
    .A(_04196_),
    .B(\slice.sliceluroni.cc.P[1] ));
 sky130_fd_sc_hd__mux4_1 _11451_ (.A0(_04226_),
    .A1(_04233_),
    .A2(_04234_),
    .A3(_04235_),
    .S0(clb_west_in[4]),
    .S1(clb_west_in[5]),
    .X(_04218_));
 transmission_gate_cell _11452_ (.Cnot(_00073_),
    .C(_04222_),
    .A(_04218_),
    .B(clb_west_out[1]));
 sky130_fd_sc_hd__mux4_1 _11453_ (.A0(_04236_),
    .A1(_04237_),
    .A2(_04238_),
    .A3(_04239_),
    .S0(clb_west_in[4]),
    .S1(clb_west_in[5]),
    .X(_04219_));
 transmission_gate_cell _11454_ (.Cnot(_00074_),
    .C(_04223_),
    .A(_04219_),
    .B(clb_west_out[1]));
 sky130_fd_sc_hd__mux4_1 _11455_ (.A0(_04240_),
    .A1(_04241_),
    .A2(_04227_),
    .A3(_04228_),
    .S0(clb_west_in[4]),
    .S1(clb_west_in[5]),
    .X(_04220_));
 transmission_gate_cell _11456_ (.Cnot(_00075_),
    .C(_04224_),
    .A(_04220_),
    .B(clb_west_out[1]));
 sky130_fd_sc_hd__mux4_1 _11457_ (.A0(_04229_),
    .A1(_04230_),
    .A2(_04231_),
    .A3(_04232_),
    .S0(clb_west_in[4]),
    .S1(clb_west_in[5]),
    .X(_04221_));
 transmission_gate_cell _11458_ (.Cnot(_00076_),
    .C(_04225_),
    .A(_04221_),
    .B(clb_west_out[1]));
 sky130_fd_sc_hd__mux4_1 _11459_ (.A0(_04250_),
    .A1(_04257_),
    .A2(_04258_),
    .A3(_04259_),
    .S0(clb_west_in[0]),
    .S1(clb_west_in[1]),
    .X(_04242_));
 transmission_gate_cell _11460_ (.Cnot(_00077_),
    .C(_04246_),
    .A(_04242_),
    .B(\slice.sliceluroni.cc.P[2] ));
 sky130_fd_sc_hd__mux4_1 _11461_ (.A0(_04260_),
    .A1(_04261_),
    .A2(_04262_),
    .A3(_04263_),
    .S0(clb_west_in[0]),
    .S1(clb_west_in[1]),
    .X(_04243_));
 transmission_gate_cell _11462_ (.Cnot(_00078_),
    .C(_04247_),
    .A(_04243_),
    .B(\slice.sliceluroni.cc.P[2] ));
 sky130_fd_sc_hd__mux4_1 _11463_ (.A0(_04264_),
    .A1(_04265_),
    .A2(_04251_),
    .A3(_04252_),
    .S0(clb_west_in[0]),
    .S1(clb_west_in[1]),
    .X(_04244_));
 transmission_gate_cell _11464_ (.Cnot(_00079_),
    .C(_04248_),
    .A(_04244_),
    .B(\slice.sliceluroni.cc.P[2] ));
 sky130_fd_sc_hd__mux4_1 _11465_ (.A0(_04253_),
    .A1(_04254_),
    .A2(_04255_),
    .A3(_04256_),
    .S0(clb_west_in[0]),
    .S1(clb_west_in[1]),
    .X(_04245_));
 transmission_gate_cell _11466_ (.Cnot(_00080_),
    .C(_04249_),
    .A(_04245_),
    .B(\slice.sliceluroni.cc.P[2] ));
 sky130_fd_sc_hd__mux4_1 _11467_ (.A0(_04275_),
    .A1(_04282_),
    .A2(_04283_),
    .A3(_04284_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04267_));
 transmission_gate_cell _11468_ (.Cnot(_00081_),
    .C(_04271_),
    .A(_04267_),
    .B(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11469_ (.A0(_04285_),
    .A1(_04286_),
    .A2(_04287_),
    .A3(_04288_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04268_));
 transmission_gate_cell _11470_ (.Cnot(_00082_),
    .C(_04272_),
    .A(_04268_),
    .B(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11471_ (.A0(_04289_),
    .A1(_04290_),
    .A2(_04276_),
    .A3(_04277_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04269_));
 transmission_gate_cell _11472_ (.Cnot(_00083_),
    .C(_04273_),
    .A(_04269_),
    .B(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11473_ (.A0(_04278_),
    .A1(_04279_),
    .A2(_04280_),
    .A3(_04281_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[4].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[5].directs[0].s.a ),
    .X(_04270_));
 transmission_gate_cell _11474_ (.Cnot(_00084_),
    .C(_04274_),
    .A(_04270_),
    .B(\cb_north.inst.connectaroni.clb0_outputs[1].doubles[0].s.b ));
 sky130_fd_sc_hd__mux4_1 _11475_ (.A0(_04299_),
    .A1(_04306_),
    .A2(_04307_),
    .A3(_04308_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04291_));
 transmission_gate_cell _11476_ (.Cnot(_00085_),
    .C(_04295_),
    .A(_04291_),
    .B(\slice.sliceluroni.cc.P[3] ));
 sky130_fd_sc_hd__mux4_1 _11477_ (.A0(_04309_),
    .A1(_04310_),
    .A2(_04311_),
    .A3(_04312_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04292_));
 transmission_gate_cell _11478_ (.Cnot(_00086_),
    .C(_04296_),
    .A(_04292_),
    .B(\slice.sliceluroni.cc.P[3] ));
 sky130_fd_sc_hd__mux4_1 _11479_ (.A0(_04313_),
    .A1(_04314_),
    .A2(_04300_),
    .A3(_04301_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04293_));
 transmission_gate_cell _11480_ (.Cnot(_00087_),
    .C(_04297_),
    .A(_04293_),
    .B(\slice.sliceluroni.cc.P[3] ));
 sky130_fd_sc_hd__mux4_1 _11481_ (.A0(_04302_),
    .A1(_04303_),
    .A2(_04304_),
    .A3(_04305_),
    .S0(\cb_north.inst.connectaroni.clb0_inputs[0].directs[0].s.a ),
    .S1(\cb_north.inst.connectaroni.clb0_inputs[1].directs[0].s.a ),
    .X(_04294_));
 transmission_gate_cell _11482_ (.Cnot(_00088_),
    .C(_04298_),
    .A(_04294_),
    .B(\slice.sliceluroni.cc.P[3] ));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.e0s1.impl  (.Cnot(_00001_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e0s1.c ),
    .A(south_double[5]),
    .B(east_double[4]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.e1s0.impl  (.Cnot(_00002_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1s0.c ),
    .A(south_double[4]),
    .B(east_double[5]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.e1w1.impl  (.Cnot(_00003_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.e1w1.c ),
    .A(west_double[1]),
    .B(east_double[5]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.n0e0.impl  (.Cnot(_00004_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0e0.c ),
    .A(east_double[4]),
    .B(north_double[0]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.n0s0.impl  (.Cnot(_00005_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n0s0.c ),
    .A(south_double[4]),
    .B(north_double[0]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.n1e1.impl  (.Cnot(_00006_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.n1e1.c ),
    .A(east_double[5]),
    .B(north_double[1]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.s0w0.impl  (.Cnot(_00007_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s0w0.c ),
    .A(west_double[0]),
    .B(south_double[4]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.s1n1.impl  (.Cnot(_00008_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1n1.c ),
    .A(north_double[1]),
    .B(south_double[5]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.s1w1.impl  (.Cnot(_00009_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.s1w1.c ),
    .A(west_double[1]),
    .B(south_double[5]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.w0e0.impl  (.Cnot(_00010_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0e0.c ),
    .A(east_double[4]),
    .B(west_double[0]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.w0n1.impl  (.Cnot(_00011_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w0n1.c ),
    .A(north_double[1]),
    .B(west_double[0]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[0].elem.w1n0.impl  (.Cnot(_00012_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[0].elem.w1n0.c ),
    .A(north_double[0]),
    .B(west_double[1]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.e0s1.impl  (.Cnot(_00013_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e0s1.c ),
    .A(south_double[7]),
    .B(east_double[6]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.e1s0.impl  (.Cnot(_00014_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1s0.c ),
    .A(south_double[6]),
    .B(east_double[7]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.e1w1.impl  (.Cnot(_00015_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.e1w1.c ),
    .A(west_double[3]),
    .B(east_double[7]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.n0e0.impl  (.Cnot(_00016_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0e0.c ),
    .A(east_double[6]),
    .B(north_double[2]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.n0s0.impl  (.Cnot(_00017_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n0s0.c ),
    .A(south_double[6]),
    .B(north_double[2]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.n1e1.impl  (.Cnot(_00018_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.n1e1.c ),
    .A(east_double[7]),
    .B(north_double[3]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.s0w0.impl  (.Cnot(_00019_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s0w0.c ),
    .A(west_double[2]),
    .B(south_double[6]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.s1n1.impl  (.Cnot(_00020_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1n1.c ),
    .A(north_double[3]),
    .B(south_double[7]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.s1w1.impl  (.Cnot(_00021_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.s1w1.c ),
    .A(west_double[3]),
    .B(south_double[7]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.w0e0.impl  (.Cnot(_00022_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0e0.c ),
    .A(east_double[6]),
    .B(west_double[2]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.w0n1.impl  (.Cnot(_00023_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w0n1.c ),
    .A(north_double[3]),
    .B(west_double[2]));
 transmission_gate_cell \sb.switcharoni.dusb.switch_box_element_two[1].elem.w1n0.impl  (.Cnot(_00024_),
    .C(\sb.switcharoni.dusb.switch_box_element_two[1].elem.w1n0.c ),
    .A(north_double[2]),
    .B(west_double[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.e0s1.impl  (.Cnot(_00025_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.e0s1.c ),
    .A(south_single[1]),
    .B(east_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.e1s0.impl  (.Cnot(_00026_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1s0.c ),
    .A(south_single[0]),
    .B(east_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.e1w1.impl  (.Cnot(_00027_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.e1w1.c ),
    .A(west_single[1]),
    .B(east_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.n0e0.impl  (.Cnot(_00028_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0e0.c ),
    .A(east_single[0]),
    .B(north_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.n0s0.impl  (.Cnot(_00029_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.n0s0.c ),
    .A(south_single[0]),
    .B(north_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.n1e1.impl  (.Cnot(_00030_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.n1e1.c ),
    .A(east_single[1]),
    .B(north_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.s0w0.impl  (.Cnot(_00031_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.s0w0.c ),
    .A(west_single[0]),
    .B(south_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.s1n1.impl  (.Cnot(_00032_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1n1.c ),
    .A(north_single[1]),
    .B(south_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.s1w1.impl  (.Cnot(_00033_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.s1w1.c ),
    .A(west_single[1]),
    .B(south_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.w0e0.impl  (.Cnot(_00034_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0e0.c ),
    .A(east_single[0]),
    .B(west_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.w0n1.impl  (.Cnot(_00035_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.w0n1.c ),
    .A(north_single[1]),
    .B(west_single[0]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[0].elem.w1n0.impl  (.Cnot(_00036_),
    .C(\sb.switcharoni.susb.switch_box_element_two[0].elem.w1n0.c ),
    .A(north_single[0]),
    .B(west_single[1]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.e0s1.impl  (.Cnot(_00037_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.e0s1.c ),
    .A(south_single[3]),
    .B(east_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.e1s0.impl  (.Cnot(_00038_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1s0.c ),
    .A(south_single[2]),
    .B(east_single[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.e1w1.impl  (.Cnot(_00039_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.e1w1.c ),
    .A(west_single[3]),
    .B(east_single[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.n0e0.impl  (.Cnot(_00040_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0e0.c ),
    .A(east_single[2]),
    .B(north_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.n0s0.impl  (.Cnot(_00041_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.n0s0.c ),
    .A(south_single[2]),
    .B(north_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.n1e1.impl  (.Cnot(_00042_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.n1e1.c ),
    .A(east_single[3]),
    .B(north_single[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.s0w0.impl  (.Cnot(_00043_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.s0w0.c ),
    .A(west_single[2]),
    .B(south_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.s1n1.impl  (.Cnot(_00044_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1n1.c ),
    .A(north_single[3]),
    .B(south_single[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.s1w1.impl  (.Cnot(_00045_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.s1w1.c ),
    .A(west_single[3]),
    .B(south_single[3]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.w0e0.impl  (.Cnot(_00046_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0e0.c ),
    .A(east_single[2]),
    .B(west_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.w0n1.impl  (.Cnot(_00047_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.w0n1.c ),
    .A(north_single[3]),
    .B(west_single[2]));
 transmission_gate_cell \sb.switcharoni.susb.switch_box_element_two[1].elem.w1n0.impl  (.Cnot(_00048_),
    .C(\sb.switcharoni.susb.switch_box_element_two[1].elem.w1n0.c ),
    .A(north_single[2]),
    .B(west_single[3]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_0 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_0));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_1 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_1));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_2 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_2));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_3 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_3));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_4 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_4));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_5 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_5));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_6 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_6));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_7 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_7));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_8 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_8));
 sky130_fd_sc_hd__buf_8 psn_inst_psn_buff_9 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_9));
 sky130_fd_sc_hd__buf_8 psn_inst_psn_buff_10 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_10));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_11 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_11));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_12 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_12));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_13 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_13));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_14 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_14));
 sky130_fd_sc_hd__buf_8 psn_inst_psn_buff_15 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_15));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_16 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_16));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_17 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_17));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_18 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_18));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_19 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_19));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_20 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_20));
 sky130_fd_sc_hd__buf_4 psn_inst_psn_buff_21 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_21));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_22 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_22));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_23 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_23));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_24 (.A(\cb_east.inst.configuroni.comb_shifter.head_bit.shift_enable ),
    .X(psn_net_24));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_0_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_1_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_2_0_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_3_0_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_4_0_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_5_0_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_6_0_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_7_0_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_8_0_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_9_0_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_10_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_11_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_12_0_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_13_0_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_14_0_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_15_0_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_16_0_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_17_0_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_18_0_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_19_0_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_20_0_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_21_0_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_22_0_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_23_0_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_24_0_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_25_0_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_26_0_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_27_0_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_28_0_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_29_0_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_30_0_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_31_0_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_32_0_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_33_0_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_34_0_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_35_0_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_36_0_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_37_0_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_38_0_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_39_0_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_40_0_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_41_0_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_42_0_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_43_0_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_44_0_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_45_0_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_46_0_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_47_0_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_48_0_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_49_0_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_50_0_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_51_0_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_52_0_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_53_0_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_54_0_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_55_0_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_56_0_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_57_0_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_58_0_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_59_0_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_60_0_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_61_0_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_62_0_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_63_0_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_0_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_7_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_1_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_7_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_2_0_clk (.A(clknet_6_1_0_clk),
    .X(clknet_7_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_3_0_clk (.A(clknet_6_1_0_clk),
    .X(clknet_7_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_4_0_clk (.A(clknet_6_2_0_clk),
    .X(clknet_7_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_5_0_clk (.A(clknet_6_2_0_clk),
    .X(clknet_7_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_6_0_clk (.A(clknet_6_3_0_clk),
    .X(clknet_7_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_7_0_clk (.A(clknet_6_3_0_clk),
    .X(clknet_7_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_8_0_clk (.A(clknet_6_4_0_clk),
    .X(clknet_7_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_9_0_clk (.A(clknet_6_4_0_clk),
    .X(clknet_7_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_10_0_clk (.A(clknet_6_5_0_clk),
    .X(clknet_7_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_11_0_clk (.A(clknet_6_5_0_clk),
    .X(clknet_7_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_12_0_clk (.A(clknet_6_6_0_clk),
    .X(clknet_7_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_13_0_clk (.A(clknet_6_6_0_clk),
    .X(clknet_7_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_14_0_clk (.A(clknet_6_7_0_clk),
    .X(clknet_7_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_15_0_clk (.A(clknet_6_7_0_clk),
    .X(clknet_7_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_16_0_clk (.A(clknet_6_8_0_clk),
    .X(clknet_7_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_17_0_clk (.A(clknet_6_8_0_clk),
    .X(clknet_7_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_18_0_clk (.A(clknet_6_9_0_clk),
    .X(clknet_7_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_19_0_clk (.A(clknet_6_9_0_clk),
    .X(clknet_7_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_20_0_clk (.A(clknet_6_10_0_clk),
    .X(clknet_7_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_21_0_clk (.A(clknet_6_10_0_clk),
    .X(clknet_7_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_22_0_clk (.A(clknet_6_11_0_clk),
    .X(clknet_7_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_23_0_clk (.A(clknet_6_11_0_clk),
    .X(clknet_7_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_24_0_clk (.A(clknet_6_12_0_clk),
    .X(clknet_7_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_25_0_clk (.A(clknet_6_12_0_clk),
    .X(clknet_7_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_26_0_clk (.A(clknet_6_13_0_clk),
    .X(clknet_7_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_27_0_clk (.A(clknet_6_13_0_clk),
    .X(clknet_7_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_28_0_clk (.A(clknet_6_14_0_clk),
    .X(clknet_7_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_29_0_clk (.A(clknet_6_14_0_clk),
    .X(clknet_7_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_30_0_clk (.A(clknet_6_15_0_clk),
    .X(clknet_7_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_31_0_clk (.A(clknet_6_15_0_clk),
    .X(clknet_7_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_32_0_clk (.A(clknet_6_16_0_clk),
    .X(clknet_7_32_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_33_0_clk (.A(clknet_6_16_0_clk),
    .X(clknet_7_33_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_34_0_clk (.A(clknet_6_17_0_clk),
    .X(clknet_7_34_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_35_0_clk (.A(clknet_6_17_0_clk),
    .X(clknet_7_35_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_36_0_clk (.A(clknet_6_18_0_clk),
    .X(clknet_7_36_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_37_0_clk (.A(clknet_6_18_0_clk),
    .X(clknet_7_37_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_38_0_clk (.A(clknet_6_19_0_clk),
    .X(clknet_7_38_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_39_0_clk (.A(clknet_6_19_0_clk),
    .X(clknet_7_39_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_40_0_clk (.A(clknet_6_20_0_clk),
    .X(clknet_7_40_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_41_0_clk (.A(clknet_6_20_0_clk),
    .X(clknet_7_41_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_42_0_clk (.A(clknet_6_21_0_clk),
    .X(clknet_7_42_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_43_0_clk (.A(clknet_6_21_0_clk),
    .X(clknet_7_43_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_44_0_clk (.A(clknet_6_22_0_clk),
    .X(clknet_7_44_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_45_0_clk (.A(clknet_6_22_0_clk),
    .X(clknet_7_45_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_46_0_clk (.A(clknet_6_23_0_clk),
    .X(clknet_7_46_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_47_0_clk (.A(clknet_6_23_0_clk),
    .X(clknet_7_47_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_48_0_clk (.A(clknet_6_24_0_clk),
    .X(clknet_7_48_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_49_0_clk (.A(clknet_6_24_0_clk),
    .X(clknet_7_49_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_50_0_clk (.A(clknet_6_25_0_clk),
    .X(clknet_7_50_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_51_0_clk (.A(clknet_6_25_0_clk),
    .X(clknet_7_51_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_52_0_clk (.A(clknet_6_26_0_clk),
    .X(clknet_7_52_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_53_0_clk (.A(clknet_6_26_0_clk),
    .X(clknet_7_53_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_54_0_clk (.A(clknet_6_27_0_clk),
    .X(clknet_7_54_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_55_0_clk (.A(clknet_6_27_0_clk),
    .X(clknet_7_55_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_56_0_clk (.A(clknet_6_28_0_clk),
    .X(clknet_7_56_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_57_0_clk (.A(clknet_6_28_0_clk),
    .X(clknet_7_57_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_58_0_clk (.A(clknet_6_29_0_clk),
    .X(clknet_7_58_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_59_0_clk (.A(clknet_6_29_0_clk),
    .X(clknet_7_59_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_60_0_clk (.A(clknet_6_30_0_clk),
    .X(clknet_7_60_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_61_0_clk (.A(clknet_6_30_0_clk),
    .X(clknet_7_61_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_62_0_clk (.A(clknet_6_31_0_clk),
    .X(clknet_7_62_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_63_0_clk (.A(clknet_6_31_0_clk),
    .X(clknet_7_63_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_64_0_clk (.A(clknet_6_32_0_clk),
    .X(clknet_7_64_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_65_0_clk (.A(clknet_6_32_0_clk),
    .X(clknet_7_65_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_66_0_clk (.A(clknet_6_33_0_clk),
    .X(clknet_7_66_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_67_0_clk (.A(clknet_6_33_0_clk),
    .X(clknet_7_67_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_68_0_clk (.A(clknet_6_34_0_clk),
    .X(clknet_7_68_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_69_0_clk (.A(clknet_6_34_0_clk),
    .X(clknet_7_69_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_70_0_clk (.A(clknet_6_35_0_clk),
    .X(clknet_7_70_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_71_0_clk (.A(clknet_6_35_0_clk),
    .X(clknet_7_71_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_72_0_clk (.A(clknet_6_36_0_clk),
    .X(clknet_7_72_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_73_0_clk (.A(clknet_6_36_0_clk),
    .X(clknet_7_73_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_74_0_clk (.A(clknet_6_37_0_clk),
    .X(clknet_7_74_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_75_0_clk (.A(clknet_6_37_0_clk),
    .X(clknet_7_75_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_76_0_clk (.A(clknet_6_38_0_clk),
    .X(clknet_7_76_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_77_0_clk (.A(clknet_6_38_0_clk),
    .X(clknet_7_77_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_78_0_clk (.A(clknet_6_39_0_clk),
    .X(clknet_7_78_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_79_0_clk (.A(clknet_6_39_0_clk),
    .X(clknet_7_79_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_80_0_clk (.A(clknet_6_40_0_clk),
    .X(clknet_7_80_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_81_0_clk (.A(clknet_6_40_0_clk),
    .X(clknet_7_81_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_82_0_clk (.A(clknet_6_41_0_clk),
    .X(clknet_7_82_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_83_0_clk (.A(clknet_6_41_0_clk),
    .X(clknet_7_83_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_84_0_clk (.A(clknet_6_42_0_clk),
    .X(clknet_7_84_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_85_0_clk (.A(clknet_6_42_0_clk),
    .X(clknet_7_85_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_86_0_clk (.A(clknet_6_43_0_clk),
    .X(clknet_7_86_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_87_0_clk (.A(clknet_6_43_0_clk),
    .X(clknet_7_87_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_88_0_clk (.A(clknet_6_44_0_clk),
    .X(clknet_7_88_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_89_0_clk (.A(clknet_6_44_0_clk),
    .X(clknet_7_89_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_90_0_clk (.A(clknet_6_45_0_clk),
    .X(clknet_7_90_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_91_0_clk (.A(clknet_6_45_0_clk),
    .X(clknet_7_91_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_92_0_clk (.A(clknet_6_46_0_clk),
    .X(clknet_7_92_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_93_0_clk (.A(clknet_6_46_0_clk),
    .X(clknet_7_93_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_94_0_clk (.A(clknet_6_47_0_clk),
    .X(clknet_7_94_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_95_0_clk (.A(clknet_6_47_0_clk),
    .X(clknet_7_95_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_96_0_clk (.A(clknet_6_48_0_clk),
    .X(clknet_7_96_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_97_0_clk (.A(clknet_6_48_0_clk),
    .X(clknet_7_97_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_98_0_clk (.A(clknet_6_49_0_clk),
    .X(clknet_7_98_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_99_0_clk (.A(clknet_6_49_0_clk),
    .X(clknet_7_99_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_100_0_clk (.A(clknet_6_50_0_clk),
    .X(clknet_7_100_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_101_0_clk (.A(clknet_6_50_0_clk),
    .X(clknet_7_101_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_102_0_clk (.A(clknet_6_51_0_clk),
    .X(clknet_7_102_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_103_0_clk (.A(clknet_6_51_0_clk),
    .X(clknet_7_103_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_104_0_clk (.A(clknet_6_52_0_clk),
    .X(clknet_7_104_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_105_0_clk (.A(clknet_6_52_0_clk),
    .X(clknet_7_105_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_106_0_clk (.A(clknet_6_53_0_clk),
    .X(clknet_7_106_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_107_0_clk (.A(clknet_6_53_0_clk),
    .X(clknet_7_107_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_108_0_clk (.A(clknet_6_54_0_clk),
    .X(clknet_7_108_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_109_0_clk (.A(clknet_6_54_0_clk),
    .X(clknet_7_109_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_110_0_clk (.A(clknet_6_55_0_clk),
    .X(clknet_7_110_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_111_0_clk (.A(clknet_6_55_0_clk),
    .X(clknet_7_111_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_112_0_clk (.A(clknet_6_56_0_clk),
    .X(clknet_7_112_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_113_0_clk (.A(clknet_6_56_0_clk),
    .X(clknet_7_113_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_114_0_clk (.A(clknet_6_57_0_clk),
    .X(clknet_7_114_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_115_0_clk (.A(clknet_6_57_0_clk),
    .X(clknet_7_115_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_116_0_clk (.A(clknet_6_58_0_clk),
    .X(clknet_7_116_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_117_0_clk (.A(clknet_6_58_0_clk),
    .X(clknet_7_117_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_118_0_clk (.A(clknet_6_59_0_clk),
    .X(clknet_7_118_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_119_0_clk (.A(clknet_6_59_0_clk),
    .X(clknet_7_119_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_120_0_clk (.A(clknet_6_60_0_clk),
    .X(clknet_7_120_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_121_0_clk (.A(clknet_6_60_0_clk),
    .X(clknet_7_121_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_122_0_clk (.A(clknet_6_61_0_clk),
    .X(clknet_7_122_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_123_0_clk (.A(clknet_6_61_0_clk),
    .X(clknet_7_123_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_124_0_clk (.A(clknet_6_62_0_clk),
    .X(clknet_7_124_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_125_0_clk (.A(clknet_6_62_0_clk),
    .X(clknet_7_125_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_126_0_clk (.A(clknet_6_63_0_clk),
    .X(clknet_7_126_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_127_0_clk (.A(clknet_6_63_0_clk),
    .X(clknet_7_127_0_clk));
endmodule
