VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_slicel
  CLASS BLOCK ;
  FOREIGN baked_slicel ;
  ORIGIN 0.000 0.000 ;
  SIZE 191.080 BY 201.800 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 182.280 191.080 182.880 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END carry_out
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 197.800 172.870 201.800 ;
    END
  END clk
  PIN comb_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 187.080 131.960 191.080 132.560 ;
    END
  END comb_output[0]
  PIN comb_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 187.080 144.880 191.080 145.480 ;
    END
  END comb_output[1]
  PIN comb_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END comb_output[2]
  PIN comb_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END comb_output[3]
  PIN comb_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END comb_output[4]
  PIN comb_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END comb_output[5]
  PIN comb_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 197.800 101.110 201.800 ;
    END
  END comb_output[6]
  PIN comb_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 197.800 113.070 201.800 ;
    END
  END comb_output[7]
  PIN higher_order_address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 6.160 191.080 6.760 ;
    END
  END higher_order_address[0]
  PIN higher_order_address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 18.400 191.080 19.000 ;
    END
  END higher_order_address[1]
  PIN luts_input[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 31.320 191.080 31.920 ;
    END
  END luts_input[0]
  PIN luts_input[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END luts_input[10]
  PIN luts_input[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END luts_input[11]
  PIN luts_input[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END luts_input[12]
  PIN luts_input[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END luts_input[13]
  PIN luts_input[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END luts_input[14]
  PIN luts_input[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END luts_input[15]
  PIN luts_input[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END luts_input[16]
  PIN luts_input[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END luts_input[17]
  PIN luts_input[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END luts_input[18]
  PIN luts_input[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END luts_input[19]
  PIN luts_input[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 43.560 191.080 44.160 ;
    END
  END luts_input[1]
  PIN luts_input[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END luts_input[20]
  PIN luts_input[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END luts_input[21]
  PIN luts_input[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END luts_input[22]
  PIN luts_input[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END luts_input[23]
  PIN luts_input[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 197.800 5.890 201.800 ;
    END
  END luts_input[24]
  PIN luts_input[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 197.800 17.390 201.800 ;
    END
  END luts_input[25]
  PIN luts_input[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 197.800 29.350 201.800 ;
    END
  END luts_input[26]
  PIN luts_input[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 197.800 41.310 201.800 ;
    END
  END luts_input[27]
  PIN luts_input[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 197.800 53.270 201.800 ;
    END
  END luts_input[28]
  PIN luts_input[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 197.800 65.230 201.800 ;
    END
  END luts_input[29]
  PIN luts_input[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 56.480 191.080 57.080 ;
    END
  END luts_input[2]
  PIN luts_input[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 197.800 77.190 201.800 ;
    END
  END luts_input[30]
  PIN luts_input[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 197.800 89.150 201.800 ;
    END
  END luts_input[31]
  PIN luts_input[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 68.720 191.080 69.320 ;
    END
  END luts_input[3]
  PIN luts_input[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 81.640 191.080 82.240 ;
    END
  END luts_input[4]
  PIN luts_input[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 93.880 191.080 94.480 ;
    END
  END luts_input[5]
  PIN luts_input[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 106.800 191.080 107.400 ;
    END
  END luts_input[6]
  PIN luts_input[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 119.720 191.080 120.320 ;
    END
  END luts_input[7]
  PIN luts_input[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END luts_input[8]
  PIN luts_input[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END luts_input[9]
  PIN reg_we
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.550 197.800 184.830 201.800 ;
    END
  END reg_we
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 187.080 195.200 191.080 195.800 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END set_in
  PIN set_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END set_in_soft
  PIN set_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.630 197.800 160.910 201.800 ;
    END
  END set_out
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END shift_in
  PIN shift_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END shift_in_soft
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.670 197.800 148.950 201.800 ;
    END
  END shift_out
  PIN sync_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 187.080 157.120 191.080 157.720 ;
    END
  END sync_output[0]
  PIN sync_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 187.080 170.040 191.080 170.640 ;
    END
  END sync_output[1]
  PIN sync_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END sync_output[2]
  PIN sync_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END sync_output[3]
  PIN sync_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END sync_output[4]
  PIN sync_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END sync_output[5]
  PIN sync_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 197.800 125.030 201.800 ;
    END
  END sync_output[6]
  PIN sync_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.710 197.800 136.990 201.800 ;
    END
  END sync_output[7]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 190.640 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 190.640 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 185.380 190.485 ;
      LAYER met1 ;
        RECT 5.520 10.640 185.380 193.420 ;
      LAYER met2 ;
        RECT 6.170 197.520 16.830 197.800 ;
        RECT 17.670 197.520 28.790 197.800 ;
        RECT 29.630 197.520 40.750 197.800 ;
        RECT 41.590 197.520 52.710 197.800 ;
        RECT 53.550 197.520 64.670 197.800 ;
        RECT 65.510 197.520 76.630 197.800 ;
        RECT 77.470 197.520 88.590 197.800 ;
        RECT 89.430 197.520 100.550 197.800 ;
        RECT 101.390 197.520 112.510 197.800 ;
        RECT 113.350 197.520 124.470 197.800 ;
        RECT 125.310 197.520 136.430 197.800 ;
        RECT 137.270 197.520 148.390 197.800 ;
        RECT 149.230 197.520 160.350 197.800 ;
        RECT 161.190 197.520 172.310 197.800 ;
        RECT 173.150 197.520 184.270 197.800 ;
        RECT 5.620 4.280 184.820 197.520 ;
        RECT 6.170 4.000 16.830 4.280 ;
        RECT 17.670 4.000 28.790 4.280 ;
        RECT 29.630 4.000 40.750 4.280 ;
        RECT 41.590 4.000 52.710 4.280 ;
        RECT 53.550 4.000 64.670 4.280 ;
        RECT 65.510 4.000 76.630 4.280 ;
        RECT 77.470 4.000 88.590 4.280 ;
        RECT 89.430 4.000 100.550 4.280 ;
        RECT 101.390 4.000 112.510 4.280 ;
        RECT 113.350 4.000 124.470 4.280 ;
        RECT 125.310 4.000 136.430 4.280 ;
        RECT 137.270 4.000 148.390 4.280 ;
        RECT 149.230 4.000 160.350 4.280 ;
        RECT 161.190 4.000 172.310 4.280 ;
        RECT 173.150 4.000 184.270 4.280 ;
      LAYER met3 ;
        RECT 4.000 194.840 186.680 195.665 ;
        RECT 4.400 194.800 186.680 194.840 ;
        RECT 4.400 193.440 187.080 194.800 ;
        RECT 4.000 183.280 187.080 193.440 ;
        RECT 4.000 181.880 186.680 183.280 ;
        RECT 4.000 180.560 187.080 181.880 ;
        RECT 4.400 179.160 187.080 180.560 ;
        RECT 4.000 171.040 187.080 179.160 ;
        RECT 4.000 169.640 186.680 171.040 ;
        RECT 4.000 166.280 187.080 169.640 ;
        RECT 4.400 164.880 187.080 166.280 ;
        RECT 4.000 158.120 187.080 164.880 ;
        RECT 4.000 156.720 186.680 158.120 ;
        RECT 4.000 152.000 187.080 156.720 ;
        RECT 4.400 150.600 187.080 152.000 ;
        RECT 4.000 145.880 187.080 150.600 ;
        RECT 4.000 144.480 186.680 145.880 ;
        RECT 4.000 137.040 187.080 144.480 ;
        RECT 4.400 135.640 187.080 137.040 ;
        RECT 4.000 132.960 187.080 135.640 ;
        RECT 4.000 131.560 186.680 132.960 ;
        RECT 4.000 122.760 187.080 131.560 ;
        RECT 4.400 121.360 187.080 122.760 ;
        RECT 4.000 120.720 187.080 121.360 ;
        RECT 4.000 119.320 186.680 120.720 ;
        RECT 4.000 108.480 187.080 119.320 ;
        RECT 4.400 107.800 187.080 108.480 ;
        RECT 4.400 107.080 186.680 107.800 ;
        RECT 4.000 106.400 186.680 107.080 ;
        RECT 4.000 94.880 187.080 106.400 ;
        RECT 4.000 94.200 186.680 94.880 ;
        RECT 4.400 93.480 186.680 94.200 ;
        RECT 4.400 92.800 187.080 93.480 ;
        RECT 4.000 82.640 187.080 92.800 ;
        RECT 4.000 81.240 186.680 82.640 ;
        RECT 4.000 79.920 187.080 81.240 ;
        RECT 4.400 78.520 187.080 79.920 ;
        RECT 4.000 69.720 187.080 78.520 ;
        RECT 4.000 68.320 186.680 69.720 ;
        RECT 4.000 64.960 187.080 68.320 ;
        RECT 4.400 63.560 187.080 64.960 ;
        RECT 4.000 57.480 187.080 63.560 ;
        RECT 4.000 56.080 186.680 57.480 ;
        RECT 4.000 50.680 187.080 56.080 ;
        RECT 4.400 49.280 187.080 50.680 ;
        RECT 4.000 44.560 187.080 49.280 ;
        RECT 4.000 43.160 186.680 44.560 ;
        RECT 4.000 36.400 187.080 43.160 ;
        RECT 4.400 35.000 187.080 36.400 ;
        RECT 4.000 32.320 187.080 35.000 ;
        RECT 4.000 30.920 186.680 32.320 ;
        RECT 4.000 22.120 187.080 30.920 ;
        RECT 4.400 20.720 187.080 22.120 ;
        RECT 4.000 19.400 187.080 20.720 ;
        RECT 4.000 18.000 186.680 19.400 ;
        RECT 4.000 7.840 187.080 18.000 ;
        RECT 4.400 7.160 187.080 7.840 ;
        RECT 4.400 6.440 186.680 7.160 ;
        RECT 4.000 5.760 186.680 6.440 ;
        RECT 4.000 4.255 187.080 5.760 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 190.640 ;
  END
END baked_slicel
END LIBRARY

