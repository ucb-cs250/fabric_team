VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_slicel
  CLASS BLOCK ;
  FOREIGN baked_slicel ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.615 BY 234.335 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.750 230.335 217.030 234.335 ;
    END
  END carry_out
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 8.880 223.615 9.480 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END clk
  PIN comb_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 230.335 137.910 234.335 ;
    END
  END comb_output[0]
  PIN comb_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 230.335 151.250 234.335 ;
    END
  END comb_output[1]
  PIN comb_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END comb_output[2]
  PIN comb_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END comb_output[3]
  PIN comb_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 219.615 170.720 223.615 171.320 ;
    END
  END comb_output[4]
  PIN comb_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 219.615 189.080 223.615 189.680 ;
    END
  END comb_output[5]
  PIN comb_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END comb_output[6]
  PIN comb_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END comb_output[7]
  PIN higher_order_address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 230.335 6.810 234.335 ;
    END
  END higher_order_address[0]
  PIN higher_order_address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 230.335 19.690 234.335 ;
    END
  END higher_order_address[1]
  PIN luts_input[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 230.335 33.030 234.335 ;
    END
  END luts_input[0]
  PIN luts_input[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END luts_input[10]
  PIN luts_input[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END luts_input[11]
  PIN luts_input[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END luts_input[12]
  PIN luts_input[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END luts_input[13]
  PIN luts_input[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END luts_input[14]
  PIN luts_input[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END luts_input[15]
  PIN luts_input[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 26.560 223.615 27.160 ;
    END
  END luts_input[16]
  PIN luts_input[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 44.920 223.615 45.520 ;
    END
  END luts_input[17]
  PIN luts_input[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 62.600 223.615 63.200 ;
    END
  END luts_input[18]
  PIN luts_input[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 80.960 223.615 81.560 ;
    END
  END luts_input[19]
  PIN luts_input[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 230.335 45.910 234.335 ;
    END
  END luts_input[1]
  PIN luts_input[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 98.640 223.615 99.240 ;
    END
  END luts_input[20]
  PIN luts_input[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 117.000 223.615 117.600 ;
    END
  END luts_input[21]
  PIN luts_input[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 134.680 223.615 135.280 ;
    END
  END luts_input[22]
  PIN luts_input[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 219.615 153.040 223.615 153.640 ;
    END
  END luts_input[23]
  PIN luts_input[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END luts_input[24]
  PIN luts_input[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END luts_input[25]
  PIN luts_input[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END luts_input[26]
  PIN luts_input[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END luts_input[27]
  PIN luts_input[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END luts_input[28]
  PIN luts_input[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END luts_input[29]
  PIN luts_input[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 230.335 59.250 234.335 ;
    END
  END luts_input[2]
  PIN luts_input[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END luts_input[30]
  PIN luts_input[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END luts_input[31]
  PIN luts_input[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 230.335 72.130 234.335 ;
    END
  END luts_input[3]
  PIN luts_input[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 230.335 85.470 234.335 ;
    END
  END luts_input[4]
  PIN luts_input[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 230.335 98.810 234.335 ;
    END
  END luts_input[5]
  PIN luts_input[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 230.335 111.690 234.335 ;
    END
  END luts_input[6]
  PIN luts_input[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 230.335 125.030 234.335 ;
    END
  END luts_input[7]
  PIN luts_input[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END luts_input[8]
  PIN luts_input[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END luts_input[9]
  PIN reg_we
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END reg_we
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END set_in
  PIN set_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END set_in_soft
  PIN set_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.410 230.335 203.690 234.335 ;
    END
  END set_out
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END shift_in
  PIN shift_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END shift_in_soft
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 230.335 190.810 234.335 ;
    END
  END shift_out
  PIN sync_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.310 230.335 164.590 234.335 ;
    END
  END sync_output[0]
  PIN sync_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.190 230.335 177.470 234.335 ;
    END
  END sync_output[1]
  PIN sync_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END sync_output[2]
  PIN sync_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END sync_output[3]
  PIN sync_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 219.615 206.760 223.615 207.360 ;
    END
  END sync_output[4]
  PIN sync_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 219.615 225.120 223.615 225.720 ;
    END
  END sync_output[5]
  PIN sync_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END sync_output[6]
  PIN sync_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END sync_output[7]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 223.280 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 223.280 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 218.040 223.125 ;
      LAYER met1 ;
        RECT 5.520 5.480 218.040 223.280 ;
      LAYER met2 ;
        RECT 7.090 230.055 19.130 230.335 ;
        RECT 19.970 230.055 32.470 230.335 ;
        RECT 33.310 230.055 45.350 230.335 ;
        RECT 46.190 230.055 58.690 230.335 ;
        RECT 59.530 230.055 71.570 230.335 ;
        RECT 72.410 230.055 84.910 230.335 ;
        RECT 85.750 230.055 98.250 230.335 ;
        RECT 99.090 230.055 111.130 230.335 ;
        RECT 111.970 230.055 124.470 230.335 ;
        RECT 125.310 230.055 137.350 230.335 ;
        RECT 138.190 230.055 150.690 230.335 ;
        RECT 151.530 230.055 164.030 230.335 ;
        RECT 164.870 230.055 176.910 230.335 ;
        RECT 177.750 230.055 190.250 230.335 ;
        RECT 191.090 230.055 203.130 230.335 ;
        RECT 203.970 230.055 216.470 230.335 ;
        RECT 6.540 4.280 217.030 230.055 ;
        RECT 7.090 4.000 19.130 4.280 ;
        RECT 19.970 4.000 32.470 4.280 ;
        RECT 33.310 4.000 45.350 4.280 ;
        RECT 46.190 4.000 58.690 4.280 ;
        RECT 59.530 4.000 71.570 4.280 ;
        RECT 72.410 4.000 84.910 4.280 ;
        RECT 85.750 4.000 98.250 4.280 ;
        RECT 99.090 4.000 111.130 4.280 ;
        RECT 111.970 4.000 124.470 4.280 ;
        RECT 125.310 4.000 137.350 4.280 ;
        RECT 138.190 4.000 150.690 4.280 ;
        RECT 151.530 4.000 164.030 4.280 ;
        RECT 164.870 4.000 176.910 4.280 ;
        RECT 177.750 4.000 190.250 4.280 ;
        RECT 191.090 4.000 203.130 4.280 ;
        RECT 203.970 4.000 216.470 4.280 ;
      LAYER met3 ;
        RECT 4.400 226.120 219.615 226.945 ;
        RECT 4.400 226.080 219.215 226.120 ;
        RECT 4.000 224.720 219.215 226.080 ;
        RECT 4.000 211.840 219.615 224.720 ;
        RECT 4.400 210.440 219.615 211.840 ;
        RECT 4.000 207.760 219.615 210.440 ;
        RECT 4.000 206.360 219.215 207.760 ;
        RECT 4.000 196.200 219.615 206.360 ;
        RECT 4.400 194.800 219.615 196.200 ;
        RECT 4.000 190.080 219.615 194.800 ;
        RECT 4.000 188.680 219.215 190.080 ;
        RECT 4.000 180.560 219.615 188.680 ;
        RECT 4.400 179.160 219.615 180.560 ;
        RECT 4.000 171.720 219.615 179.160 ;
        RECT 4.000 170.320 219.215 171.720 ;
        RECT 4.000 164.920 219.615 170.320 ;
        RECT 4.400 163.520 219.615 164.920 ;
        RECT 4.000 154.040 219.615 163.520 ;
        RECT 4.000 152.640 219.215 154.040 ;
        RECT 4.000 149.280 219.615 152.640 ;
        RECT 4.400 147.880 219.615 149.280 ;
        RECT 4.000 135.680 219.615 147.880 ;
        RECT 4.000 134.280 219.215 135.680 ;
        RECT 4.000 133.640 219.615 134.280 ;
        RECT 4.400 132.240 219.615 133.640 ;
        RECT 4.000 118.000 219.615 132.240 ;
        RECT 4.400 116.600 219.215 118.000 ;
        RECT 4.000 102.360 219.615 116.600 ;
        RECT 4.400 100.960 219.615 102.360 ;
        RECT 4.000 99.640 219.615 100.960 ;
        RECT 4.000 98.240 219.215 99.640 ;
        RECT 4.000 86.720 219.615 98.240 ;
        RECT 4.400 85.320 219.615 86.720 ;
        RECT 4.000 81.960 219.615 85.320 ;
        RECT 4.000 80.560 219.215 81.960 ;
        RECT 4.000 71.080 219.615 80.560 ;
        RECT 4.400 69.680 219.615 71.080 ;
        RECT 4.000 63.600 219.615 69.680 ;
        RECT 4.000 62.200 219.215 63.600 ;
        RECT 4.000 55.440 219.615 62.200 ;
        RECT 4.400 54.040 219.615 55.440 ;
        RECT 4.000 45.920 219.615 54.040 ;
        RECT 4.000 44.520 219.215 45.920 ;
        RECT 4.000 39.800 219.615 44.520 ;
        RECT 4.400 38.400 219.615 39.800 ;
        RECT 4.000 27.560 219.615 38.400 ;
        RECT 4.000 26.160 219.215 27.560 ;
        RECT 4.000 24.160 219.615 26.160 ;
        RECT 4.400 22.760 219.615 24.160 ;
        RECT 4.000 9.880 219.615 22.760 ;
        RECT 4.000 8.520 219.215 9.880 ;
        RECT 4.400 8.480 219.215 8.520 ;
        RECT 4.400 7.120 219.615 8.480 ;
        RECT 4.000 4.255 219.615 7.120 ;
      LAYER met4 ;
        RECT 106.095 10.640 176.240 223.280 ;
  END
END baked_slicel
END LIBRARY

