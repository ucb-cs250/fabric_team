VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 752.620 BY 751.920 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 696.280 53.480 696.880 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 692.190 704.755 692.470 708.755 ;
    END
  END clk
  PIN east_clb_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 56.400 703.395 57.000 ;
    END
  END east_clb_in[0]
  PIN east_clb_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 80.880 703.395 81.480 ;
    END
  END east_clb_in[1]
  PIN east_clb_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 105.360 703.395 105.960 ;
    END
  END east_clb_in[2]
  PIN east_clb_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 129.840 703.395 130.440 ;
    END
  END east_clb_in[3]
  PIN east_clb_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 154.320 703.395 154.920 ;
    END
  END east_clb_in[4]
  PIN east_clb_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 178.800 703.395 179.400 ;
    END
  END east_clb_in[5]
  PIN east_clb_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 203.960 703.395 204.560 ;
    END
  END east_clb_in[6]
  PIN east_clb_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 228.440 703.395 229.040 ;
    END
  END east_clb_in[7]
  PIN east_clb_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 252.920 703.395 253.520 ;
    END
  END east_clb_in[8]
  PIN east_clb_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 699.395 277.400 703.395 278.000 ;
    END
  END east_clb_in[9]
  PIN east_clb_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 301.880 703.395 302.480 ;
    END
  END east_clb_out[0]
  PIN east_clb_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 327.040 703.395 327.640 ;
    END
  END east_clb_out[1]
  PIN east_clb_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 351.520 703.395 352.120 ;
    END
  END east_clb_out[2]
  PIN east_clb_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 376.000 703.395 376.600 ;
    END
  END east_clb_out[3]
  PIN east_clb_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 400.480 703.395 401.080 ;
    END
  END east_clb_out[4]
  PIN east_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 523.560 703.395 524.160 ;
    END
  END east_double[0]
  PIN east_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 548.040 703.395 548.640 ;
    END
  END east_double[1]
  PIN east_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 572.520 703.395 573.120 ;
    END
  END east_double[2]
  PIN east_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 597.680 703.395 598.280 ;
    END
  END east_double[3]
  PIN east_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 622.160 703.395 622.760 ;
    END
  END east_double[4]
  PIN east_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 646.640 703.395 647.240 ;
    END
  END east_double[5]
  PIN east_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 671.120 703.395 671.720 ;
    END
  END east_double[6]
  PIN east_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 695.600 703.395 696.200 ;
    END
  END east_double[7]
  PIN east_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 424.960 703.395 425.560 ;
    END
  END east_single[0]
  PIN east_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 449.440 703.395 450.040 ;
    END
  END east_single[1]
  PIN east_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 474.600 703.395 475.200 ;
    END
  END east_single[2]
  PIN east_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 699.395 499.080 703.395 499.680 ;
    END
  END east_single[3]
  PIN north_clb_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.150 704.755 60.430 708.755 ;
    END
  END north_clb_in[0]
  PIN north_clb_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.770 704.755 82.050 708.755 ;
    END
  END north_clb_in[1]
  PIN north_clb_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.390 704.755 103.670 708.755 ;
    END
  END north_clb_in[2]
  PIN north_clb_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.470 704.755 125.750 708.755 ;
    END
  END north_clb_in[3]
  PIN north_clb_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.090 704.755 147.370 708.755 ;
    END
  END north_clb_in[4]
  PIN north_clb_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.170 704.755 169.450 708.755 ;
    END
  END north_clb_in[5]
  PIN north_clb_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.790 704.755 191.070 708.755 ;
    END
  END north_clb_in[6]
  PIN north_clb_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.410 704.755 212.690 708.755 ;
    END
  END north_clb_in[7]
  PIN north_clb_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.490 704.755 234.770 708.755 ;
    END
  END north_clb_in[8]
  PIN north_clb_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.110 704.755 256.390 708.755 ;
    END
  END north_clb_in[9]
  PIN north_clb_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.190 704.755 278.470 708.755 ;
    END
  END north_clb_out[0]
  PIN north_clb_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.810 704.755 300.090 708.755 ;
    END
  END north_clb_out[1]
  PIN north_clb_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.430 704.755 321.710 708.755 ;
    END
  END north_clb_out[2]
  PIN north_clb_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.510 704.755 343.790 708.755 ;
    END
  END north_clb_out[3]
  PIN north_clb_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.130 704.755 365.410 708.755 ;
    END
  END north_clb_out[4]
  PIN north_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 474.150 704.755 474.430 708.755 ;
    END
  END north_double[0]
  PIN north_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 496.230 704.755 496.510 708.755 ;
    END
  END north_double[1]
  PIN north_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 517.850 704.755 518.130 708.755 ;
    END
  END north_double[2]
  PIN north_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 539.470 704.755 539.750 708.755 ;
    END
  END north_double[3]
  PIN north_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 561.550 704.755 561.830 708.755 ;
    END
  END north_double[4]
  PIN north_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 583.170 704.755 583.450 708.755 ;
    END
  END north_double[5]
  PIN north_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.250 704.755 605.530 708.755 ;
    END
  END north_double[6]
  PIN north_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 626.870 704.755 627.150 708.755 ;
    END
  END north_double[7]
  PIN north_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 387.210 704.755 387.490 708.755 ;
    END
  END north_single[0]
  PIN north_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 408.830 704.755 409.110 708.755 ;
    END
  END north_single[1]
  PIN north_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 430.450 704.755 430.730 708.755 ;
    END
  END north_single[2]
  PIN north_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 452.530 704.755 452.810 708.755 ;
    END
  END north_single[3]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 692.190 44.120 692.470 48.120 ;
    END
  END rst
  PIN set_in_from_north
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.570 704.755 670.850 708.755 ;
    END
  END set_in_from_north
  PIN set_out_to_south
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.570 44.120 670.850 48.120 ;
    END
  END set_out_to_south
  PIN shift_in_from_north
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.490 704.755 648.770 708.755 ;
    END
  END shift_in_from_north
  PIN shift_out_to_south
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 648.490 44.120 648.770 48.120 ;
    END
  END shift_out_to_south
  PIN south_clb_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.150 44.120 60.430 48.120 ;
    END
  END south_clb_in[0]
  PIN south_clb_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.770 44.120 82.050 48.120 ;
    END
  END south_clb_in[1]
  PIN south_clb_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.390 44.120 103.670 48.120 ;
    END
  END south_clb_in[2]
  PIN south_clb_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.470 44.120 125.750 48.120 ;
    END
  END south_clb_in[3]
  PIN south_clb_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.090 44.120 147.370 48.120 ;
    END
  END south_clb_in[4]
  PIN south_clb_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.170 44.120 169.450 48.120 ;
    END
  END south_clb_in[5]
  PIN south_clb_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.790 44.120 191.070 48.120 ;
    END
  END south_clb_in[6]
  PIN south_clb_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.410 44.120 212.690 48.120 ;
    END
  END south_clb_in[7]
  PIN south_clb_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.490 44.120 234.770 48.120 ;
    END
  END south_clb_in[8]
  PIN south_clb_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.110 44.120 256.390 48.120 ;
    END
  END south_clb_in[9]
  PIN south_clb_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.190 44.120 278.470 48.120 ;
    END
  END south_clb_out[0]
  PIN south_clb_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 299.810 44.120 300.090 48.120 ;
    END
  END south_clb_out[1]
  PIN south_clb_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.430 44.120 321.710 48.120 ;
    END
  END south_clb_out[2]
  PIN south_clb_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.510 44.120 343.790 48.120 ;
    END
  END south_clb_out[3]
  PIN south_clb_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.130 44.120 365.410 48.120 ;
    END
  END south_clb_out[4]
  PIN south_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 474.150 44.120 474.430 48.120 ;
    END
  END south_double[0]
  PIN south_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 496.230 44.120 496.510 48.120 ;
    END
  END south_double[1]
  PIN south_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 517.850 44.120 518.130 48.120 ;
    END
  END south_double[2]
  PIN south_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 539.470 44.120 539.750 48.120 ;
    END
  END south_double[3]
  PIN south_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 561.550 44.120 561.830 48.120 ;
    END
  END south_double[4]
  PIN south_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 583.170 44.120 583.450 48.120 ;
    END
  END south_double[5]
  PIN south_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.250 44.120 605.530 48.120 ;
    END
  END south_double[6]
  PIN south_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 626.870 44.120 627.150 48.120 ;
    END
  END south_double[7]
  PIN south_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 387.210 44.120 387.490 48.120 ;
    END
  END south_single[0]
  PIN south_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 408.830 44.120 409.110 48.120 ;
    END
  END south_single[1]
  PIN south_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 430.450 44.120 430.730 48.120 ;
    END
  END south_single[2]
  PIN south_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 452.530 44.120 452.810 48.120 ;
    END
  END south_single[3]
  PIN west_clb_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 55.720 53.480 56.320 ;
    END
  END west_clb_in[0]
  PIN west_clb_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 78.840 53.480 79.440 ;
    END
  END west_clb_in[1]
  PIN west_clb_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 102.640 53.480 103.240 ;
    END
  END west_clb_in[2]
  PIN west_clb_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 126.440 53.480 127.040 ;
    END
  END west_clb_in[3]
  PIN west_clb_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 150.240 53.480 150.840 ;
    END
  END west_clb_in[4]
  PIN west_clb_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 174.040 53.480 174.640 ;
    END
  END west_clb_in[5]
  PIN west_clb_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 197.840 53.480 198.440 ;
    END
  END west_clb_in[6]
  PIN west_clb_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 221.640 53.480 222.240 ;
    END
  END west_clb_in[7]
  PIN west_clb_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 245.440 53.480 246.040 ;
    END
  END west_clb_in[8]
  PIN west_clb_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 269.240 53.480 269.840 ;
    END
  END west_clb_in[9]
  PIN west_clb_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 292.360 53.480 292.960 ;
    END
  END west_clb_out[0]
  PIN west_clb_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 316.160 53.480 316.760 ;
    END
  END west_clb_out[1]
  PIN west_clb_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 339.960 53.480 340.560 ;
    END
  END west_clb_out[2]
  PIN west_clb_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 363.760 53.480 364.360 ;
    END
  END west_clb_out[3]
  PIN west_clb_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 387.560 53.480 388.160 ;
    END
  END west_clb_out[4]
  PIN west_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 505.880 53.480 506.480 ;
    END
  END west_double[0]
  PIN west_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 529.680 53.480 530.280 ;
    END
  END west_double[1]
  PIN west_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 553.480 53.480 554.080 ;
    END
  END west_double[2]
  PIN west_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 577.280 53.480 577.880 ;
    END
  END west_double[3]
  PIN west_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 601.080 53.480 601.680 ;
    END
  END west_double[4]
  PIN west_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 624.880 53.480 625.480 ;
    END
  END west_double[5]
  PIN west_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 648.680 53.480 649.280 ;
    END
  END west_double[6]
  PIN west_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 672.480 53.480 673.080 ;
    END
  END west_double[7]
  PIN west_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 411.360 53.480 411.960 ;
    END
  END west_single[0]
  PIN west_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 435.160 53.480 435.760 ;
    END
  END west_single[1]
  PIN west_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 458.960 53.480 459.560 ;
    END
  END west_single[2]
  PIN west_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 482.760 53.480 483.360 ;
    END
  END west_single[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 727.620 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 752.620 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 697.620 697.005 ;
      LAYER met1 ;
        RECT 55.000 48.580 697.620 697.160 ;
      LAYER met2 ;
        RECT 60.710 704.475 81.490 704.810 ;
        RECT 82.330 704.475 103.110 704.810 ;
        RECT 103.950 704.475 125.190 704.810 ;
        RECT 126.030 704.475 146.810 704.810 ;
        RECT 147.650 704.475 168.890 704.810 ;
        RECT 169.730 704.475 190.510 704.810 ;
        RECT 191.350 704.475 212.130 704.810 ;
        RECT 212.970 704.475 234.210 704.810 ;
        RECT 235.050 704.475 255.830 704.810 ;
        RECT 256.670 704.475 277.910 704.810 ;
        RECT 278.750 704.475 299.530 704.810 ;
        RECT 300.370 704.475 321.150 704.810 ;
        RECT 321.990 704.475 343.230 704.810 ;
        RECT 344.070 704.475 364.850 704.810 ;
        RECT 365.690 704.475 386.930 704.810 ;
        RECT 387.770 704.475 408.550 704.810 ;
        RECT 409.390 704.475 430.170 704.810 ;
        RECT 431.010 704.475 452.250 704.810 ;
        RECT 453.090 704.475 473.870 704.810 ;
        RECT 474.710 704.475 495.950 704.810 ;
        RECT 496.790 704.475 517.570 704.810 ;
        RECT 518.410 704.475 539.190 704.810 ;
        RECT 540.030 704.475 561.270 704.810 ;
        RECT 562.110 704.475 582.890 704.810 ;
        RECT 583.730 704.475 604.970 704.810 ;
        RECT 605.810 704.475 626.590 704.810 ;
        RECT 627.430 704.475 648.210 704.810 ;
        RECT 649.050 704.475 670.290 704.810 ;
        RECT 671.130 704.475 691.910 704.810 ;
        RECT 692.750 704.475 693.380 704.810 ;
        RECT 60.160 48.400 693.380 704.475 ;
        RECT 60.710 48.120 81.490 48.400 ;
        RECT 82.330 48.120 103.110 48.400 ;
        RECT 103.950 48.120 125.190 48.400 ;
        RECT 126.030 48.120 146.810 48.400 ;
        RECT 147.650 48.120 168.890 48.400 ;
        RECT 169.730 48.120 190.510 48.400 ;
        RECT 191.350 48.120 212.130 48.400 ;
        RECT 212.970 48.120 234.210 48.400 ;
        RECT 235.050 48.120 255.830 48.400 ;
        RECT 256.670 48.120 277.910 48.400 ;
        RECT 278.750 48.120 299.530 48.400 ;
        RECT 300.370 48.120 321.150 48.400 ;
        RECT 321.990 48.120 343.230 48.400 ;
        RECT 344.070 48.120 364.850 48.400 ;
        RECT 365.690 48.120 386.930 48.400 ;
        RECT 387.770 48.120 408.550 48.400 ;
        RECT 409.390 48.120 430.170 48.400 ;
        RECT 431.010 48.120 452.250 48.400 ;
        RECT 453.090 48.120 473.870 48.400 ;
        RECT 474.710 48.120 495.950 48.400 ;
        RECT 496.790 48.120 517.570 48.400 ;
        RECT 518.410 48.120 539.190 48.400 ;
        RECT 540.030 48.120 561.270 48.400 ;
        RECT 562.110 48.120 582.890 48.400 ;
        RECT 583.730 48.120 604.970 48.400 ;
        RECT 605.810 48.120 626.590 48.400 ;
        RECT 627.430 48.120 648.210 48.400 ;
        RECT 649.050 48.120 670.290 48.400 ;
        RECT 671.130 48.120 691.910 48.400 ;
        RECT 692.750 48.120 693.380 48.400 ;
      LAYER met3 ;
        RECT 53.880 696.600 699.395 697.085 ;
        RECT 53.880 695.880 698.995 696.600 ;
        RECT 53.480 695.200 698.995 695.880 ;
        RECT 53.480 673.480 699.395 695.200 ;
        RECT 53.880 672.120 699.395 673.480 ;
        RECT 53.880 672.080 698.995 672.120 ;
        RECT 53.480 670.720 698.995 672.080 ;
        RECT 53.480 649.680 699.395 670.720 ;
        RECT 53.880 648.280 699.395 649.680 ;
        RECT 53.480 647.640 699.395 648.280 ;
        RECT 53.480 646.240 698.995 647.640 ;
        RECT 53.480 625.880 699.395 646.240 ;
        RECT 53.880 624.480 699.395 625.880 ;
        RECT 53.480 623.160 699.395 624.480 ;
        RECT 53.480 621.760 698.995 623.160 ;
        RECT 53.480 602.080 699.395 621.760 ;
        RECT 53.880 600.680 699.395 602.080 ;
        RECT 53.480 598.680 699.395 600.680 ;
        RECT 53.480 597.280 698.995 598.680 ;
        RECT 53.480 578.280 699.395 597.280 ;
        RECT 53.880 576.880 699.395 578.280 ;
        RECT 53.480 573.520 699.395 576.880 ;
        RECT 53.480 572.120 698.995 573.520 ;
        RECT 53.480 554.480 699.395 572.120 ;
        RECT 53.880 553.080 699.395 554.480 ;
        RECT 53.480 549.040 699.395 553.080 ;
        RECT 53.480 547.640 698.995 549.040 ;
        RECT 53.480 530.680 699.395 547.640 ;
        RECT 53.880 529.280 699.395 530.680 ;
        RECT 53.480 524.560 699.395 529.280 ;
        RECT 53.480 523.160 698.995 524.560 ;
        RECT 53.480 506.880 699.395 523.160 ;
        RECT 53.880 505.480 699.395 506.880 ;
        RECT 53.480 500.080 699.395 505.480 ;
        RECT 53.480 498.680 698.995 500.080 ;
        RECT 53.480 483.760 699.395 498.680 ;
        RECT 53.880 482.360 699.395 483.760 ;
        RECT 53.480 475.600 699.395 482.360 ;
        RECT 53.480 474.200 698.995 475.600 ;
        RECT 53.480 459.960 699.395 474.200 ;
        RECT 53.880 458.560 699.395 459.960 ;
        RECT 53.480 450.440 699.395 458.560 ;
        RECT 53.480 449.040 698.995 450.440 ;
        RECT 53.480 436.160 699.395 449.040 ;
        RECT 53.880 434.760 699.395 436.160 ;
        RECT 53.480 425.960 699.395 434.760 ;
        RECT 53.480 424.560 698.995 425.960 ;
        RECT 53.480 412.360 699.395 424.560 ;
        RECT 53.880 410.960 699.395 412.360 ;
        RECT 53.480 401.480 699.395 410.960 ;
        RECT 53.480 400.080 698.995 401.480 ;
        RECT 53.480 388.560 699.395 400.080 ;
        RECT 53.880 387.160 699.395 388.560 ;
        RECT 53.480 377.000 699.395 387.160 ;
        RECT 53.480 375.600 698.995 377.000 ;
        RECT 53.480 364.760 699.395 375.600 ;
        RECT 53.880 363.360 699.395 364.760 ;
        RECT 53.480 352.520 699.395 363.360 ;
        RECT 53.480 351.120 698.995 352.520 ;
        RECT 53.480 340.960 699.395 351.120 ;
        RECT 53.880 339.560 699.395 340.960 ;
        RECT 53.480 328.040 699.395 339.560 ;
        RECT 53.480 326.640 698.995 328.040 ;
        RECT 53.480 317.160 699.395 326.640 ;
        RECT 53.880 315.760 699.395 317.160 ;
        RECT 53.480 302.880 699.395 315.760 ;
        RECT 53.480 301.480 698.995 302.880 ;
        RECT 53.480 293.360 699.395 301.480 ;
        RECT 53.880 291.960 699.395 293.360 ;
        RECT 53.480 278.400 699.395 291.960 ;
        RECT 53.480 277.000 698.995 278.400 ;
        RECT 53.480 270.240 699.395 277.000 ;
        RECT 53.880 268.840 699.395 270.240 ;
        RECT 53.480 253.920 699.395 268.840 ;
        RECT 53.480 252.520 698.995 253.920 ;
        RECT 53.480 246.440 699.395 252.520 ;
        RECT 53.880 245.040 699.395 246.440 ;
        RECT 53.480 229.440 699.395 245.040 ;
        RECT 53.480 228.040 698.995 229.440 ;
        RECT 53.480 222.640 699.395 228.040 ;
        RECT 53.880 221.240 699.395 222.640 ;
        RECT 53.480 204.960 699.395 221.240 ;
        RECT 53.480 203.560 698.995 204.960 ;
        RECT 53.480 198.840 699.395 203.560 ;
        RECT 53.880 197.440 699.395 198.840 ;
        RECT 53.480 179.800 699.395 197.440 ;
        RECT 53.480 178.400 698.995 179.800 ;
        RECT 53.480 175.040 699.395 178.400 ;
        RECT 53.880 173.640 699.395 175.040 ;
        RECT 53.480 155.320 699.395 173.640 ;
        RECT 53.480 153.920 698.995 155.320 ;
        RECT 53.480 151.240 699.395 153.920 ;
        RECT 53.880 149.840 699.395 151.240 ;
        RECT 53.480 130.840 699.395 149.840 ;
        RECT 53.480 129.440 698.995 130.840 ;
        RECT 53.480 127.440 699.395 129.440 ;
        RECT 53.880 126.040 699.395 127.440 ;
        RECT 53.480 106.360 699.395 126.040 ;
        RECT 53.480 104.960 698.995 106.360 ;
        RECT 53.480 103.640 699.395 104.960 ;
        RECT 53.880 102.240 699.395 103.640 ;
        RECT 53.480 81.880 699.395 102.240 ;
        RECT 53.480 80.480 698.995 81.880 ;
        RECT 53.480 79.840 699.395 80.480 ;
        RECT 53.880 78.440 699.395 79.840 ;
        RECT 53.480 57.400 699.395 78.440 ;
        RECT 53.480 56.720 698.995 57.400 ;
        RECT 53.880 56.000 698.995 56.720 ;
        RECT 53.880 55.320 699.395 56.000 ;
        RECT 53.480 54.835 699.395 55.320 ;
      LAYER met4 ;
        RECT 0.000 0.000 752.620 751.920 ;
      LAYER met5 ;
        RECT 0.000 70.610 752.620 751.920 ;
  END
END clb_tile
END LIBRARY

