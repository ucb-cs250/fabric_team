VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 678.560 BY 727.440 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.110 680.120 601.390 684.120 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 619.510 44.120 619.790 48.120 ;
    END
  END carry_out
  PIN cb_east_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 55.720 629.480 56.320 ;
    END
  END cb_east_in[0]
  PIN cb_east_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 78.840 629.480 79.440 ;
    END
  END cb_east_in[1]
  PIN cb_east_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 102.640 629.480 103.240 ;
    END
  END cb_east_in[2]
  PIN cb_east_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 126.440 629.480 127.040 ;
    END
  END cb_east_in[3]
  PIN cb_east_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 150.240 629.480 150.840 ;
    END
  END cb_east_in[4]
  PIN cb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 174.040 629.480 174.640 ;
    END
  END cb_east_out[0]
  PIN cb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 197.840 629.480 198.440 ;
    END
  END cb_east_out[1]
  PIN cb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 220.960 629.480 221.560 ;
    END
  END cb_east_out[2]
  PIN cb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 244.760 629.480 245.360 ;
    END
  END cb_east_out[3]
  PIN cb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 268.560 629.480 269.160 ;
    END
  END cb_east_out[4]
  PIN cb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 292.360 629.480 292.960 ;
    END
  END cb_east_out[5]
  PIN cb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 316.160 629.480 316.760 ;
    END
  END cb_east_out[6]
  PIN cb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 339.960 629.480 340.560 ;
    END
  END cb_east_out[7]
  PIN cb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 363.760 629.480 364.360 ;
    END
  END cb_east_out[8]
  PIN cb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 386.880 629.480 387.480 ;
    END
  END cb_east_out[9]
  PIN cb_north_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.770 680.120 59.050 684.120 ;
    END
  END cb_north_in[0]
  PIN cb_north_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.170 680.120 77.450 684.120 ;
    END
  END cb_north_in[1]
  PIN cb_north_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.030 680.120 96.310 684.120 ;
    END
  END cb_north_in[2]
  PIN cb_north_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.890 680.120 115.170 684.120 ;
    END
  END cb_north_in[3]
  PIN cb_north_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.290 680.120 133.570 684.120 ;
    END
  END cb_north_in[4]
  PIN cb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.150 680.120 152.430 684.120 ;
    END
  END cb_north_out[0]
  PIN cb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 171.010 680.120 171.290 684.120 ;
    END
  END cb_north_out[1]
  PIN cb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.410 680.120 189.690 684.120 ;
    END
  END cb_north_out[2]
  PIN cb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.270 680.120 208.550 684.120 ;
    END
  END cb_north_out[3]
  PIN cb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.130 680.120 227.410 684.120 ;
    END
  END cb_north_out[4]
  PIN cb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.530 680.120 245.810 684.120 ;
    END
  END cb_north_out[5]
  PIN cb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.390 680.120 264.670 684.120 ;
    END
  END cb_north_out[6]
  PIN cb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.250 680.120 283.530 684.120 ;
    END
  END cb_north_out[7]
  PIN cb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.650 680.120 301.930 684.120 ;
    END
  END cb_north_out[8]
  PIN cb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.510 680.120 320.790 684.120 ;
    END
  END cb_north_out[9]
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.970 680.120 620.250 684.120 ;
    END
  END cen
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.230 44.120 59.510 48.120 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.550 44.120 78.830 48.120 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.870 44.120 98.150 48.120 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.190 44.120 117.470 48.120 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.510 44.120 136.790 48.120 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.830 44.120 156.110 48.120 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.150 44.120 175.430 48.120 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.470 44.120 194.750 48.120 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.790 44.120 214.070 48.120 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.110 44.120 233.390 48.120 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.430 44.120 252.710 48.120 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 271.750 44.120 272.030 48.120 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.070 44.120 291.350 48.120 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 310.390 44.120 310.670 48.120 ;
    END
  END clb_south_out[3]
  PIN clb_south_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.710 44.120 329.990 48.120 ;
    END
  END clb_south_out[4]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 55.040 53.480 55.640 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 76.800 53.480 77.400 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 98.560 53.480 99.160 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 121.000 53.480 121.600 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 142.760 53.480 143.360 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 165.200 53.480 165.800 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 186.960 53.480 187.560 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 209.400 53.480 210.000 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 231.160 53.480 231.760 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 253.600 53.480 254.200 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 275.360 53.480 275.960 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 297.120 53.480 297.720 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 319.560 53.480 320.160 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 341.320 53.480 341.920 ;
    END
  END clb_west_out[3]
  PIN clb_west_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 363.760 53.480 364.360 ;
    END
  END clb_west_out[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 650.720 53.480 651.320 ;
    END
  END clk
  PIN east_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 505.880 629.480 506.480 ;
    END
  END east_double[0]
  PIN east_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 529.680 629.480 530.280 ;
    END
  END east_double[1]
  PIN east_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 552.800 629.480 553.400 ;
    END
  END east_double[2]
  PIN east_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 576.600 629.480 577.200 ;
    END
  END east_double[3]
  PIN east_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 600.400 629.480 601.000 ;
    END
  END east_double[4]
  PIN east_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 624.200 629.480 624.800 ;
    END
  END east_double[5]
  PIN east_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 648.000 629.480 648.600 ;
    END
  END east_double[6]
  PIN east_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 671.800 629.480 672.400 ;
    END
  END east_double[7]
  PIN east_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 410.680 629.480 411.280 ;
    END
  END east_single[0]
  PIN east_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 434.480 629.480 435.080 ;
    END
  END east_single[1]
  PIN east_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 458.280 629.480 458.880 ;
    END
  END east_single[2]
  PIN east_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 482.080 629.480 482.680 ;
    END
  END east_single[3]
  PIN north_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 413.890 680.120 414.170 684.120 ;
    END
  END north_double[0]
  PIN north_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 432.750 680.120 433.030 684.120 ;
    END
  END north_double[1]
  PIN north_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 451.610 680.120 451.890 684.120 ;
    END
  END north_double[2]
  PIN north_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 470.010 680.120 470.290 684.120 ;
    END
  END north_double[3]
  PIN north_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 488.870 680.120 489.150 684.120 ;
    END
  END north_double[4]
  PIN north_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 507.730 680.120 508.010 684.120 ;
    END
  END north_double[5]
  PIN north_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 526.130 680.120 526.410 684.120 ;
    END
  END north_double[6]
  PIN north_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 544.990 680.120 545.270 684.120 ;
    END
  END north_double[7]
  PIN north_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 339.370 680.120 339.650 684.120 ;
    END
  END north_single[0]
  PIN north_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 357.770 680.120 358.050 684.120 ;
    END
  END north_single[1]
  PIN north_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 376.630 680.120 376.910 684.120 ;
    END
  END north_single[2]
  PIN north_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 395.490 680.120 395.770 684.120 ;
    END
  END north_single[3]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 672.480 53.480 673.080 ;
    END
  END rst
  PIN set_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 600.190 44.120 600.470 48.120 ;
    END
  END set_in_hard
  PIN set_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.250 680.120 582.530 684.120 ;
    END
  END set_out_hard
  PIN shift_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.870 44.120 581.150 48.120 ;
    END
  END shift_in_hard
  PIN shift_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.850 680.120 564.130 684.120 ;
    END
  END shift_out_hard
  PIN south_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 426.310 44.120 426.590 48.120 ;
    END
  END south_double[0]
  PIN south_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 445.630 44.120 445.910 48.120 ;
    END
  END south_double[1]
  PIN south_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 464.950 44.120 465.230 48.120 ;
    END
  END south_double[2]
  PIN south_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 484.270 44.120 484.550 48.120 ;
    END
  END south_double[3]
  PIN south_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 503.590 44.120 503.870 48.120 ;
    END
  END south_double[4]
  PIN south_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 522.910 44.120 523.190 48.120 ;
    END
  END south_double[5]
  PIN south_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 542.230 44.120 542.510 48.120 ;
    END
  END south_double[6]
  PIN south_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 561.550 44.120 561.830 48.120 ;
    END
  END south_double[7]
  PIN south_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 349.030 44.120 349.310 48.120 ;
    END
  END south_single[0]
  PIN south_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 368.350 44.120 368.630 48.120 ;
    END
  END south_single[1]
  PIN south_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 387.670 44.120 387.950 48.120 ;
    END
  END south_single[2]
  PIN south_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 406.990 44.120 407.270 48.120 ;
    END
  END south_single[3]
  PIN west_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 473.920 53.480 474.520 ;
    END
  END west_double[0]
  PIN west_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 495.680 53.480 496.280 ;
    END
  END west_double[1]
  PIN west_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 518.120 53.480 518.720 ;
    END
  END west_double[2]
  PIN west_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 539.880 53.480 540.480 ;
    END
  END west_double[3]
  PIN west_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 562.320 53.480 562.920 ;
    END
  END west_double[4]
  PIN west_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 584.080 53.480 584.680 ;
    END
  END west_double[5]
  PIN west_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 606.520 53.480 607.120 ;
    END
  END west_double[6]
  PIN west_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 628.280 53.480 628.880 ;
    END
  END west_double[7]
  PIN west_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 385.520 53.480 386.120 ;
    END
  END west_single[0]
  PIN west_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 407.960 53.480 408.560 ;
    END
  END west_single[1]
  PIN west_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 429.720 53.480 430.320 ;
    END
  END west_single[2]
  PIN west_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 452.160 53.480 452.760 ;
    END
  END west_single[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 653.560 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 678.560 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 623.560 672.525 ;
      LAYER met1 ;
        RECT 55.000 54.760 623.560 679.880 ;
      LAYER met2 ;
        RECT 56.940 679.840 58.490 680.120 ;
        RECT 59.330 679.840 76.890 680.120 ;
        RECT 77.730 679.840 95.750 680.120 ;
        RECT 96.590 679.840 114.610 680.120 ;
        RECT 115.450 679.840 133.010 680.120 ;
        RECT 133.850 679.840 151.870 680.120 ;
        RECT 152.710 679.840 170.730 680.120 ;
        RECT 171.570 679.840 189.130 680.120 ;
        RECT 189.970 679.840 207.990 680.120 ;
        RECT 208.830 679.840 226.850 680.120 ;
        RECT 227.690 679.840 245.250 680.120 ;
        RECT 246.090 679.840 264.110 680.120 ;
        RECT 264.950 679.840 282.970 680.120 ;
        RECT 283.810 679.840 301.370 680.120 ;
        RECT 302.210 679.840 320.230 680.120 ;
        RECT 321.070 679.840 339.090 680.120 ;
        RECT 339.930 679.840 357.490 680.120 ;
        RECT 358.330 679.840 376.350 680.120 ;
        RECT 377.190 679.840 395.210 680.120 ;
        RECT 396.050 679.840 413.610 680.120 ;
        RECT 414.450 679.840 432.470 680.120 ;
        RECT 433.310 679.840 451.330 680.120 ;
        RECT 452.170 679.840 469.730 680.120 ;
        RECT 470.570 679.840 488.590 680.120 ;
        RECT 489.430 679.840 507.450 680.120 ;
        RECT 508.290 679.840 525.850 680.120 ;
        RECT 526.690 679.840 544.710 680.120 ;
        RECT 545.550 679.840 563.570 680.120 ;
        RECT 564.410 679.840 581.970 680.120 ;
        RECT 582.810 679.840 600.830 680.120 ;
        RECT 601.670 679.840 619.690 680.120 ;
        RECT 56.940 48.400 620.180 679.840 ;
        RECT 56.940 48.120 58.950 48.400 ;
        RECT 59.790 48.120 78.270 48.400 ;
        RECT 79.110 48.120 97.590 48.400 ;
        RECT 98.430 48.120 116.910 48.400 ;
        RECT 117.750 48.120 136.230 48.400 ;
        RECT 137.070 48.120 155.550 48.400 ;
        RECT 156.390 48.120 174.870 48.400 ;
        RECT 175.710 48.120 194.190 48.400 ;
        RECT 195.030 48.120 213.510 48.400 ;
        RECT 214.350 48.120 232.830 48.400 ;
        RECT 233.670 48.120 252.150 48.400 ;
        RECT 252.990 48.120 271.470 48.400 ;
        RECT 272.310 48.120 290.790 48.400 ;
        RECT 291.630 48.120 310.110 48.400 ;
        RECT 310.950 48.120 329.430 48.400 ;
        RECT 330.270 48.120 348.750 48.400 ;
        RECT 349.590 48.120 368.070 48.400 ;
        RECT 368.910 48.120 387.390 48.400 ;
        RECT 388.230 48.120 406.710 48.400 ;
        RECT 407.550 48.120 426.030 48.400 ;
        RECT 426.870 48.120 445.350 48.400 ;
        RECT 446.190 48.120 464.670 48.400 ;
        RECT 465.510 48.120 483.990 48.400 ;
        RECT 484.830 48.120 503.310 48.400 ;
        RECT 504.150 48.120 522.630 48.400 ;
        RECT 523.470 48.120 541.950 48.400 ;
        RECT 542.790 48.120 561.270 48.400 ;
        RECT 562.110 48.120 580.590 48.400 ;
        RECT 581.430 48.120 599.910 48.400 ;
        RECT 600.750 48.120 619.230 48.400 ;
        RECT 620.070 48.120 620.180 48.400 ;
      LAYER met3 ;
        RECT 53.880 672.800 625.480 672.945 ;
        RECT 53.880 672.080 625.080 672.800 ;
        RECT 53.480 671.400 625.080 672.080 ;
        RECT 53.480 651.720 625.480 671.400 ;
        RECT 53.880 650.320 625.480 651.720 ;
        RECT 53.480 649.000 625.480 650.320 ;
        RECT 53.480 647.600 625.080 649.000 ;
        RECT 53.480 629.280 625.480 647.600 ;
        RECT 53.880 627.880 625.480 629.280 ;
        RECT 53.480 625.200 625.480 627.880 ;
        RECT 53.480 623.800 625.080 625.200 ;
        RECT 53.480 607.520 625.480 623.800 ;
        RECT 53.880 606.120 625.480 607.520 ;
        RECT 53.480 601.400 625.480 606.120 ;
        RECT 53.480 600.000 625.080 601.400 ;
        RECT 53.480 585.080 625.480 600.000 ;
        RECT 53.880 583.680 625.480 585.080 ;
        RECT 53.480 577.600 625.480 583.680 ;
        RECT 53.480 576.200 625.080 577.600 ;
        RECT 53.480 563.320 625.480 576.200 ;
        RECT 53.880 561.920 625.480 563.320 ;
        RECT 53.480 553.800 625.480 561.920 ;
        RECT 53.480 552.400 625.080 553.800 ;
        RECT 53.480 540.880 625.480 552.400 ;
        RECT 53.880 539.480 625.480 540.880 ;
        RECT 53.480 530.680 625.480 539.480 ;
        RECT 53.480 529.280 625.080 530.680 ;
        RECT 53.480 519.120 625.480 529.280 ;
        RECT 53.880 517.720 625.480 519.120 ;
        RECT 53.480 506.880 625.480 517.720 ;
        RECT 53.480 505.480 625.080 506.880 ;
        RECT 53.480 496.680 625.480 505.480 ;
        RECT 53.880 495.280 625.480 496.680 ;
        RECT 53.480 483.080 625.480 495.280 ;
        RECT 53.480 481.680 625.080 483.080 ;
        RECT 53.480 474.920 625.480 481.680 ;
        RECT 53.880 473.520 625.480 474.920 ;
        RECT 53.480 459.280 625.480 473.520 ;
        RECT 53.480 457.880 625.080 459.280 ;
        RECT 53.480 453.160 625.480 457.880 ;
        RECT 53.880 451.760 625.480 453.160 ;
        RECT 53.480 435.480 625.480 451.760 ;
        RECT 53.480 434.080 625.080 435.480 ;
        RECT 53.480 430.720 625.480 434.080 ;
        RECT 53.880 429.320 625.480 430.720 ;
        RECT 53.480 411.680 625.480 429.320 ;
        RECT 53.480 410.280 625.080 411.680 ;
        RECT 53.480 408.960 625.480 410.280 ;
        RECT 53.880 407.560 625.480 408.960 ;
        RECT 53.480 387.880 625.480 407.560 ;
        RECT 53.480 386.520 625.080 387.880 ;
        RECT 53.880 386.480 625.080 386.520 ;
        RECT 53.880 385.120 625.480 386.480 ;
        RECT 53.480 364.760 625.480 385.120 ;
        RECT 53.880 363.360 625.080 364.760 ;
        RECT 53.480 342.320 625.480 363.360 ;
        RECT 53.880 340.960 625.480 342.320 ;
        RECT 53.880 340.920 625.080 340.960 ;
        RECT 53.480 339.560 625.080 340.920 ;
        RECT 53.480 320.560 625.480 339.560 ;
        RECT 53.880 319.160 625.480 320.560 ;
        RECT 53.480 317.160 625.480 319.160 ;
        RECT 53.480 315.760 625.080 317.160 ;
        RECT 53.480 298.120 625.480 315.760 ;
        RECT 53.880 296.720 625.480 298.120 ;
        RECT 53.480 293.360 625.480 296.720 ;
        RECT 53.480 291.960 625.080 293.360 ;
        RECT 53.480 276.360 625.480 291.960 ;
        RECT 53.880 274.960 625.480 276.360 ;
        RECT 53.480 269.560 625.480 274.960 ;
        RECT 53.480 268.160 625.080 269.560 ;
        RECT 53.480 254.600 625.480 268.160 ;
        RECT 53.880 253.200 625.480 254.600 ;
        RECT 53.480 245.760 625.480 253.200 ;
        RECT 53.480 244.360 625.080 245.760 ;
        RECT 53.480 232.160 625.480 244.360 ;
        RECT 53.880 230.760 625.480 232.160 ;
        RECT 53.480 221.960 625.480 230.760 ;
        RECT 53.480 220.560 625.080 221.960 ;
        RECT 53.480 210.400 625.480 220.560 ;
        RECT 53.880 209.000 625.480 210.400 ;
        RECT 53.480 198.840 625.480 209.000 ;
        RECT 53.480 197.440 625.080 198.840 ;
        RECT 53.480 187.960 625.480 197.440 ;
        RECT 53.880 186.560 625.480 187.960 ;
        RECT 53.480 175.040 625.480 186.560 ;
        RECT 53.480 173.640 625.080 175.040 ;
        RECT 53.480 166.200 625.480 173.640 ;
        RECT 53.880 164.800 625.480 166.200 ;
        RECT 53.480 151.240 625.480 164.800 ;
        RECT 53.480 149.840 625.080 151.240 ;
        RECT 53.480 143.760 625.480 149.840 ;
        RECT 53.880 142.360 625.480 143.760 ;
        RECT 53.480 127.440 625.480 142.360 ;
        RECT 53.480 126.040 625.080 127.440 ;
        RECT 53.480 122.000 625.480 126.040 ;
        RECT 53.880 120.600 625.480 122.000 ;
        RECT 53.480 103.640 625.480 120.600 ;
        RECT 53.480 102.240 625.080 103.640 ;
        RECT 53.480 99.560 625.480 102.240 ;
        RECT 53.880 98.160 625.480 99.560 ;
        RECT 53.480 79.840 625.480 98.160 ;
        RECT 53.480 78.440 625.080 79.840 ;
        RECT 53.480 77.800 625.480 78.440 ;
        RECT 53.880 76.400 625.480 77.800 ;
        RECT 53.480 56.720 625.480 76.400 ;
        RECT 53.480 56.040 625.080 56.720 ;
        RECT 53.880 55.320 625.080 56.040 ;
        RECT 53.880 54.835 625.480 55.320 ;
      LAYER met4 ;
        RECT 0.000 0.000 678.560 727.440 ;
      LAYER met5 ;
        RECT 0.000 70.610 678.560 727.440 ;
  END
END clb_tile
END LIBRARY

