VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_data_connection_block
  CLASS BLOCK ;
  FOREIGN baked_data_connection_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 1196.000 15.090 1200.000 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 1196.000 3.130 1200.000 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 1196.000 21.070 1200.000 ;
    END
  END cset
  PIN cset_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1194.800 1200.000 1195.400 ;
    END
  END cset_out
  PIN data_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 4.120 1200.000 4.720 ;
    END
  END data_input[0]
  PIN data_input[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 96.600 1200.000 97.200 ;
    END
  END data_input[10]
  PIN data_input[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 106.120 1200.000 106.720 ;
    END
  END data_input[11]
  PIN data_input[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 115.640 1200.000 116.240 ;
    END
  END data_input[12]
  PIN data_input[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 124.480 1200.000 125.080 ;
    END
  END data_input[13]
  PIN data_input[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 134.000 1200.000 134.600 ;
    END
  END data_input[14]
  PIN data_input[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 143.520 1200.000 144.120 ;
    END
  END data_input[15]
  PIN data_input[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 152.360 1200.000 152.960 ;
    END
  END data_input[16]
  PIN data_input[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 161.880 1200.000 162.480 ;
    END
  END data_input[17]
  PIN data_input[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 171.400 1200.000 172.000 ;
    END
  END data_input[18]
  PIN data_input[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 180.240 1200.000 180.840 ;
    END
  END data_input[19]
  PIN data_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 12.960 1200.000 13.560 ;
    END
  END data_input[1]
  PIN data_input[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 189.760 1200.000 190.360 ;
    END
  END data_input[20]
  PIN data_input[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 199.280 1200.000 199.880 ;
    END
  END data_input[21]
  PIN data_input[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 208.800 1200.000 209.400 ;
    END
  END data_input[22]
  PIN data_input[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 217.640 1200.000 218.240 ;
    END
  END data_input[23]
  PIN data_input[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 227.160 1200.000 227.760 ;
    END
  END data_input[24]
  PIN data_input[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 236.680 1200.000 237.280 ;
    END
  END data_input[25]
  PIN data_input[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 245.520 1200.000 246.120 ;
    END
  END data_input[26]
  PIN data_input[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 255.040 1200.000 255.640 ;
    END
  END data_input[27]
  PIN data_input[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 264.560 1200.000 265.160 ;
    END
  END data_input[28]
  PIN data_input[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 273.400 1200.000 274.000 ;
    END
  END data_input[29]
  PIN data_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 22.480 1200.000 23.080 ;
    END
  END data_input[2]
  PIN data_input[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 282.920 1200.000 283.520 ;
    END
  END data_input[30]
  PIN data_input[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 292.440 1200.000 293.040 ;
    END
  END data_input[31]
  PIN data_input[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 301.280 1200.000 301.880 ;
    END
  END data_input[32]
  PIN data_input[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 310.800 1200.000 311.400 ;
    END
  END data_input[33]
  PIN data_input[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 320.320 1200.000 320.920 ;
    END
  END data_input[34]
  PIN data_input[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 329.160 1200.000 329.760 ;
    END
  END data_input[35]
  PIN data_input[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 338.680 1200.000 339.280 ;
    END
  END data_input[36]
  PIN data_input[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 348.200 1200.000 348.800 ;
    END
  END data_input[37]
  PIN data_input[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 357.040 1200.000 357.640 ;
    END
  END data_input[38]
  PIN data_input[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 366.560 1200.000 367.160 ;
    END
  END data_input[39]
  PIN data_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 32.000 1200.000 32.600 ;
    END
  END data_input[3]
  PIN data_input[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 376.080 1200.000 376.680 ;
    END
  END data_input[40]
  PIN data_input[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 384.920 1200.000 385.520 ;
    END
  END data_input[41]
  PIN data_input[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 394.440 1200.000 395.040 ;
    END
  END data_input[42]
  PIN data_input[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 403.960 1200.000 404.560 ;
    END
  END data_input[43]
  PIN data_input[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 413.480 1200.000 414.080 ;
    END
  END data_input[44]
  PIN data_input[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 422.320 1200.000 422.920 ;
    END
  END data_input[45]
  PIN data_input[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 431.840 1200.000 432.440 ;
    END
  END data_input[46]
  PIN data_input[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 441.360 1200.000 441.960 ;
    END
  END data_input[47]
  PIN data_input[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 450.200 1200.000 450.800 ;
    END
  END data_input[48]
  PIN data_input[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 459.720 1200.000 460.320 ;
    END
  END data_input[49]
  PIN data_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 40.840 1200.000 41.440 ;
    END
  END data_input[4]
  PIN data_input[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 469.240 1200.000 469.840 ;
    END
  END data_input[50]
  PIN data_input[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 478.080 1200.000 478.680 ;
    END
  END data_input[51]
  PIN data_input[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 487.600 1200.000 488.200 ;
    END
  END data_input[52]
  PIN data_input[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 497.120 1200.000 497.720 ;
    END
  END data_input[53]
  PIN data_input[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 505.960 1200.000 506.560 ;
    END
  END data_input[54]
  PIN data_input[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 515.480 1200.000 516.080 ;
    END
  END data_input[55]
  PIN data_input[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 525.000 1200.000 525.600 ;
    END
  END data_input[56]
  PIN data_input[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.840 1200.000 534.440 ;
    END
  END data_input[57]
  PIN data_input[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 543.360 1200.000 543.960 ;
    END
  END data_input[58]
  PIN data_input[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 552.880 1200.000 553.480 ;
    END
  END data_input[59]
  PIN data_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 50.360 1200.000 50.960 ;
    END
  END data_input[5]
  PIN data_input[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 561.720 1200.000 562.320 ;
    END
  END data_input[60]
  PIN data_input[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 571.240 1200.000 571.840 ;
    END
  END data_input[61]
  PIN data_input[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 580.760 1200.000 581.360 ;
    END
  END data_input[62]
  PIN data_input[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 589.600 1200.000 590.200 ;
    END
  END data_input[63]
  PIN data_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 59.880 1200.000 60.480 ;
    END
  END data_input[6]
  PIN data_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 68.720 1200.000 69.320 ;
    END
  END data_input[7]
  PIN data_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 78.240 1200.000 78.840 ;
    END
  END data_input[8]
  PIN data_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 87.760 1200.000 88.360 ;
    END
  END data_input[9]
  PIN data_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 599.120 1200.000 599.720 ;
    END
  END data_output[0]
  PIN data_output[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 692.280 1200.000 692.880 ;
    END
  END data_output[10]
  PIN data_output[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 701.800 1200.000 702.400 ;
    END
  END data_output[11]
  PIN data_output[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 710.640 1200.000 711.240 ;
    END
  END data_output[12]
  PIN data_output[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 720.160 1200.000 720.760 ;
    END
  END data_output[13]
  PIN data_output[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 729.680 1200.000 730.280 ;
    END
  END data_output[14]
  PIN data_output[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 738.520 1200.000 739.120 ;
    END
  END data_output[15]
  PIN data_output[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 748.040 1200.000 748.640 ;
    END
  END data_output[16]
  PIN data_output[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 757.560 1200.000 758.160 ;
    END
  END data_output[17]
  PIN data_output[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 766.400 1200.000 767.000 ;
    END
  END data_output[18]
  PIN data_output[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 775.920 1200.000 776.520 ;
    END
  END data_output[19]
  PIN data_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 608.640 1200.000 609.240 ;
    END
  END data_output[1]
  PIN data_output[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 785.440 1200.000 786.040 ;
    END
  END data_output[20]
  PIN data_output[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 794.280 1200.000 794.880 ;
    END
  END data_output[21]
  PIN data_output[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 803.800 1200.000 804.400 ;
    END
  END data_output[22]
  PIN data_output[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 813.320 1200.000 813.920 ;
    END
  END data_output[23]
  PIN data_output[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 822.840 1200.000 823.440 ;
    END
  END data_output[24]
  PIN data_output[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 831.680 1200.000 832.280 ;
    END
  END data_output[25]
  PIN data_output[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 841.200 1200.000 841.800 ;
    END
  END data_output[26]
  PIN data_output[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 850.720 1200.000 851.320 ;
    END
  END data_output[27]
  PIN data_output[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 859.560 1200.000 860.160 ;
    END
  END data_output[28]
  PIN data_output[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 869.080 1200.000 869.680 ;
    END
  END data_output[29]
  PIN data_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 618.160 1200.000 618.760 ;
    END
  END data_output[2]
  PIN data_output[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 878.600 1200.000 879.200 ;
    END
  END data_output[30]
  PIN data_output[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 887.440 1200.000 888.040 ;
    END
  END data_output[31]
  PIN data_output[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 896.960 1200.000 897.560 ;
    END
  END data_output[32]
  PIN data_output[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 906.480 1200.000 907.080 ;
    END
  END data_output[33]
  PIN data_output[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 915.320 1200.000 915.920 ;
    END
  END data_output[34]
  PIN data_output[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 924.840 1200.000 925.440 ;
    END
  END data_output[35]
  PIN data_output[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 934.360 1200.000 934.960 ;
    END
  END data_output[36]
  PIN data_output[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 943.200 1200.000 943.800 ;
    END
  END data_output[37]
  PIN data_output[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 952.720 1200.000 953.320 ;
    END
  END data_output[38]
  PIN data_output[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 962.240 1200.000 962.840 ;
    END
  END data_output[39]
  PIN data_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 627.000 1200.000 627.600 ;
    END
  END data_output[3]
  PIN data_output[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 971.080 1200.000 971.680 ;
    END
  END data_output[40]
  PIN data_output[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 980.600 1200.000 981.200 ;
    END
  END data_output[41]
  PIN data_output[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 990.120 1200.000 990.720 ;
    END
  END data_output[42]
  PIN data_output[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 998.960 1200.000 999.560 ;
    END
  END data_output[43]
  PIN data_output[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1008.480 1200.000 1009.080 ;
    END
  END data_output[44]
  PIN data_output[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1018.000 1200.000 1018.600 ;
    END
  END data_output[45]
  PIN data_output[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1027.520 1200.000 1028.120 ;
    END
  END data_output[46]
  PIN data_output[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1036.360 1200.000 1036.960 ;
    END
  END data_output[47]
  PIN data_output[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1045.880 1200.000 1046.480 ;
    END
  END data_output[48]
  PIN data_output[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1055.400 1200.000 1056.000 ;
    END
  END data_output[49]
  PIN data_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 636.520 1200.000 637.120 ;
    END
  END data_output[4]
  PIN data_output[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1064.240 1200.000 1064.840 ;
    END
  END data_output[50]
  PIN data_output[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1073.760 1200.000 1074.360 ;
    END
  END data_output[51]
  PIN data_output[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1083.280 1200.000 1083.880 ;
    END
  END data_output[52]
  PIN data_output[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1092.120 1200.000 1092.720 ;
    END
  END data_output[53]
  PIN data_output[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1101.640 1200.000 1102.240 ;
    END
  END data_output[54]
  PIN data_output[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1111.160 1200.000 1111.760 ;
    END
  END data_output[55]
  PIN data_output[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1120.000 1200.000 1120.600 ;
    END
  END data_output[56]
  PIN data_output[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1129.520 1200.000 1130.120 ;
    END
  END data_output[57]
  PIN data_output[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1139.040 1200.000 1139.640 ;
    END
  END data_output[58]
  PIN data_output[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1147.880 1200.000 1148.480 ;
    END
  END data_output[59]
  PIN data_output[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 646.040 1200.000 646.640 ;
    END
  END data_output[5]
  PIN data_output[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1157.400 1200.000 1158.000 ;
    END
  END data_output[60]
  PIN data_output[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1166.920 1200.000 1167.520 ;
    END
  END data_output[61]
  PIN data_output[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1175.760 1200.000 1176.360 ;
    END
  END data_output[62]
  PIN data_output[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1185.280 1200.000 1185.880 ;
    END
  END data_output[63]
  PIN data_output[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 654.880 1200.000 655.480 ;
    END
  END data_output[6]
  PIN data_output[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 664.400 1200.000 665.000 ;
    END
  END data_output[7]
  PIN data_output[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 673.920 1200.000 674.520 ;
    END
  END data_output[8]
  PIN data_output[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 682.760 1200.000 683.360 ;
    END
  END data_output[9]
  PIN north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 1196.000 33.030 1200.000 ;
    END
  END north[0]
  PIN north[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 639.030 1196.000 639.310 1200.000 ;
    END
  END north[100]
  PIN north[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 645.010 1196.000 645.290 1200.000 ;
    END
  END north[101]
  PIN north[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 650.990 1196.000 651.270 1200.000 ;
    END
  END north[102]
  PIN north[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 657.430 1196.000 657.710 1200.000 ;
    END
  END north[103]
  PIN north[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 663.410 1196.000 663.690 1200.000 ;
    END
  END north[104]
  PIN north[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 669.390 1196.000 669.670 1200.000 ;
    END
  END north[105]
  PIN north[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 675.370 1196.000 675.650 1200.000 ;
    END
  END north[106]
  PIN north[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 681.350 1196.000 681.630 1200.000 ;
    END
  END north[107]
  PIN north[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 687.330 1196.000 687.610 1200.000 ;
    END
  END north[108]
  PIN north[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 693.770 1196.000 694.050 1200.000 ;
    END
  END north[109]
  PIN north[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 1196.000 93.750 1200.000 ;
    END
  END north[10]
  PIN north[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 699.750 1196.000 700.030 1200.000 ;
    END
  END north[110]
  PIN north[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 705.730 1196.000 706.010 1200.000 ;
    END
  END north[111]
  PIN north[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 711.710 1196.000 711.990 1200.000 ;
    END
  END north[112]
  PIN north[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 1196.000 717.970 1200.000 ;
    END
  END north[113]
  PIN north[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 724.130 1196.000 724.410 1200.000 ;
    END
  END north[114]
  PIN north[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 730.110 1196.000 730.390 1200.000 ;
    END
  END north[115]
  PIN north[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 736.090 1196.000 736.370 1200.000 ;
    END
  END north[116]
  PIN north[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 742.070 1196.000 742.350 1200.000 ;
    END
  END north[117]
  PIN north[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 748.050 1196.000 748.330 1200.000 ;
    END
  END north[118]
  PIN north[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 754.030 1196.000 754.310 1200.000 ;
    END
  END north[119]
  PIN north[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 1196.000 99.730 1200.000 ;
    END
  END north[11]
  PIN north[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 760.470 1196.000 760.750 1200.000 ;
    END
  END north[120]
  PIN north[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 1196.000 766.730 1200.000 ;
    END
  END north[121]
  PIN north[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 772.430 1196.000 772.710 1200.000 ;
    END
  END north[122]
  PIN north[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 778.410 1196.000 778.690 1200.000 ;
    END
  END north[123]
  PIN north[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 784.390 1196.000 784.670 1200.000 ;
    END
  END north[124]
  PIN north[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 790.370 1196.000 790.650 1200.000 ;
    END
  END north[125]
  PIN north[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 796.810 1196.000 797.090 1200.000 ;
    END
  END north[126]
  PIN north[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 802.790 1196.000 803.070 1200.000 ;
    END
  END north[127]
  PIN north[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 808.770 1196.000 809.050 1200.000 ;
    END
  END north[128]
  PIN north[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 814.750 1196.000 815.030 1200.000 ;
    END
  END north[129]
  PIN north[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 1196.000 106.170 1200.000 ;
    END
  END north[12]
  PIN north[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 820.730 1196.000 821.010 1200.000 ;
    END
  END north[130]
  PIN north[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 827.170 1196.000 827.450 1200.000 ;
    END
  END north[131]
  PIN north[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 833.150 1196.000 833.430 1200.000 ;
    END
  END north[132]
  PIN north[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 839.130 1196.000 839.410 1200.000 ;
    END
  END north[133]
  PIN north[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 845.110 1196.000 845.390 1200.000 ;
    END
  END north[134]
  PIN north[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 851.090 1196.000 851.370 1200.000 ;
    END
  END north[135]
  PIN north[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 857.070 1196.000 857.350 1200.000 ;
    END
  END north[136]
  PIN north[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 863.510 1196.000 863.790 1200.000 ;
    END
  END north[137]
  PIN north[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 869.490 1196.000 869.770 1200.000 ;
    END
  END north[138]
  PIN north[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 875.470 1196.000 875.750 1200.000 ;
    END
  END north[139]
  PIN north[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 111.870 1196.000 112.150 1200.000 ;
    END
  END north[13]
  PIN north[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 881.450 1196.000 881.730 1200.000 ;
    END
  END north[140]
  PIN north[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 887.430 1196.000 887.710 1200.000 ;
    END
  END north[141]
  PIN north[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 893.410 1196.000 893.690 1200.000 ;
    END
  END north[142]
  PIN north[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 899.850 1196.000 900.130 1200.000 ;
    END
  END north[143]
  PIN north[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 905.830 1196.000 906.110 1200.000 ;
    END
  END north[144]
  PIN north[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 911.810 1196.000 912.090 1200.000 ;
    END
  END north[145]
  PIN north[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 917.790 1196.000 918.070 1200.000 ;
    END
  END north[146]
  PIN north[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 923.770 1196.000 924.050 1200.000 ;
    END
  END north[147]
  PIN north[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 930.210 1196.000 930.490 1200.000 ;
    END
  END north[148]
  PIN north[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 936.190 1196.000 936.470 1200.000 ;
    END
  END north[149]
  PIN north[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 1196.000 118.130 1200.000 ;
    END
  END north[14]
  PIN north[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 942.170 1196.000 942.450 1200.000 ;
    END
  END north[150]
  PIN north[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 948.150 1196.000 948.430 1200.000 ;
    END
  END north[151]
  PIN north[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 954.130 1196.000 954.410 1200.000 ;
    END
  END north[152]
  PIN north[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 960.110 1196.000 960.390 1200.000 ;
    END
  END north[153]
  PIN north[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 966.550 1196.000 966.830 1200.000 ;
    END
  END north[154]
  PIN north[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 972.530 1196.000 972.810 1200.000 ;
    END
  END north[155]
  PIN north[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 978.510 1196.000 978.790 1200.000 ;
    END
  END north[156]
  PIN north[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 984.490 1196.000 984.770 1200.000 ;
    END
  END north[157]
  PIN north[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 990.470 1196.000 990.750 1200.000 ;
    END
  END north[158]
  PIN north[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 996.450 1196.000 996.730 1200.000 ;
    END
  END north[159]
  PIN north[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 123.830 1196.000 124.110 1200.000 ;
    END
  END north[15]
  PIN north[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1002.890 1196.000 1003.170 1200.000 ;
    END
  END north[160]
  PIN north[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1008.870 1196.000 1009.150 1200.000 ;
    END
  END north[161]
  PIN north[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1014.850 1196.000 1015.130 1200.000 ;
    END
  END north[162]
  PIN north[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1196.000 1021.110 1200.000 ;
    END
  END north[163]
  PIN north[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1026.810 1196.000 1027.090 1200.000 ;
    END
  END north[164]
  PIN north[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1196.000 1033.530 1200.000 ;
    END
  END north[165]
  PIN north[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1039.230 1196.000 1039.510 1200.000 ;
    END
  END north[166]
  PIN north[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1045.210 1196.000 1045.490 1200.000 ;
    END
  END north[167]
  PIN north[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1051.190 1196.000 1051.470 1200.000 ;
    END
  END north[168]
  PIN north[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1057.170 1196.000 1057.450 1200.000 ;
    END
  END north[169]
  PIN north[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 1196.000 130.090 1200.000 ;
    END
  END north[16]
  PIN north[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1063.150 1196.000 1063.430 1200.000 ;
    END
  END north[170]
  PIN north[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 1196.000 1069.870 1200.000 ;
    END
  END north[171]
  PIN north[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 1196.000 1075.850 1200.000 ;
    END
  END north[172]
  PIN north[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1081.550 1196.000 1081.830 1200.000 ;
    END
  END north[173]
  PIN north[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1087.530 1196.000 1087.810 1200.000 ;
    END
  END north[174]
  PIN north[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1093.510 1196.000 1093.790 1200.000 ;
    END
  END north[175]
  PIN north[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1099.490 1196.000 1099.770 1200.000 ;
    END
  END north[176]
  PIN north[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1105.930 1196.000 1106.210 1200.000 ;
    END
  END north[177]
  PIN north[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1111.910 1196.000 1112.190 1200.000 ;
    END
  END north[178]
  PIN north[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1117.890 1196.000 1118.170 1200.000 ;
    END
  END north[179]
  PIN north[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 1196.000 136.070 1200.000 ;
    END
  END north[17]
  PIN north[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1196.000 1124.150 1200.000 ;
    END
  END north[180]
  PIN north[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1129.850 1196.000 1130.130 1200.000 ;
    END
  END north[181]
  PIN north[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1136.290 1196.000 1136.570 1200.000 ;
    END
  END north[182]
  PIN north[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1142.270 1196.000 1142.550 1200.000 ;
    END
  END north[183]
  PIN north[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1148.250 1196.000 1148.530 1200.000 ;
    END
  END north[184]
  PIN north[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1154.230 1196.000 1154.510 1200.000 ;
    END
  END north[185]
  PIN north[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 1196.000 1160.490 1200.000 ;
    END
  END north[186]
  PIN north[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1166.190 1196.000 1166.470 1200.000 ;
    END
  END north[187]
  PIN north[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1172.630 1196.000 1172.910 1200.000 ;
    END
  END north[188]
  PIN north[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1196.000 1178.890 1200.000 ;
    END
  END north[189]
  PIN north[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 142.230 1196.000 142.510 1200.000 ;
    END
  END north[18]
  PIN north[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1184.590 1196.000 1184.870 1200.000 ;
    END
  END north[190]
  PIN north[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1190.570 1196.000 1190.850 1200.000 ;
    END
  END north[191]
  PIN north[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 1196.000 148.490 1200.000 ;
    END
  END north[19]
  PIN north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 1196.000 39.470 1200.000 ;
    END
  END north[1]
  PIN north[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 1196.000 154.470 1200.000 ;
    END
  END north[20]
  PIN north[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 1196.000 160.450 1200.000 ;
    END
  END north[21]
  PIN north[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 166.150 1196.000 166.430 1200.000 ;
    END
  END north[22]
  PIN north[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 1196.000 172.410 1200.000 ;
    END
  END north[23]
  PIN north[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 1196.000 178.850 1200.000 ;
    END
  END north[24]
  PIN north[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 184.550 1196.000 184.830 1200.000 ;
    END
  END north[25]
  PIN north[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 1196.000 190.810 1200.000 ;
    END
  END north[26]
  PIN north[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 196.510 1196.000 196.790 1200.000 ;
    END
  END north[27]
  PIN north[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 1196.000 202.770 1200.000 ;
    END
  END north[28]
  PIN north[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 1196.000 209.210 1200.000 ;
    END
  END north[29]
  PIN north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 1196.000 45.450 1200.000 ;
    END
  END north[2]
  PIN north[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 214.910 1196.000 215.190 1200.000 ;
    END
  END north[30]
  PIN north[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 220.890 1196.000 221.170 1200.000 ;
    END
  END north[31]
  PIN north[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 226.870 1196.000 227.150 1200.000 ;
    END
  END north[32]
  PIN north[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 1196.000 233.130 1200.000 ;
    END
  END north[33]
  PIN north[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 238.830 1196.000 239.110 1200.000 ;
    END
  END north[34]
  PIN north[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 245.270 1196.000 245.550 1200.000 ;
    END
  END north[35]
  PIN north[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 251.250 1196.000 251.530 1200.000 ;
    END
  END north[36]
  PIN north[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 257.230 1196.000 257.510 1200.000 ;
    END
  END north[37]
  PIN north[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 1196.000 263.490 1200.000 ;
    END
  END north[38]
  PIN north[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 1196.000 269.470 1200.000 ;
    END
  END north[39]
  PIN north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 1196.000 51.430 1200.000 ;
    END
  END north[3]
  PIN north[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 275.170 1196.000 275.450 1200.000 ;
    END
  END north[40]
  PIN north[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 1196.000 281.890 1200.000 ;
    END
  END north[41]
  PIN north[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 287.590 1196.000 287.870 1200.000 ;
    END
  END north[42]
  PIN north[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 293.570 1196.000 293.850 1200.000 ;
    END
  END north[43]
  PIN north[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 299.550 1196.000 299.830 1200.000 ;
    END
  END north[44]
  PIN north[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 305.530 1196.000 305.810 1200.000 ;
    END
  END north[45]
  PIN north[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 311.970 1196.000 312.250 1200.000 ;
    END
  END north[46]
  PIN north[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 317.950 1196.000 318.230 1200.000 ;
    END
  END north[47]
  PIN north[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 1196.000 324.210 1200.000 ;
    END
  END north[48]
  PIN north[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 329.910 1196.000 330.190 1200.000 ;
    END
  END north[49]
  PIN north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 1196.000 57.410 1200.000 ;
    END
  END north[4]
  PIN north[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 335.890 1196.000 336.170 1200.000 ;
    END
  END north[50]
  PIN north[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 341.870 1196.000 342.150 1200.000 ;
    END
  END north[51]
  PIN north[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 348.310 1196.000 348.590 1200.000 ;
    END
  END north[52]
  PIN north[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 354.290 1196.000 354.570 1200.000 ;
    END
  END north[53]
  PIN north[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 360.270 1196.000 360.550 1200.000 ;
    END
  END north[54]
  PIN north[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 366.250 1196.000 366.530 1200.000 ;
    END
  END north[55]
  PIN north[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 372.230 1196.000 372.510 1200.000 ;
    END
  END north[56]
  PIN north[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 378.210 1196.000 378.490 1200.000 ;
    END
  END north[57]
  PIN north[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 384.650 1196.000 384.930 1200.000 ;
    END
  END north[58]
  PIN north[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 390.630 1196.000 390.910 1200.000 ;
    END
  END north[59]
  PIN north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 1196.000 63.390 1200.000 ;
    END
  END north[5]
  PIN north[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 396.610 1196.000 396.890 1200.000 ;
    END
  END north[60]
  PIN north[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 402.590 1196.000 402.870 1200.000 ;
    END
  END north[61]
  PIN north[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 1196.000 408.850 1200.000 ;
    END
  END north[62]
  PIN north[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 415.010 1196.000 415.290 1200.000 ;
    END
  END north[63]
  PIN north[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 420.990 1196.000 421.270 1200.000 ;
    END
  END north[64]
  PIN north[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 426.970 1196.000 427.250 1200.000 ;
    END
  END north[65]
  PIN north[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 1196.000 433.230 1200.000 ;
    END
  END north[66]
  PIN north[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 438.930 1196.000 439.210 1200.000 ;
    END
  END north[67]
  PIN north[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 444.910 1196.000 445.190 1200.000 ;
    END
  END north[68]
  PIN north[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 451.350 1196.000 451.630 1200.000 ;
    END
  END north[69]
  PIN north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 1196.000 69.370 1200.000 ;
    END
  END north[6]
  PIN north[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 457.330 1196.000 457.610 1200.000 ;
    END
  END north[70]
  PIN north[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 1196.000 463.590 1200.000 ;
    END
  END north[71]
  PIN north[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 469.290 1196.000 469.570 1200.000 ;
    END
  END north[72]
  PIN north[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 475.270 1196.000 475.550 1200.000 ;
    END
  END north[73]
  PIN north[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 1196.000 481.530 1200.000 ;
    END
  END north[74]
  PIN north[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 487.690 1196.000 487.970 1200.000 ;
    END
  END north[75]
  PIN north[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 493.670 1196.000 493.950 1200.000 ;
    END
  END north[76]
  PIN north[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 499.650 1196.000 499.930 1200.000 ;
    END
  END north[77]
  PIN north[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 505.630 1196.000 505.910 1200.000 ;
    END
  END north[78]
  PIN north[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 511.610 1196.000 511.890 1200.000 ;
    END
  END north[79]
  PIN north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 1196.000 75.810 1200.000 ;
    END
  END north[7]
  PIN north[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 518.050 1196.000 518.330 1200.000 ;
    END
  END north[80]
  PIN north[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 524.030 1196.000 524.310 1200.000 ;
    END
  END north[81]
  PIN north[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 530.010 1196.000 530.290 1200.000 ;
    END
  END north[82]
  PIN north[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 535.990 1196.000 536.270 1200.000 ;
    END
  END north[83]
  PIN north[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 541.970 1196.000 542.250 1200.000 ;
    END
  END north[84]
  PIN north[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 547.950 1196.000 548.230 1200.000 ;
    END
  END north[85]
  PIN north[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 554.390 1196.000 554.670 1200.000 ;
    END
  END north[86]
  PIN north[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 560.370 1196.000 560.650 1200.000 ;
    END
  END north[87]
  PIN north[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 566.350 1196.000 566.630 1200.000 ;
    END
  END north[88]
  PIN north[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 572.330 1196.000 572.610 1200.000 ;
    END
  END north[89]
  PIN north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 1196.000 81.790 1200.000 ;
    END
  END north[8]
  PIN north[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 578.310 1196.000 578.590 1200.000 ;
    END
  END north[90]
  PIN north[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 584.290 1196.000 584.570 1200.000 ;
    END
  END north[91]
  PIN north[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 590.730 1196.000 591.010 1200.000 ;
    END
  END north[92]
  PIN north[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 596.710 1196.000 596.990 1200.000 ;
    END
  END north[93]
  PIN north[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 602.690 1196.000 602.970 1200.000 ;
    END
  END north[94]
  PIN north[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.670 1196.000 608.950 1200.000 ;
    END
  END north[95]
  PIN north[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 614.650 1196.000 614.930 1200.000 ;
    END
  END north[96]
  PIN north[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 621.090 1196.000 621.370 1200.000 ;
    END
  END north[97]
  PIN north[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 627.070 1196.000 627.350 1200.000 ;
    END
  END north[98]
  PIN north[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 633.050 1196.000 633.330 1200.000 ;
    END
  END north[99]
  PIN north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 1196.000 87.770 1200.000 ;
    END
  END north[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 1196.000 9.110 1200.000 ;
    END
  END rst
  PIN set_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END set_soft
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 1196.000 27.050 1200.000 ;
    END
  END shift_in
  PIN shift_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END shift_in_soft
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1196.550 1196.000 1196.830 1200.000 ;
    END
  END shift_out
  PIN south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END south[0]
  PIN south[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END south[100]
  PIN south[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END south[101]
  PIN south[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END south[102]
  PIN south[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END south[103]
  PIN south[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END south[104]
  PIN south[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END south[105]
  PIN south[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END south[106]
  PIN south[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END south[107]
  PIN south[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END south[108]
  PIN south[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END south[109]
  PIN south[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END south[10]
  PIN south[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END south[110]
  PIN south[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END south[111]
  PIN south[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END south[112]
  PIN south[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END south[113]
  PIN south[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END south[114]
  PIN south[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END south[115]
  PIN south[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END south[116]
  PIN south[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END south[117]
  PIN south[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END south[118]
  PIN south[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END south[119]
  PIN south[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END south[11]
  PIN south[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END south[120]
  PIN south[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END south[121]
  PIN south[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END south[122]
  PIN south[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END south[123]
  PIN south[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END south[124]
  PIN south[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END south[125]
  PIN south[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END south[126]
  PIN south[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END south[127]
  PIN south[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END south[128]
  PIN south[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END south[129]
  PIN south[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END south[12]
  PIN south[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END south[130]
  PIN south[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END south[131]
  PIN south[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END south[132]
  PIN south[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END south[133]
  PIN south[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 835.910 0.000 836.190 4.000 ;
    END
  END south[134]
  PIN south[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END south[135]
  PIN south[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END south[136]
  PIN south[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END south[137]
  PIN south[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END south[138]
  PIN south[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END south[139]
  PIN south[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END south[13]
  PIN south[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END south[140]
  PIN south[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END south[141]
  PIN south[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END south[142]
  PIN south[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END south[143]
  PIN south[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END south[144]
  PIN south[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END south[145]
  PIN south[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END south[146]
  PIN south[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END south[147]
  PIN south[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END south[148]
  PIN south[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END south[149]
  PIN south[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END south[14]
  PIN south[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 935.270 0.000 935.550 4.000 ;
    END
  END south[150]
  PIN south[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END south[151]
  PIN south[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END south[152]
  PIN south[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END south[153]
  PIN south[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END south[154]
  PIN south[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END south[155]
  PIN south[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END south[156]
  PIN south[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END south[157]
  PIN south[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END south[158]
  PIN south[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END south[159]
  PIN south[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END south[15]
  PIN south[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END south[160]
  PIN south[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 4.000 ;
    END
  END south[161]
  PIN south[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END south[162]
  PIN south[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END south[163]
  PIN south[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 4.000 ;
    END
  END south[164]
  PIN south[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END south[165]
  PIN south[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END south[166]
  PIN south[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END south[167]
  PIN south[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 4.000 ;
    END
  END south[168]
  PIN south[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1053.490 0.000 1053.770 4.000 ;
    END
  END south[169]
  PIN south[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END south[16]
  PIN south[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1059.930 0.000 1060.210 4.000 ;
    END
  END south[170]
  PIN south[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END south[171]
  PIN south[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END south[172]
  PIN south[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1078.330 0.000 1078.610 4.000 ;
    END
  END south[173]
  PIN south[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END south[174]
  PIN south[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END south[175]
  PIN south[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 4.000 ;
    END
  END south[176]
  PIN south[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1103.170 0.000 1103.450 4.000 ;
    END
  END south[177]
  PIN south[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END south[178]
  PIN south[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 4.000 ;
    END
  END south[179]
  PIN south[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END south[17]
  PIN south[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1122.030 0.000 1122.310 4.000 ;
    END
  END south[180]
  PIN south[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END south[181]
  PIN south[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END south[182]
  PIN south[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1140.430 0.000 1140.710 4.000 ;
    END
  END south[183]
  PIN south[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1146.870 0.000 1147.150 4.000 ;
    END
  END south[184]
  PIN south[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END south[185]
  PIN south[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END south[186]
  PIN south[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1165.270 0.000 1165.550 4.000 ;
    END
  END south[187]
  PIN south[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1171.710 0.000 1171.990 4.000 ;
    END
  END south[188]
  PIN south[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 4.000 ;
    END
  END south[189]
  PIN south[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END south[18]
  PIN south[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END south[190]
  PIN south[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END south[191]
  PIN south[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END south[19]
  PIN south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END south[1]
  PIN south[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END south[20]
  PIN south[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END south[21]
  PIN south[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END south[22]
  PIN south[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END south[23]
  PIN south[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END south[24]
  PIN south[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END south[25]
  PIN south[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END south[26]
  PIN south[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END south[27]
  PIN south[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END south[28]
  PIN south[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END south[29]
  PIN south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END south[2]
  PIN south[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END south[30]
  PIN south[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END south[31]
  PIN south[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END south[32]
  PIN south[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END south[33]
  PIN south[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END south[34]
  PIN south[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END south[35]
  PIN south[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END south[36]
  PIN south[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END south[37]
  PIN south[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END south[38]
  PIN south[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END south[39]
  PIN south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END south[3]
  PIN south[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END south[40]
  PIN south[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END south[41]
  PIN south[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END south[42]
  PIN south[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END south[43]
  PIN south[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END south[44]
  PIN south[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END south[45]
  PIN south[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END south[46]
  PIN south[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END south[47]
  PIN south[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END south[48]
  PIN south[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END south[49]
  PIN south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END south[4]
  PIN south[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END south[50]
  PIN south[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END south[51]
  PIN south[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END south[52]
  PIN south[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END south[53]
  PIN south[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END south[54]
  PIN south[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END south[55]
  PIN south[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END south[56]
  PIN south[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END south[57]
  PIN south[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END south[58]
  PIN south[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END south[59]
  PIN south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END south[5]
  PIN south[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END south[60]
  PIN south[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END south[61]
  PIN south[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END south[62]
  PIN south[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END south[63]
  PIN south[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END south[64]
  PIN south[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END south[65]
  PIN south[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END south[66]
  PIN south[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END south[67]
  PIN south[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END south[68]
  PIN south[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END south[69]
  PIN south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END south[6]
  PIN south[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END south[70]
  PIN south[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END south[71]
  PIN south[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END south[72]
  PIN south[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END south[73]
  PIN south[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END south[74]
  PIN south[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END south[75]
  PIN south[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END south[76]
  PIN south[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END south[77]
  PIN south[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END south[78]
  PIN south[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END south[79]
  PIN south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END south[7]
  PIN south[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END south[80]
  PIN south[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END south[81]
  PIN south[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END south[82]
  PIN south[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END south[83]
  PIN south[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END south[84]
  PIN south[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END south[85]
  PIN south[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END south[86]
  PIN south[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END south[87]
  PIN south[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END south[88]
  PIN south[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END south[89]
  PIN south[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END south[8]
  PIN south[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END south[90]
  PIN south[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END south[91]
  PIN south[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END south[92]
  PIN south[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END south[93]
  PIN south[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END south[94]
  PIN south[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END south[95]
  PIN south[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END south[96]
  PIN south[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END south[97]
  PIN south[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END south[98]
  PIN south[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END south[99]
  PIN south[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END south[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1194.160 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1194.160 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 2.830 5.820 1196.850 1189.620 ;
      LAYER met2 ;
        RECT 0.090 1195.720 2.570 1196.000 ;
        RECT 3.410 1195.720 8.550 1196.000 ;
        RECT 9.390 1195.720 14.530 1196.000 ;
        RECT 15.370 1195.720 20.510 1196.000 ;
        RECT 21.350 1195.720 26.490 1196.000 ;
        RECT 27.330 1195.720 32.470 1196.000 ;
        RECT 33.310 1195.720 38.910 1196.000 ;
        RECT 39.750 1195.720 44.890 1196.000 ;
        RECT 45.730 1195.720 50.870 1196.000 ;
        RECT 51.710 1195.720 56.850 1196.000 ;
        RECT 57.690 1195.720 62.830 1196.000 ;
        RECT 63.670 1195.720 68.810 1196.000 ;
        RECT 69.650 1195.720 75.250 1196.000 ;
        RECT 76.090 1195.720 81.230 1196.000 ;
        RECT 82.070 1195.720 87.210 1196.000 ;
        RECT 88.050 1195.720 93.190 1196.000 ;
        RECT 94.030 1195.720 99.170 1196.000 ;
        RECT 100.010 1195.720 105.610 1196.000 ;
        RECT 106.450 1195.720 111.590 1196.000 ;
        RECT 112.430 1195.720 117.570 1196.000 ;
        RECT 118.410 1195.720 123.550 1196.000 ;
        RECT 124.390 1195.720 129.530 1196.000 ;
        RECT 130.370 1195.720 135.510 1196.000 ;
        RECT 136.350 1195.720 141.950 1196.000 ;
        RECT 142.790 1195.720 147.930 1196.000 ;
        RECT 148.770 1195.720 153.910 1196.000 ;
        RECT 154.750 1195.720 159.890 1196.000 ;
        RECT 160.730 1195.720 165.870 1196.000 ;
        RECT 166.710 1195.720 171.850 1196.000 ;
        RECT 172.690 1195.720 178.290 1196.000 ;
        RECT 179.130 1195.720 184.270 1196.000 ;
        RECT 185.110 1195.720 190.250 1196.000 ;
        RECT 191.090 1195.720 196.230 1196.000 ;
        RECT 197.070 1195.720 202.210 1196.000 ;
        RECT 203.050 1195.720 208.650 1196.000 ;
        RECT 209.490 1195.720 214.630 1196.000 ;
        RECT 215.470 1195.720 220.610 1196.000 ;
        RECT 221.450 1195.720 226.590 1196.000 ;
        RECT 227.430 1195.720 232.570 1196.000 ;
        RECT 233.410 1195.720 238.550 1196.000 ;
        RECT 239.390 1195.720 244.990 1196.000 ;
        RECT 245.830 1195.720 250.970 1196.000 ;
        RECT 251.810 1195.720 256.950 1196.000 ;
        RECT 257.790 1195.720 262.930 1196.000 ;
        RECT 263.770 1195.720 268.910 1196.000 ;
        RECT 269.750 1195.720 274.890 1196.000 ;
        RECT 275.730 1195.720 281.330 1196.000 ;
        RECT 282.170 1195.720 287.310 1196.000 ;
        RECT 288.150 1195.720 293.290 1196.000 ;
        RECT 294.130 1195.720 299.270 1196.000 ;
        RECT 300.110 1195.720 305.250 1196.000 ;
        RECT 306.090 1195.720 311.690 1196.000 ;
        RECT 312.530 1195.720 317.670 1196.000 ;
        RECT 318.510 1195.720 323.650 1196.000 ;
        RECT 324.490 1195.720 329.630 1196.000 ;
        RECT 330.470 1195.720 335.610 1196.000 ;
        RECT 336.450 1195.720 341.590 1196.000 ;
        RECT 342.430 1195.720 348.030 1196.000 ;
        RECT 348.870 1195.720 354.010 1196.000 ;
        RECT 354.850 1195.720 359.990 1196.000 ;
        RECT 360.830 1195.720 365.970 1196.000 ;
        RECT 366.810 1195.720 371.950 1196.000 ;
        RECT 372.790 1195.720 377.930 1196.000 ;
        RECT 378.770 1195.720 384.370 1196.000 ;
        RECT 385.210 1195.720 390.350 1196.000 ;
        RECT 391.190 1195.720 396.330 1196.000 ;
        RECT 397.170 1195.720 402.310 1196.000 ;
        RECT 403.150 1195.720 408.290 1196.000 ;
        RECT 409.130 1195.720 414.730 1196.000 ;
        RECT 415.570 1195.720 420.710 1196.000 ;
        RECT 421.550 1195.720 426.690 1196.000 ;
        RECT 427.530 1195.720 432.670 1196.000 ;
        RECT 433.510 1195.720 438.650 1196.000 ;
        RECT 439.490 1195.720 444.630 1196.000 ;
        RECT 445.470 1195.720 451.070 1196.000 ;
        RECT 451.910 1195.720 457.050 1196.000 ;
        RECT 457.890 1195.720 463.030 1196.000 ;
        RECT 463.870 1195.720 469.010 1196.000 ;
        RECT 469.850 1195.720 474.990 1196.000 ;
        RECT 475.830 1195.720 480.970 1196.000 ;
        RECT 481.810 1195.720 487.410 1196.000 ;
        RECT 488.250 1195.720 493.390 1196.000 ;
        RECT 494.230 1195.720 499.370 1196.000 ;
        RECT 500.210 1195.720 505.350 1196.000 ;
        RECT 506.190 1195.720 511.330 1196.000 ;
        RECT 512.170 1195.720 517.770 1196.000 ;
        RECT 518.610 1195.720 523.750 1196.000 ;
        RECT 524.590 1195.720 529.730 1196.000 ;
        RECT 530.570 1195.720 535.710 1196.000 ;
        RECT 536.550 1195.720 541.690 1196.000 ;
        RECT 542.530 1195.720 547.670 1196.000 ;
        RECT 548.510 1195.720 554.110 1196.000 ;
        RECT 554.950 1195.720 560.090 1196.000 ;
        RECT 560.930 1195.720 566.070 1196.000 ;
        RECT 566.910 1195.720 572.050 1196.000 ;
        RECT 572.890 1195.720 578.030 1196.000 ;
        RECT 578.870 1195.720 584.010 1196.000 ;
        RECT 584.850 1195.720 590.450 1196.000 ;
        RECT 591.290 1195.720 596.430 1196.000 ;
        RECT 597.270 1195.720 602.410 1196.000 ;
        RECT 603.250 1195.720 608.390 1196.000 ;
        RECT 609.230 1195.720 614.370 1196.000 ;
        RECT 615.210 1195.720 620.810 1196.000 ;
        RECT 621.650 1195.720 626.790 1196.000 ;
        RECT 627.630 1195.720 632.770 1196.000 ;
        RECT 633.610 1195.720 638.750 1196.000 ;
        RECT 639.590 1195.720 644.730 1196.000 ;
        RECT 645.570 1195.720 650.710 1196.000 ;
        RECT 651.550 1195.720 657.150 1196.000 ;
        RECT 657.990 1195.720 663.130 1196.000 ;
        RECT 663.970 1195.720 669.110 1196.000 ;
        RECT 669.950 1195.720 675.090 1196.000 ;
        RECT 675.930 1195.720 681.070 1196.000 ;
        RECT 681.910 1195.720 687.050 1196.000 ;
        RECT 687.890 1195.720 693.490 1196.000 ;
        RECT 694.330 1195.720 699.470 1196.000 ;
        RECT 700.310 1195.720 705.450 1196.000 ;
        RECT 706.290 1195.720 711.430 1196.000 ;
        RECT 712.270 1195.720 717.410 1196.000 ;
        RECT 718.250 1195.720 723.850 1196.000 ;
        RECT 724.690 1195.720 729.830 1196.000 ;
        RECT 730.670 1195.720 735.810 1196.000 ;
        RECT 736.650 1195.720 741.790 1196.000 ;
        RECT 742.630 1195.720 747.770 1196.000 ;
        RECT 748.610 1195.720 753.750 1196.000 ;
        RECT 754.590 1195.720 760.190 1196.000 ;
        RECT 761.030 1195.720 766.170 1196.000 ;
        RECT 767.010 1195.720 772.150 1196.000 ;
        RECT 772.990 1195.720 778.130 1196.000 ;
        RECT 778.970 1195.720 784.110 1196.000 ;
        RECT 784.950 1195.720 790.090 1196.000 ;
        RECT 790.930 1195.720 796.530 1196.000 ;
        RECT 797.370 1195.720 802.510 1196.000 ;
        RECT 803.350 1195.720 808.490 1196.000 ;
        RECT 809.330 1195.720 814.470 1196.000 ;
        RECT 815.310 1195.720 820.450 1196.000 ;
        RECT 821.290 1195.720 826.890 1196.000 ;
        RECT 827.730 1195.720 832.870 1196.000 ;
        RECT 833.710 1195.720 838.850 1196.000 ;
        RECT 839.690 1195.720 844.830 1196.000 ;
        RECT 845.670 1195.720 850.810 1196.000 ;
        RECT 851.650 1195.720 856.790 1196.000 ;
        RECT 857.630 1195.720 863.230 1196.000 ;
        RECT 864.070 1195.720 869.210 1196.000 ;
        RECT 870.050 1195.720 875.190 1196.000 ;
        RECT 876.030 1195.720 881.170 1196.000 ;
        RECT 882.010 1195.720 887.150 1196.000 ;
        RECT 887.990 1195.720 893.130 1196.000 ;
        RECT 893.970 1195.720 899.570 1196.000 ;
        RECT 900.410 1195.720 905.550 1196.000 ;
        RECT 906.390 1195.720 911.530 1196.000 ;
        RECT 912.370 1195.720 917.510 1196.000 ;
        RECT 918.350 1195.720 923.490 1196.000 ;
        RECT 924.330 1195.720 929.930 1196.000 ;
        RECT 930.770 1195.720 935.910 1196.000 ;
        RECT 936.750 1195.720 941.890 1196.000 ;
        RECT 942.730 1195.720 947.870 1196.000 ;
        RECT 948.710 1195.720 953.850 1196.000 ;
        RECT 954.690 1195.720 959.830 1196.000 ;
        RECT 960.670 1195.720 966.270 1196.000 ;
        RECT 967.110 1195.720 972.250 1196.000 ;
        RECT 973.090 1195.720 978.230 1196.000 ;
        RECT 979.070 1195.720 984.210 1196.000 ;
        RECT 985.050 1195.720 990.190 1196.000 ;
        RECT 991.030 1195.720 996.170 1196.000 ;
        RECT 997.010 1195.720 1002.610 1196.000 ;
        RECT 1003.450 1195.720 1008.590 1196.000 ;
        RECT 1009.430 1195.720 1014.570 1196.000 ;
        RECT 1015.410 1195.720 1020.550 1196.000 ;
        RECT 1021.390 1195.720 1026.530 1196.000 ;
        RECT 1027.370 1195.720 1032.970 1196.000 ;
        RECT 1033.810 1195.720 1038.950 1196.000 ;
        RECT 1039.790 1195.720 1044.930 1196.000 ;
        RECT 1045.770 1195.720 1050.910 1196.000 ;
        RECT 1051.750 1195.720 1056.890 1196.000 ;
        RECT 1057.730 1195.720 1062.870 1196.000 ;
        RECT 1063.710 1195.720 1069.310 1196.000 ;
        RECT 1070.150 1195.720 1075.290 1196.000 ;
        RECT 1076.130 1195.720 1081.270 1196.000 ;
        RECT 1082.110 1195.720 1087.250 1196.000 ;
        RECT 1088.090 1195.720 1093.230 1196.000 ;
        RECT 1094.070 1195.720 1099.210 1196.000 ;
        RECT 1100.050 1195.720 1105.650 1196.000 ;
        RECT 1106.490 1195.720 1111.630 1196.000 ;
        RECT 1112.470 1195.720 1117.610 1196.000 ;
        RECT 1118.450 1195.720 1123.590 1196.000 ;
        RECT 1124.430 1195.720 1129.570 1196.000 ;
        RECT 1130.410 1195.720 1136.010 1196.000 ;
        RECT 1136.850 1195.720 1141.990 1196.000 ;
        RECT 1142.830 1195.720 1147.970 1196.000 ;
        RECT 1148.810 1195.720 1153.950 1196.000 ;
        RECT 1154.790 1195.720 1159.930 1196.000 ;
        RECT 1160.770 1195.720 1165.910 1196.000 ;
        RECT 1166.750 1195.720 1172.350 1196.000 ;
        RECT 1173.190 1195.720 1178.330 1196.000 ;
        RECT 1179.170 1195.720 1184.310 1196.000 ;
        RECT 1185.150 1195.720 1190.290 1196.000 ;
        RECT 1191.130 1195.720 1196.270 1196.000 ;
        RECT 0.090 4.280 1196.830 1195.720 ;
        RECT 0.090 4.000 2.570 4.280 ;
        RECT 3.410 4.000 8.550 4.280 ;
        RECT 9.390 4.000 14.990 4.280 ;
        RECT 15.830 4.000 20.970 4.280 ;
        RECT 21.810 4.000 27.410 4.280 ;
        RECT 28.250 4.000 33.390 4.280 ;
        RECT 34.230 4.000 39.830 4.280 ;
        RECT 40.670 4.000 45.810 4.280 ;
        RECT 46.650 4.000 52.250 4.280 ;
        RECT 53.090 4.000 58.230 4.280 ;
        RECT 59.070 4.000 64.670 4.280 ;
        RECT 65.510 4.000 70.650 4.280 ;
        RECT 71.490 4.000 77.090 4.280 ;
        RECT 77.930 4.000 83.070 4.280 ;
        RECT 83.910 4.000 89.510 4.280 ;
        RECT 90.350 4.000 95.490 4.280 ;
        RECT 96.330 4.000 101.930 4.280 ;
        RECT 102.770 4.000 107.910 4.280 ;
        RECT 108.750 4.000 114.350 4.280 ;
        RECT 115.190 4.000 120.330 4.280 ;
        RECT 121.170 4.000 126.770 4.280 ;
        RECT 127.610 4.000 132.750 4.280 ;
        RECT 133.590 4.000 139.190 4.280 ;
        RECT 140.030 4.000 145.170 4.280 ;
        RECT 146.010 4.000 151.610 4.280 ;
        RECT 152.450 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.010 4.280 ;
        RECT 170.850 4.000 176.450 4.280 ;
        RECT 177.290 4.000 182.890 4.280 ;
        RECT 183.730 4.000 188.870 4.280 ;
        RECT 189.710 4.000 195.310 4.280 ;
        RECT 196.150 4.000 201.290 4.280 ;
        RECT 202.130 4.000 207.730 4.280 ;
        RECT 208.570 4.000 213.710 4.280 ;
        RECT 214.550 4.000 220.150 4.280 ;
        RECT 220.990 4.000 226.130 4.280 ;
        RECT 226.970 4.000 232.570 4.280 ;
        RECT 233.410 4.000 238.550 4.280 ;
        RECT 239.390 4.000 244.990 4.280 ;
        RECT 245.830 4.000 250.970 4.280 ;
        RECT 251.810 4.000 257.410 4.280 ;
        RECT 258.250 4.000 263.390 4.280 ;
        RECT 264.230 4.000 269.830 4.280 ;
        RECT 270.670 4.000 275.810 4.280 ;
        RECT 276.650 4.000 282.250 4.280 ;
        RECT 283.090 4.000 288.230 4.280 ;
        RECT 289.070 4.000 294.670 4.280 ;
        RECT 295.510 4.000 300.650 4.280 ;
        RECT 301.490 4.000 307.090 4.280 ;
        RECT 307.930 4.000 313.070 4.280 ;
        RECT 313.910 4.000 319.510 4.280 ;
        RECT 320.350 4.000 325.490 4.280 ;
        RECT 326.330 4.000 331.930 4.280 ;
        RECT 332.770 4.000 337.910 4.280 ;
        RECT 338.750 4.000 344.350 4.280 ;
        RECT 345.190 4.000 350.790 4.280 ;
        RECT 351.630 4.000 356.770 4.280 ;
        RECT 357.610 4.000 363.210 4.280 ;
        RECT 364.050 4.000 369.190 4.280 ;
        RECT 370.030 4.000 375.630 4.280 ;
        RECT 376.470 4.000 381.610 4.280 ;
        RECT 382.450 4.000 388.050 4.280 ;
        RECT 388.890 4.000 394.030 4.280 ;
        RECT 394.870 4.000 400.470 4.280 ;
        RECT 401.310 4.000 406.450 4.280 ;
        RECT 407.290 4.000 412.890 4.280 ;
        RECT 413.730 4.000 418.870 4.280 ;
        RECT 419.710 4.000 425.310 4.280 ;
        RECT 426.150 4.000 431.290 4.280 ;
        RECT 432.130 4.000 437.730 4.280 ;
        RECT 438.570 4.000 443.710 4.280 ;
        RECT 444.550 4.000 450.150 4.280 ;
        RECT 450.990 4.000 456.130 4.280 ;
        RECT 456.970 4.000 462.570 4.280 ;
        RECT 463.410 4.000 468.550 4.280 ;
        RECT 469.390 4.000 474.990 4.280 ;
        RECT 475.830 4.000 480.970 4.280 ;
        RECT 481.810 4.000 487.410 4.280 ;
        RECT 488.250 4.000 493.390 4.280 ;
        RECT 494.230 4.000 499.830 4.280 ;
        RECT 500.670 4.000 505.810 4.280 ;
        RECT 506.650 4.000 512.250 4.280 ;
        RECT 513.090 4.000 518.690 4.280 ;
        RECT 519.530 4.000 524.670 4.280 ;
        RECT 525.510 4.000 531.110 4.280 ;
        RECT 531.950 4.000 537.090 4.280 ;
        RECT 537.930 4.000 543.530 4.280 ;
        RECT 544.370 4.000 549.510 4.280 ;
        RECT 550.350 4.000 555.950 4.280 ;
        RECT 556.790 4.000 561.930 4.280 ;
        RECT 562.770 4.000 568.370 4.280 ;
        RECT 569.210 4.000 574.350 4.280 ;
        RECT 575.190 4.000 580.790 4.280 ;
        RECT 581.630 4.000 586.770 4.280 ;
        RECT 587.610 4.000 593.210 4.280 ;
        RECT 594.050 4.000 599.190 4.280 ;
        RECT 600.030 4.000 605.630 4.280 ;
        RECT 606.470 4.000 611.610 4.280 ;
        RECT 612.450 4.000 618.050 4.280 ;
        RECT 618.890 4.000 624.030 4.280 ;
        RECT 624.870 4.000 630.470 4.280 ;
        RECT 631.310 4.000 636.450 4.280 ;
        RECT 637.290 4.000 642.890 4.280 ;
        RECT 643.730 4.000 648.870 4.280 ;
        RECT 649.710 4.000 655.310 4.280 ;
        RECT 656.150 4.000 661.290 4.280 ;
        RECT 662.130 4.000 667.730 4.280 ;
        RECT 668.570 4.000 673.710 4.280 ;
        RECT 674.550 4.000 680.150 4.280 ;
        RECT 680.990 4.000 686.130 4.280 ;
        RECT 686.970 4.000 692.570 4.280 ;
        RECT 693.410 4.000 699.010 4.280 ;
        RECT 699.850 4.000 704.990 4.280 ;
        RECT 705.830 4.000 711.430 4.280 ;
        RECT 712.270 4.000 717.410 4.280 ;
        RECT 718.250 4.000 723.850 4.280 ;
        RECT 724.690 4.000 729.830 4.280 ;
        RECT 730.670 4.000 736.270 4.280 ;
        RECT 737.110 4.000 742.250 4.280 ;
        RECT 743.090 4.000 748.690 4.280 ;
        RECT 749.530 4.000 754.670 4.280 ;
        RECT 755.510 4.000 761.110 4.280 ;
        RECT 761.950 4.000 767.090 4.280 ;
        RECT 767.930 4.000 773.530 4.280 ;
        RECT 774.370 4.000 779.510 4.280 ;
        RECT 780.350 4.000 785.950 4.280 ;
        RECT 786.790 4.000 791.930 4.280 ;
        RECT 792.770 4.000 798.370 4.280 ;
        RECT 799.210 4.000 804.350 4.280 ;
        RECT 805.190 4.000 810.790 4.280 ;
        RECT 811.630 4.000 816.770 4.280 ;
        RECT 817.610 4.000 823.210 4.280 ;
        RECT 824.050 4.000 829.190 4.280 ;
        RECT 830.030 4.000 835.630 4.280 ;
        RECT 836.470 4.000 841.610 4.280 ;
        RECT 842.450 4.000 848.050 4.280 ;
        RECT 848.890 4.000 854.030 4.280 ;
        RECT 854.870 4.000 860.470 4.280 ;
        RECT 861.310 4.000 866.910 4.280 ;
        RECT 867.750 4.000 872.890 4.280 ;
        RECT 873.730 4.000 879.330 4.280 ;
        RECT 880.170 4.000 885.310 4.280 ;
        RECT 886.150 4.000 891.750 4.280 ;
        RECT 892.590 4.000 897.730 4.280 ;
        RECT 898.570 4.000 904.170 4.280 ;
        RECT 905.010 4.000 910.150 4.280 ;
        RECT 910.990 4.000 916.590 4.280 ;
        RECT 917.430 4.000 922.570 4.280 ;
        RECT 923.410 4.000 929.010 4.280 ;
        RECT 929.850 4.000 934.990 4.280 ;
        RECT 935.830 4.000 941.430 4.280 ;
        RECT 942.270 4.000 947.410 4.280 ;
        RECT 948.250 4.000 953.850 4.280 ;
        RECT 954.690 4.000 959.830 4.280 ;
        RECT 960.670 4.000 966.270 4.280 ;
        RECT 967.110 4.000 972.250 4.280 ;
        RECT 973.090 4.000 978.690 4.280 ;
        RECT 979.530 4.000 984.670 4.280 ;
        RECT 985.510 4.000 991.110 4.280 ;
        RECT 991.950 4.000 997.090 4.280 ;
        RECT 997.930 4.000 1003.530 4.280 ;
        RECT 1004.370 4.000 1009.510 4.280 ;
        RECT 1010.350 4.000 1015.950 4.280 ;
        RECT 1016.790 4.000 1021.930 4.280 ;
        RECT 1022.770 4.000 1028.370 4.280 ;
        RECT 1029.210 4.000 1034.810 4.280 ;
        RECT 1035.650 4.000 1040.790 4.280 ;
        RECT 1041.630 4.000 1047.230 4.280 ;
        RECT 1048.070 4.000 1053.210 4.280 ;
        RECT 1054.050 4.000 1059.650 4.280 ;
        RECT 1060.490 4.000 1065.630 4.280 ;
        RECT 1066.470 4.000 1072.070 4.280 ;
        RECT 1072.910 4.000 1078.050 4.280 ;
        RECT 1078.890 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1090.470 4.280 ;
        RECT 1091.310 4.000 1096.910 4.280 ;
        RECT 1097.750 4.000 1102.890 4.280 ;
        RECT 1103.730 4.000 1109.330 4.280 ;
        RECT 1110.170 4.000 1115.310 4.280 ;
        RECT 1116.150 4.000 1121.750 4.280 ;
        RECT 1122.590 4.000 1127.730 4.280 ;
        RECT 1128.570 4.000 1134.170 4.280 ;
        RECT 1135.010 4.000 1140.150 4.280 ;
        RECT 1140.990 4.000 1146.590 4.280 ;
        RECT 1147.430 4.000 1152.570 4.280 ;
        RECT 1153.410 4.000 1159.010 4.280 ;
        RECT 1159.850 4.000 1164.990 4.280 ;
        RECT 1165.830 4.000 1171.430 4.280 ;
        RECT 1172.270 4.000 1177.410 4.280 ;
        RECT 1178.250 4.000 1183.850 4.280 ;
        RECT 1184.690 4.000 1189.830 4.280 ;
        RECT 1190.670 4.000 1196.270 4.280 ;
      LAYER met3 ;
        RECT 0.065 1194.400 1195.600 1195.265 ;
        RECT 0.065 1186.280 1196.855 1194.400 ;
        RECT 0.065 1184.880 1195.600 1186.280 ;
        RECT 0.065 1176.760 1196.855 1184.880 ;
        RECT 0.065 1175.360 1195.600 1176.760 ;
        RECT 0.065 1167.920 1196.855 1175.360 ;
        RECT 0.065 1166.520 1195.600 1167.920 ;
        RECT 0.065 1158.400 1196.855 1166.520 ;
        RECT 0.065 1157.000 1195.600 1158.400 ;
        RECT 0.065 1148.880 1196.855 1157.000 ;
        RECT 0.065 1147.480 1195.600 1148.880 ;
        RECT 0.065 1140.040 1196.855 1147.480 ;
        RECT 0.065 1138.640 1195.600 1140.040 ;
        RECT 0.065 1130.520 1196.855 1138.640 ;
        RECT 0.065 1129.120 1195.600 1130.520 ;
        RECT 0.065 1121.000 1196.855 1129.120 ;
        RECT 0.065 1119.600 1195.600 1121.000 ;
        RECT 0.065 1112.160 1196.855 1119.600 ;
        RECT 0.065 1110.760 1195.600 1112.160 ;
        RECT 0.065 1102.640 1196.855 1110.760 ;
        RECT 0.065 1101.240 1195.600 1102.640 ;
        RECT 0.065 1093.120 1196.855 1101.240 ;
        RECT 0.065 1091.720 1195.600 1093.120 ;
        RECT 0.065 1084.280 1196.855 1091.720 ;
        RECT 0.065 1082.880 1195.600 1084.280 ;
        RECT 0.065 1074.760 1196.855 1082.880 ;
        RECT 0.065 1073.360 1195.600 1074.760 ;
        RECT 0.065 1065.240 1196.855 1073.360 ;
        RECT 0.065 1063.840 1195.600 1065.240 ;
        RECT 0.065 1056.400 1196.855 1063.840 ;
        RECT 0.065 1055.000 1195.600 1056.400 ;
        RECT 0.065 1046.880 1196.855 1055.000 ;
        RECT 0.065 1045.480 1195.600 1046.880 ;
        RECT 0.065 1037.360 1196.855 1045.480 ;
        RECT 0.065 1035.960 1195.600 1037.360 ;
        RECT 0.065 1028.520 1196.855 1035.960 ;
        RECT 0.065 1027.120 1195.600 1028.520 ;
        RECT 0.065 1019.000 1196.855 1027.120 ;
        RECT 0.065 1017.600 1195.600 1019.000 ;
        RECT 0.065 1009.480 1196.855 1017.600 ;
        RECT 0.065 1008.080 1195.600 1009.480 ;
        RECT 0.065 999.960 1196.855 1008.080 ;
        RECT 0.065 998.560 1195.600 999.960 ;
        RECT 0.065 991.120 1196.855 998.560 ;
        RECT 0.065 989.720 1195.600 991.120 ;
        RECT 0.065 981.600 1196.855 989.720 ;
        RECT 0.065 980.200 1195.600 981.600 ;
        RECT 0.065 972.080 1196.855 980.200 ;
        RECT 0.065 970.680 1195.600 972.080 ;
        RECT 0.065 963.240 1196.855 970.680 ;
        RECT 0.065 961.840 1195.600 963.240 ;
        RECT 0.065 953.720 1196.855 961.840 ;
        RECT 0.065 952.320 1195.600 953.720 ;
        RECT 0.065 944.200 1196.855 952.320 ;
        RECT 0.065 942.800 1195.600 944.200 ;
        RECT 0.065 935.360 1196.855 942.800 ;
        RECT 0.065 933.960 1195.600 935.360 ;
        RECT 0.065 925.840 1196.855 933.960 ;
        RECT 0.065 924.440 1195.600 925.840 ;
        RECT 0.065 916.320 1196.855 924.440 ;
        RECT 0.065 914.920 1195.600 916.320 ;
        RECT 0.065 907.480 1196.855 914.920 ;
        RECT 0.065 906.080 1195.600 907.480 ;
        RECT 0.065 897.960 1196.855 906.080 ;
        RECT 0.065 896.560 1195.600 897.960 ;
        RECT 0.065 888.440 1196.855 896.560 ;
        RECT 0.065 887.040 1195.600 888.440 ;
        RECT 0.065 879.600 1196.855 887.040 ;
        RECT 0.065 878.200 1195.600 879.600 ;
        RECT 0.065 870.080 1196.855 878.200 ;
        RECT 0.065 868.680 1195.600 870.080 ;
        RECT 0.065 860.560 1196.855 868.680 ;
        RECT 0.065 859.160 1195.600 860.560 ;
        RECT 0.065 851.720 1196.855 859.160 ;
        RECT 0.065 850.320 1195.600 851.720 ;
        RECT 0.065 842.200 1196.855 850.320 ;
        RECT 0.065 840.800 1195.600 842.200 ;
        RECT 0.065 832.680 1196.855 840.800 ;
        RECT 0.065 831.280 1195.600 832.680 ;
        RECT 0.065 823.840 1196.855 831.280 ;
        RECT 0.065 822.440 1195.600 823.840 ;
        RECT 0.065 814.320 1196.855 822.440 ;
        RECT 0.065 812.920 1195.600 814.320 ;
        RECT 0.065 804.800 1196.855 812.920 ;
        RECT 0.065 803.400 1195.600 804.800 ;
        RECT 0.065 795.280 1196.855 803.400 ;
        RECT 0.065 793.880 1195.600 795.280 ;
        RECT 0.065 786.440 1196.855 793.880 ;
        RECT 0.065 785.040 1195.600 786.440 ;
        RECT 0.065 776.920 1196.855 785.040 ;
        RECT 0.065 775.520 1195.600 776.920 ;
        RECT 0.065 767.400 1196.855 775.520 ;
        RECT 0.065 766.000 1195.600 767.400 ;
        RECT 0.065 758.560 1196.855 766.000 ;
        RECT 0.065 757.160 1195.600 758.560 ;
        RECT 0.065 749.040 1196.855 757.160 ;
        RECT 0.065 747.640 1195.600 749.040 ;
        RECT 0.065 739.520 1196.855 747.640 ;
        RECT 0.065 738.120 1195.600 739.520 ;
        RECT 0.065 730.680 1196.855 738.120 ;
        RECT 0.065 729.280 1195.600 730.680 ;
        RECT 0.065 721.160 1196.855 729.280 ;
        RECT 0.065 719.760 1195.600 721.160 ;
        RECT 0.065 711.640 1196.855 719.760 ;
        RECT 0.065 710.240 1195.600 711.640 ;
        RECT 0.065 702.800 1196.855 710.240 ;
        RECT 0.065 701.400 1195.600 702.800 ;
        RECT 0.065 693.280 1196.855 701.400 ;
        RECT 0.065 691.880 1195.600 693.280 ;
        RECT 0.065 683.760 1196.855 691.880 ;
        RECT 0.065 682.360 1195.600 683.760 ;
        RECT 0.065 674.920 1196.855 682.360 ;
        RECT 0.065 673.520 1195.600 674.920 ;
        RECT 0.065 665.400 1196.855 673.520 ;
        RECT 0.065 664.000 1195.600 665.400 ;
        RECT 0.065 655.880 1196.855 664.000 ;
        RECT 0.065 654.480 1195.600 655.880 ;
        RECT 0.065 647.040 1196.855 654.480 ;
        RECT 0.065 645.640 1195.600 647.040 ;
        RECT 0.065 637.520 1196.855 645.640 ;
        RECT 0.065 636.120 1195.600 637.520 ;
        RECT 0.065 628.000 1196.855 636.120 ;
        RECT 0.065 626.600 1195.600 628.000 ;
        RECT 0.065 619.160 1196.855 626.600 ;
        RECT 0.065 617.760 1195.600 619.160 ;
        RECT 0.065 609.640 1196.855 617.760 ;
        RECT 0.065 608.240 1195.600 609.640 ;
        RECT 0.065 600.800 1196.855 608.240 ;
        RECT 4.400 600.120 1196.855 600.800 ;
        RECT 4.400 599.400 1195.600 600.120 ;
        RECT 0.065 598.720 1195.600 599.400 ;
        RECT 0.065 590.600 1196.855 598.720 ;
        RECT 0.065 589.200 1195.600 590.600 ;
        RECT 0.065 581.760 1196.855 589.200 ;
        RECT 0.065 580.360 1195.600 581.760 ;
        RECT 0.065 572.240 1196.855 580.360 ;
        RECT 0.065 570.840 1195.600 572.240 ;
        RECT 0.065 562.720 1196.855 570.840 ;
        RECT 0.065 561.320 1195.600 562.720 ;
        RECT 0.065 553.880 1196.855 561.320 ;
        RECT 0.065 552.480 1195.600 553.880 ;
        RECT 0.065 544.360 1196.855 552.480 ;
        RECT 0.065 542.960 1195.600 544.360 ;
        RECT 0.065 534.840 1196.855 542.960 ;
        RECT 0.065 533.440 1195.600 534.840 ;
        RECT 0.065 526.000 1196.855 533.440 ;
        RECT 0.065 524.600 1195.600 526.000 ;
        RECT 0.065 516.480 1196.855 524.600 ;
        RECT 0.065 515.080 1195.600 516.480 ;
        RECT 0.065 506.960 1196.855 515.080 ;
        RECT 0.065 505.560 1195.600 506.960 ;
        RECT 0.065 498.120 1196.855 505.560 ;
        RECT 0.065 496.720 1195.600 498.120 ;
        RECT 0.065 488.600 1196.855 496.720 ;
        RECT 0.065 487.200 1195.600 488.600 ;
        RECT 0.065 479.080 1196.855 487.200 ;
        RECT 0.065 477.680 1195.600 479.080 ;
        RECT 0.065 470.240 1196.855 477.680 ;
        RECT 0.065 468.840 1195.600 470.240 ;
        RECT 0.065 460.720 1196.855 468.840 ;
        RECT 0.065 459.320 1195.600 460.720 ;
        RECT 0.065 451.200 1196.855 459.320 ;
        RECT 0.065 449.800 1195.600 451.200 ;
        RECT 0.065 442.360 1196.855 449.800 ;
        RECT 0.065 440.960 1195.600 442.360 ;
        RECT 0.065 432.840 1196.855 440.960 ;
        RECT 0.065 431.440 1195.600 432.840 ;
        RECT 0.065 423.320 1196.855 431.440 ;
        RECT 0.065 421.920 1195.600 423.320 ;
        RECT 0.065 414.480 1196.855 421.920 ;
        RECT 0.065 413.080 1195.600 414.480 ;
        RECT 0.065 404.960 1196.855 413.080 ;
        RECT 0.065 403.560 1195.600 404.960 ;
        RECT 0.065 395.440 1196.855 403.560 ;
        RECT 0.065 394.040 1195.600 395.440 ;
        RECT 0.065 385.920 1196.855 394.040 ;
        RECT 0.065 384.520 1195.600 385.920 ;
        RECT 0.065 377.080 1196.855 384.520 ;
        RECT 0.065 375.680 1195.600 377.080 ;
        RECT 0.065 367.560 1196.855 375.680 ;
        RECT 0.065 366.160 1195.600 367.560 ;
        RECT 0.065 358.040 1196.855 366.160 ;
        RECT 0.065 356.640 1195.600 358.040 ;
        RECT 0.065 349.200 1196.855 356.640 ;
        RECT 0.065 347.800 1195.600 349.200 ;
        RECT 0.065 339.680 1196.855 347.800 ;
        RECT 0.065 338.280 1195.600 339.680 ;
        RECT 0.065 330.160 1196.855 338.280 ;
        RECT 0.065 328.760 1195.600 330.160 ;
        RECT 0.065 321.320 1196.855 328.760 ;
        RECT 0.065 319.920 1195.600 321.320 ;
        RECT 0.065 311.800 1196.855 319.920 ;
        RECT 0.065 310.400 1195.600 311.800 ;
        RECT 0.065 302.280 1196.855 310.400 ;
        RECT 0.065 300.880 1195.600 302.280 ;
        RECT 0.065 293.440 1196.855 300.880 ;
        RECT 0.065 292.040 1195.600 293.440 ;
        RECT 0.065 283.920 1196.855 292.040 ;
        RECT 0.065 282.520 1195.600 283.920 ;
        RECT 0.065 274.400 1196.855 282.520 ;
        RECT 0.065 273.000 1195.600 274.400 ;
        RECT 0.065 265.560 1196.855 273.000 ;
        RECT 0.065 264.160 1195.600 265.560 ;
        RECT 0.065 256.040 1196.855 264.160 ;
        RECT 0.065 254.640 1195.600 256.040 ;
        RECT 0.065 246.520 1196.855 254.640 ;
        RECT 0.065 245.120 1195.600 246.520 ;
        RECT 0.065 237.680 1196.855 245.120 ;
        RECT 0.065 236.280 1195.600 237.680 ;
        RECT 0.065 228.160 1196.855 236.280 ;
        RECT 0.065 226.760 1195.600 228.160 ;
        RECT 0.065 218.640 1196.855 226.760 ;
        RECT 0.065 217.240 1195.600 218.640 ;
        RECT 0.065 209.800 1196.855 217.240 ;
        RECT 0.065 208.400 1195.600 209.800 ;
        RECT 0.065 200.280 1196.855 208.400 ;
        RECT 0.065 198.880 1195.600 200.280 ;
        RECT 0.065 190.760 1196.855 198.880 ;
        RECT 0.065 189.360 1195.600 190.760 ;
        RECT 0.065 181.240 1196.855 189.360 ;
        RECT 0.065 179.840 1195.600 181.240 ;
        RECT 0.065 172.400 1196.855 179.840 ;
        RECT 0.065 171.000 1195.600 172.400 ;
        RECT 0.065 162.880 1196.855 171.000 ;
        RECT 0.065 161.480 1195.600 162.880 ;
        RECT 0.065 153.360 1196.855 161.480 ;
        RECT 0.065 151.960 1195.600 153.360 ;
        RECT 0.065 144.520 1196.855 151.960 ;
        RECT 0.065 143.120 1195.600 144.520 ;
        RECT 0.065 135.000 1196.855 143.120 ;
        RECT 0.065 133.600 1195.600 135.000 ;
        RECT 0.065 125.480 1196.855 133.600 ;
        RECT 0.065 124.080 1195.600 125.480 ;
        RECT 0.065 116.640 1196.855 124.080 ;
        RECT 0.065 115.240 1195.600 116.640 ;
        RECT 0.065 107.120 1196.855 115.240 ;
        RECT 0.065 105.720 1195.600 107.120 ;
        RECT 0.065 97.600 1196.855 105.720 ;
        RECT 0.065 96.200 1195.600 97.600 ;
        RECT 0.065 88.760 1196.855 96.200 ;
        RECT 0.065 87.360 1195.600 88.760 ;
        RECT 0.065 79.240 1196.855 87.360 ;
        RECT 0.065 77.840 1195.600 79.240 ;
        RECT 0.065 69.720 1196.855 77.840 ;
        RECT 0.065 68.320 1195.600 69.720 ;
        RECT 0.065 60.880 1196.855 68.320 ;
        RECT 0.065 59.480 1195.600 60.880 ;
        RECT 0.065 51.360 1196.855 59.480 ;
        RECT 0.065 49.960 1195.600 51.360 ;
        RECT 0.065 41.840 1196.855 49.960 ;
        RECT 0.065 40.440 1195.600 41.840 ;
        RECT 0.065 33.000 1196.855 40.440 ;
        RECT 0.065 31.600 1195.600 33.000 ;
        RECT 0.065 23.480 1196.855 31.600 ;
        RECT 0.065 22.080 1195.600 23.480 ;
        RECT 0.065 13.960 1196.855 22.080 ;
        RECT 0.065 12.560 1195.600 13.960 ;
        RECT 0.065 5.120 1196.855 12.560 ;
        RECT 0.065 4.255 1195.600 5.120 ;
      LAYER met4 ;
        RECT 14.095 10.640 1174.640 1188.880 ;
      LAYER met5 ;
        RECT 5.520 179.670 1194.160 1176.940 ;
  END
END baked_data_connection_block
END LIBRARY

