magic
tech sky130A
magscale 1 2
timestamp 1623552508
<< obsli1 >>
rect 121 1377 12483 13073
<< obsm1 >>
rect 14 892 13326 13524
<< metal2 >>
rect 754 14818 810 15618
rect 2226 14818 2282 15618
rect 3698 14818 3754 15618
rect 5170 14818 5226 15618
rect 6642 14818 6698 15618
rect 8206 14818 8262 15618
rect 9678 14818 9734 15618
rect 11150 14818 11206 15618
rect 12622 14818 12678 15618
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 386 0 442 800
rect 478 0 534 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
<< obsm2 >>
rect 20 14762 698 14818
rect 866 14762 2170 14818
rect 2338 14762 3642 14818
rect 3810 14762 5114 14818
rect 5282 14762 6586 14818
rect 6754 14762 8150 14818
rect 8318 14762 9622 14818
rect 9790 14762 11094 14818
rect 11262 14762 12566 14818
rect 12734 14762 13320 14818
rect 20 856 13320 14762
rect 314 800 330 856
rect 590 800 606 856
rect 958 800 974 856
rect 1234 800 1250 856
rect 1602 800 1618 856
rect 1878 800 1894 856
rect 2246 800 2262 856
rect 2522 800 2538 856
rect 2890 800 2906 856
rect 3166 800 3182 856
rect 3534 800 3550 856
rect 3810 800 3826 856
rect 4178 800 4194 856
rect 4454 800 4470 856
rect 4822 800 4838 856
rect 5098 800 5114 856
rect 5466 800 5482 856
rect 5742 800 5758 856
rect 6110 800 6126 856
rect 6386 800 6402 856
rect 6662 800 6678 856
rect 7030 800 7046 856
rect 7306 800 7322 856
rect 7674 800 7690 856
rect 7950 800 7966 856
rect 8318 800 8334 856
rect 8594 800 8610 856
rect 8962 800 8978 856
rect 9238 800 9254 856
rect 9606 800 9622 856
rect 9882 800 9898 856
rect 10250 800 10266 856
rect 10526 800 10542 856
rect 10894 800 10910 856
rect 11170 800 11186 856
rect 11538 800 11554 856
rect 11814 800 11830 856
rect 12182 800 12198 856
rect 12458 800 12474 856
rect 12826 800 12842 856
rect 13102 800 13118 856
<< obsm3 >>
rect 565 987 13235 13089
<< metal4 >>
rect 2815 2128 3135 13104
rect 4685 2128 5005 13104
rect 6556 2128 6876 13104
rect 8427 2128 8747 13104
rect 10297 2128 10617 13104
<< obsm4 >>
rect 979 2048 2735 13104
rect 3215 2048 4605 13104
rect 5085 2048 6476 13104
rect 6956 2048 8347 13104
rect 8827 2048 10217 13104
rect 10697 2048 10981 13104
rect 979 987 10981 2048
<< metal5 >>
rect 1104 11035 12328 11355
rect 1104 9221 12328 9541
rect 1104 7408 12328 7728
rect 1104 5595 12328 5915
rect 1104 3781 12328 4101
<< obsm5 >>
rect 1104 9861 12328 10715
rect 1104 8048 12328 8901
rect 1104 6235 12328 7088
<< labels >>
rlabel metal2 s 11150 14818 11206 15618 6 cfg_bit_out
port 1 nsew signal output
rlabel metal2 s 12622 14818 12678 15618 6 cfg_bit_out_valid
port 2 nsew signal output
rlabel metal2 s 9678 14818 9734 15618 6 cfg_out_start
port 3 nsew signal output
rlabel metal2 s 3698 14818 3754 15618 6 col_sel[0]
port 4 nsew signal output
rlabel metal2 s 5170 14818 5226 15618 6 col_sel[1]
port 5 nsew signal output
rlabel metal2 s 6642 14818 6698 15618 6 col_sel[2]
port 6 nsew signal output
rlabel metal2 s 8206 14818 8262 15618 6 col_sel[3]
port 7 nsew signal output
rlabel metal2 s 754 14818 810 15618 6 wb_clk_i
port 8 nsew signal input
rlabel metal2 s 2226 14818 2282 15618 6 wb_rst_i
port 9 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_ack_o
port 10 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[0]
port 11 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[10]
port 12 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[11]
port 13 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[12]
port 14 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[13]
port 15 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[14]
port 16 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[15]
port 17 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[16]
port 18 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[17]
port 19 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[18]
port 20 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[19]
port 21 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[1]
port 22 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[20]
port 23 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[21]
port 24 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[22]
port 25 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[23]
port 26 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[24]
port 27 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[25]
port 28 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[26]
port 29 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[27]
port 30 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[28]
port 31 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[29]
port 32 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[2]
port 33 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[30]
port 34 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[31]
port 35 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[3]
port 36 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[4]
port 37 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[5]
port 38 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[6]
port 39 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[7]
port 40 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_adr_i[8]
port 41 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[9]
port 42 nsew signal input
rlabel metal2 s 110 0 166 800 6 wbs_cyc_i
port 43 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_dat_i[0]
port 44 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[10]
port 45 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[11]
port 46 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[12]
port 47 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[13]
port 48 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[14]
port 49 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[15]
port 50 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[16]
port 51 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[17]
port 52 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[18]
port 53 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[19]
port 54 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 55 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[20]
port 56 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[21]
port 57 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[22]
port 58 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[23]
port 59 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[24]
port 60 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[25]
port 61 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[26]
port 62 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[27]
port 63 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[28]
port 64 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[29]
port 65 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_dat_i[2]
port 66 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[30]
port 67 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[31]
port 68 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_dat_i[3]
port 69 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[4]
port 70 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[5]
port 71 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[6]
port 72 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[7]
port 73 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[8]
port 74 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_i[9]
port 75 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[0]
port 76 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[10]
port 77 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[11]
port 78 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[12]
port 79 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[13]
port 80 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 81 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[15]
port 82 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[16]
port 83 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[17]
port 84 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[18]
port 85 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[19]
port 86 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[1]
port 87 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[20]
port 88 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[21]
port 89 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[22]
port 90 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[23]
port 91 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[24]
port 92 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[25]
port 93 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[26]
port 94 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[27]
port 95 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[28]
port 96 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[29]
port 97 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[2]
port 98 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[30]
port 99 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[31]
port 100 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[3]
port 101 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[4]
port 102 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 103 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[6]
port 104 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[7]
port 105 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[8]
port 106 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[9]
port 107 nsew signal output
rlabel metal2 s 386 0 442 800 6 wbs_sel_i[0]
port 108 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_sel_i[1]
port 109 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_sel_i[2]
port 110 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_sel_i[3]
port 111 nsew signal input
rlabel metal2 s 18 0 74 800 6 wbs_stb_i
port 112 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_we_i
port 113 nsew signal input
rlabel metal4 s 10297 2128 10617 13104 6 VPWR
port 114 nsew power bidirectional
rlabel metal4 s 6556 2128 6876 13104 6 VPWR
port 115 nsew power bidirectional
rlabel metal4 s 2815 2128 3135 13104 6 VPWR
port 116 nsew power bidirectional
rlabel metal5 s 1104 11035 12328 11355 6 VPWR
port 117 nsew power bidirectional
rlabel metal5 s 1104 7408 12328 7728 6 VPWR
port 118 nsew power bidirectional
rlabel metal5 s 1104 3781 12328 4101 6 VPWR
port 119 nsew power bidirectional
rlabel metal4 s 8427 2128 8747 13104 6 VGND
port 120 nsew ground bidirectional
rlabel metal4 s 4685 2128 5005 13104 6 VGND
port 121 nsew ground bidirectional
rlabel metal5 s 1104 9221 12328 9541 6 VGND
port 122 nsew ground bidirectional
rlabel metal5 s 1104 5595 12328 5915 6 VGND
port 123 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 13474 15618
string LEFview TRUE
string GDS_FILE /tools/B/tan.nqd/fabric_team/asic_config/wb_config/runs/12-06_19-45/results/magic/wb_config.gds
string GDS_END 1012174
string GDS_START 182316
<< end >>

