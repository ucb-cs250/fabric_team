VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block_east
  CLASS BLOCK ;
  FOREIGN baked_connection_block_east ;
  ORIGIN 0.000 0.000 ;
  SIZE 254.225 BY 264.945 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 6.840 254.225 7.440 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 20.440 254.225 21.040 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 34.720 254.225 35.320 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 48.320 254.225 48.920 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 62.600 254.225 63.200 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 76.200 254.225 76.800 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 90.480 254.225 91.080 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 104.080 254.225 104.680 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 118.360 254.225 118.960 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 131.960 254.225 132.560 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 146.240 254.225 146.840 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 159.840 254.225 160.440 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 174.120 254.225 174.720 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 187.720 254.225 188.320 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 202.000 254.225 202.600 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 215.600 254.225 216.200 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 229.880 254.225 230.480 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.870 260.945 227.150 264.945 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 260.945 81.790 264.945 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 260.945 99.730 264.945 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 260.945 118.130 264.945 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 260.945 136.070 264.945 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 260.945 154.470 264.945 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 260.945 172.410 264.945 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 260.945 190.810 264.945 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.470 260.945 208.750 264.945 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END double1[7]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.810 260.945 245.090 264.945 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 243.480 254.225 244.080 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 257.760 254.225 258.360 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 260.945 9.110 264.945 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 260.945 27.050 264.945 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 260.945 45.450 264.945 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 260.945 63.390 264.945 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 253.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 253.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 248.400 253.045 ;
      LAYER met1 ;
        RECT 5.520 4.460 248.400 260.740 ;
      LAYER met2 ;
        RECT 7.460 260.665 8.550 260.945 ;
        RECT 9.390 260.665 26.490 260.945 ;
        RECT 27.330 260.665 44.890 260.945 ;
        RECT 45.730 260.665 62.830 260.945 ;
        RECT 63.670 260.665 81.230 260.945 ;
        RECT 82.070 260.665 99.170 260.945 ;
        RECT 100.010 260.665 117.570 260.945 ;
        RECT 118.410 260.665 135.510 260.945 ;
        RECT 136.350 260.665 153.910 260.945 ;
        RECT 154.750 260.665 171.850 260.945 ;
        RECT 172.690 260.665 190.250 260.945 ;
        RECT 191.090 260.665 208.190 260.945 ;
        RECT 209.030 260.665 226.590 260.945 ;
        RECT 227.430 260.665 244.530 260.945 ;
        RECT 7.460 4.280 245.080 260.665 ;
        RECT 7.460 4.000 9.470 4.280 ;
        RECT 10.310 4.000 28.790 4.280 ;
        RECT 29.630 4.000 48.570 4.280 ;
        RECT 49.410 4.000 67.890 4.280 ;
        RECT 68.730 4.000 87.670 4.280 ;
        RECT 88.510 4.000 106.990 4.280 ;
        RECT 107.830 4.000 126.770 4.280 ;
        RECT 127.610 4.000 146.090 4.280 ;
        RECT 146.930 4.000 165.870 4.280 ;
        RECT 166.710 4.000 185.190 4.280 ;
        RECT 186.030 4.000 204.970 4.280 ;
        RECT 205.810 4.000 224.290 4.280 ;
        RECT 225.130 4.000 244.070 4.280 ;
        RECT 244.910 4.000 245.080 4.280 ;
      LAYER met3 ;
        RECT 4.000 258.080 249.825 258.225 ;
        RECT 4.400 257.360 249.825 258.080 ;
        RECT 4.400 256.680 250.225 257.360 ;
        RECT 4.000 244.480 250.225 256.680 ;
        RECT 4.000 243.120 249.825 244.480 ;
        RECT 4.400 243.080 249.825 243.120 ;
        RECT 4.400 241.720 250.225 243.080 ;
        RECT 4.000 230.880 250.225 241.720 ;
        RECT 4.000 229.480 249.825 230.880 ;
        RECT 4.000 228.840 250.225 229.480 ;
        RECT 4.400 227.440 250.225 228.840 ;
        RECT 4.000 216.600 250.225 227.440 ;
        RECT 4.000 215.200 249.825 216.600 ;
        RECT 4.000 213.880 250.225 215.200 ;
        RECT 4.400 212.480 250.225 213.880 ;
        RECT 4.000 203.000 250.225 212.480 ;
        RECT 4.000 201.600 249.825 203.000 ;
        RECT 4.000 198.920 250.225 201.600 ;
        RECT 4.400 197.520 250.225 198.920 ;
        RECT 4.000 188.720 250.225 197.520 ;
        RECT 4.000 187.320 249.825 188.720 ;
        RECT 4.000 184.640 250.225 187.320 ;
        RECT 4.400 183.240 250.225 184.640 ;
        RECT 4.000 175.120 250.225 183.240 ;
        RECT 4.000 173.720 249.825 175.120 ;
        RECT 4.000 169.680 250.225 173.720 ;
        RECT 4.400 168.280 250.225 169.680 ;
        RECT 4.000 160.840 250.225 168.280 ;
        RECT 4.000 159.440 249.825 160.840 ;
        RECT 4.000 154.720 250.225 159.440 ;
        RECT 4.400 153.320 250.225 154.720 ;
        RECT 4.000 147.240 250.225 153.320 ;
        RECT 4.000 145.840 249.825 147.240 ;
        RECT 4.000 140.440 250.225 145.840 ;
        RECT 4.400 139.040 250.225 140.440 ;
        RECT 4.000 132.960 250.225 139.040 ;
        RECT 4.000 131.560 249.825 132.960 ;
        RECT 4.000 125.480 250.225 131.560 ;
        RECT 4.400 124.080 250.225 125.480 ;
        RECT 4.000 119.360 250.225 124.080 ;
        RECT 4.000 117.960 249.825 119.360 ;
        RECT 4.000 110.520 250.225 117.960 ;
        RECT 4.400 109.120 250.225 110.520 ;
        RECT 4.000 105.080 250.225 109.120 ;
        RECT 4.000 103.680 249.825 105.080 ;
        RECT 4.000 96.240 250.225 103.680 ;
        RECT 4.400 94.840 250.225 96.240 ;
        RECT 4.000 91.480 250.225 94.840 ;
        RECT 4.000 90.080 249.825 91.480 ;
        RECT 4.000 81.280 250.225 90.080 ;
        RECT 4.400 79.880 250.225 81.280 ;
        RECT 4.000 77.200 250.225 79.880 ;
        RECT 4.000 75.800 249.825 77.200 ;
        RECT 4.000 66.320 250.225 75.800 ;
        RECT 4.400 64.920 250.225 66.320 ;
        RECT 4.000 63.600 250.225 64.920 ;
        RECT 4.000 62.200 249.825 63.600 ;
        RECT 4.000 52.040 250.225 62.200 ;
        RECT 4.400 50.640 250.225 52.040 ;
        RECT 4.000 49.320 250.225 50.640 ;
        RECT 4.000 47.920 249.825 49.320 ;
        RECT 4.000 37.080 250.225 47.920 ;
        RECT 4.400 35.720 250.225 37.080 ;
        RECT 4.400 35.680 249.825 35.720 ;
        RECT 4.000 34.320 249.825 35.680 ;
        RECT 4.000 22.120 250.225 34.320 ;
        RECT 4.400 21.440 250.225 22.120 ;
        RECT 4.400 20.720 249.825 21.440 ;
        RECT 4.000 20.040 249.825 20.720 ;
        RECT 4.000 7.840 250.225 20.040 ;
        RECT 4.400 6.975 249.825 7.840 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 253.200 ;
  END
END baked_connection_block_east
END LIBRARY

