VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 260.700 BY 271.420 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 267.420 242.330 271.420 ;
    END
  END COUT
  PIN cb_e_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 2.760 260.700 3.360 ;
    END
  END cb_e_clb1_input[0]
  PIN cb_e_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 8.200 260.700 8.800 ;
    END
  END cb_e_clb1_input[1]
  PIN cb_e_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 14.320 260.700 14.920 ;
    END
  END cb_e_clb1_input[2]
  PIN cb_e_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 20.440 260.700 21.040 ;
    END
  END cb_e_clb1_input[3]
  PIN cb_e_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 25.880 260.700 26.480 ;
    END
  END cb_e_clb1_input[4]
  PIN cb_e_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 32.000 260.700 32.600 ;
    END
  END cb_e_clb1_input[5]
  PIN cb_e_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 38.120 260.700 38.720 ;
    END
  END cb_e_clb1_input[6]
  PIN cb_e_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 43.560 260.700 44.160 ;
    END
  END cb_e_clb1_input[7]
  PIN cb_e_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 49.680 260.700 50.280 ;
    END
  END cb_e_clb1_input[8]
  PIN cb_e_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 55.800 260.700 56.400 ;
    END
  END cb_e_clb1_input[9]
  PIN cb_e_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 61.240 260.700 61.840 ;
    END
  END cb_e_clb1_output[0]
  PIN cb_e_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 67.360 260.700 67.960 ;
    END
  END cb_e_clb1_output[1]
  PIN cb_e_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 73.480 260.700 74.080 ;
    END
  END cb_e_clb1_output[2]
  PIN cb_e_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 78.920 260.700 79.520 ;
    END
  END cb_e_clb1_output[3]
  PIN cb_e_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END cb_e_single1_in[0]
  PIN cb_e_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END cb_e_single1_in[10]
  PIN cb_e_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END cb_e_single1_in[11]
  PIN cb_e_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cb_e_single1_in[12]
  PIN cb_e_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END cb_e_single1_in[13]
  PIN cb_e_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END cb_e_single1_in[14]
  PIN cb_e_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END cb_e_single1_in[15]
  PIN cb_e_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END cb_e_single1_in[1]
  PIN cb_e_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END cb_e_single1_in[2]
  PIN cb_e_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END cb_e_single1_in[3]
  PIN cb_e_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END cb_e_single1_in[4]
  PIN cb_e_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END cb_e_single1_in[5]
  PIN cb_e_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END cb_e_single1_in[6]
  PIN cb_e_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END cb_e_single1_in[7]
  PIN cb_e_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END cb_e_single1_in[8]
  PIN cb_e_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END cb_e_single1_in[9]
  PIN cb_e_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END cb_e_single1_out[0]
  PIN cb_e_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END cb_e_single1_out[10]
  PIN cb_e_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END cb_e_single1_out[11]
  PIN cb_e_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END cb_e_single1_out[12]
  PIN cb_e_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END cb_e_single1_out[13]
  PIN cb_e_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END cb_e_single1_out[14]
  PIN cb_e_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END cb_e_single1_out[15]
  PIN cb_e_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END cb_e_single1_out[1]
  PIN cb_e_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END cb_e_single1_out[2]
  PIN cb_e_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cb_e_single1_out[3]
  PIN cb_e_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cb_e_single1_out[4]
  PIN cb_e_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END cb_e_single1_out[5]
  PIN cb_e_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END cb_e_single1_out[6]
  PIN cb_e_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cb_e_single1_out[7]
  PIN cb_e_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END cb_e_single1_out[8]
  PIN cb_e_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END cb_e_single1_out[9]
  PIN cb_n_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 267.420 2.670 271.420 ;
    END
  END cb_n_clb1_input[0]
  PIN cb_n_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 267.420 7.730 271.420 ;
    END
  END cb_n_clb1_input[1]
  PIN cb_n_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 267.420 12.790 271.420 ;
    END
  END cb_n_clb1_input[2]
  PIN cb_n_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 267.420 18.310 271.420 ;
    END
  END cb_n_clb1_input[3]
  PIN cb_n_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 267.420 23.370 271.420 ;
    END
  END cb_n_clb1_input[4]
  PIN cb_n_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 267.420 28.430 271.420 ;
    END
  END cb_n_clb1_input[5]
  PIN cb_n_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 267.420 33.950 271.420 ;
    END
  END cb_n_clb1_input[6]
  PIN cb_n_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 267.420 39.010 271.420 ;
    END
  END cb_n_clb1_input[7]
  PIN cb_n_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 267.420 44.070 271.420 ;
    END
  END cb_n_clb1_input[8]
  PIN cb_n_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 267.420 49.590 271.420 ;
    END
  END cb_n_clb1_input[9]
  PIN cb_n_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 267.420 54.650 271.420 ;
    END
  END cb_n_clb1_output[0]
  PIN cb_n_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 267.420 59.710 271.420 ;
    END
  END cb_n_clb1_output[1]
  PIN cb_n_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 267.420 65.230 271.420 ;
    END
  END cb_n_clb1_output[2]
  PIN cb_n_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 267.420 70.290 271.420 ;
    END
  END cb_n_clb1_output[3]
  PIN cb_n_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END cb_n_single1_in[0]
  PIN cb_n_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END cb_n_single1_in[10]
  PIN cb_n_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END cb_n_single1_in[11]
  PIN cb_n_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END cb_n_single1_in[12]
  PIN cb_n_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END cb_n_single1_in[13]
  PIN cb_n_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END cb_n_single1_in[14]
  PIN cb_n_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END cb_n_single1_in[15]
  PIN cb_n_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END cb_n_single1_in[1]
  PIN cb_n_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END cb_n_single1_in[2]
  PIN cb_n_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END cb_n_single1_in[3]
  PIN cb_n_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END cb_n_single1_in[4]
  PIN cb_n_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END cb_n_single1_in[5]
  PIN cb_n_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END cb_n_single1_in[6]
  PIN cb_n_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END cb_n_single1_in[7]
  PIN cb_n_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END cb_n_single1_in[8]
  PIN cb_n_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END cb_n_single1_in[9]
  PIN cb_n_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END cb_n_single1_out[0]
  PIN cb_n_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END cb_n_single1_out[10]
  PIN cb_n_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END cb_n_single1_out[11]
  PIN cb_n_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END cb_n_single1_out[12]
  PIN cb_n_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END cb_n_single1_out[13]
  PIN cb_n_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END cb_n_single1_out[14]
  PIN cb_n_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END cb_n_single1_out[15]
  PIN cb_n_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END cb_n_single1_out[1]
  PIN cb_n_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END cb_n_single1_out[2]
  PIN cb_n_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END cb_n_single1_out[3]
  PIN cb_n_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END cb_n_single1_out[4]
  PIN cb_n_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END cb_n_single1_out[5]
  PIN cb_n_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END cb_n_single1_out[6]
  PIN cb_n_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END cb_n_single1_out[7]
  PIN cb_n_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END cb_n_single1_out[8]
  PIN cb_n_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END cb_n_single1_out[9]
  PIN cfg_bit_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END cfg_bit_in
  PIN cfg_bit_in_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END cfg_bit_in_valid
  PIN cfg_bit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 267.420 252.910 271.420 ;
    END
  END cfg_bit_out
  PIN cfg_bit_out_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 267.420 257.970 271.420 ;
    END
  END cfg_bit_out_valid
  PIN cfg_in_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END cfg_in_start
  PIN cfg_out_start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 267.420 247.390 271.420 ;
    END
  END cfg_out_start
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END clb_south_out[3]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END clb_west_out[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END clk
  PIN crst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END crst
  PIN sb_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 85.040 260.700 85.640 ;
    END
  END sb_east_in[0]
  PIN sb_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 144.200 260.700 144.800 ;
    END
  END sb_east_in[10]
  PIN sb_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 149.640 260.700 150.240 ;
    END
  END sb_east_in[11]
  PIN sb_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 155.760 260.700 156.360 ;
    END
  END sb_east_in[12]
  PIN sb_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 161.880 260.700 162.480 ;
    END
  END sb_east_in[13]
  PIN sb_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 167.320 260.700 167.920 ;
    END
  END sb_east_in[14]
  PIN sb_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 173.440 260.700 174.040 ;
    END
  END sb_east_in[15]
  PIN sb_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 91.160 260.700 91.760 ;
    END
  END sb_east_in[1]
  PIN sb_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 96.600 260.700 97.200 ;
    END
  END sb_east_in[2]
  PIN sb_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 102.720 260.700 103.320 ;
    END
  END sb_east_in[3]
  PIN sb_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 108.840 260.700 109.440 ;
    END
  END sb_east_in[4]
  PIN sb_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 114.280 260.700 114.880 ;
    END
  END sb_east_in[5]
  PIN sb_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 120.400 260.700 121.000 ;
    END
  END sb_east_in[6]
  PIN sb_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 126.520 260.700 127.120 ;
    END
  END sb_east_in[7]
  PIN sb_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 131.960 260.700 132.560 ;
    END
  END sb_east_in[8]
  PIN sb_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 138.080 260.700 138.680 ;
    END
  END sb_east_in[9]
  PIN sb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 179.560 260.700 180.160 ;
    END
  END sb_east_out[0]
  PIN sb_east_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 238.040 260.700 238.640 ;
    END
  END sb_east_out[10]
  PIN sb_east_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 244.160 260.700 244.760 ;
    END
  END sb_east_out[11]
  PIN sb_east_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 250.280 260.700 250.880 ;
    END
  END sb_east_out[12]
  PIN sb_east_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 255.720 260.700 256.320 ;
    END
  END sb_east_out[13]
  PIN sb_east_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 261.840 260.700 262.440 ;
    END
  END sb_east_out[14]
  PIN sb_east_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 267.960 260.700 268.560 ;
    END
  END sb_east_out[15]
  PIN sb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 185.000 260.700 185.600 ;
    END
  END sb_east_out[1]
  PIN sb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 191.120 260.700 191.720 ;
    END
  END sb_east_out[2]
  PIN sb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 197.240 260.700 197.840 ;
    END
  END sb_east_out[3]
  PIN sb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 202.680 260.700 203.280 ;
    END
  END sb_east_out[4]
  PIN sb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 208.800 260.700 209.400 ;
    END
  END sb_east_out[5]
  PIN sb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 214.920 260.700 215.520 ;
    END
  END sb_east_out[6]
  PIN sb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 220.360 260.700 220.960 ;
    END
  END sb_east_out[7]
  PIN sb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 226.480 260.700 227.080 ;
    END
  END sb_east_out[8]
  PIN sb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.700 232.600 260.700 233.200 ;
    END
  END sb_east_out[9]
  PIN sb_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 267.420 75.350 271.420 ;
    END
  END sb_north_in[0]
  PIN sb_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 267.420 127.790 271.420 ;
    END
  END sb_north_in[10]
  PIN sb_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 267.420 132.850 271.420 ;
    END
  END sb_north_in[11]
  PIN sb_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 267.420 137.910 271.420 ;
    END
  END sb_north_in[12]
  PIN sb_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 267.420 143.430 271.420 ;
    END
  END sb_north_in[13]
  PIN sb_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 267.420 148.490 271.420 ;
    END
  END sb_north_in[14]
  PIN sb_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 267.420 153.550 271.420 ;
    END
  END sb_north_in[15]
  PIN sb_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 267.420 80.870 271.420 ;
    END
  END sb_north_in[1]
  PIN sb_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 267.420 85.930 271.420 ;
    END
  END sb_north_in[2]
  PIN sb_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 267.420 90.990 271.420 ;
    END
  END sb_north_in[3]
  PIN sb_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 267.420 96.510 271.420 ;
    END
  END sb_north_in[4]
  PIN sb_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 267.420 101.570 271.420 ;
    END
  END sb_north_in[5]
  PIN sb_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 267.420 106.630 271.420 ;
    END
  END sb_north_in[6]
  PIN sb_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 267.420 112.150 271.420 ;
    END
  END sb_north_in[7]
  PIN sb_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 267.420 117.210 271.420 ;
    END
  END sb_north_in[8]
  PIN sb_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 267.420 122.270 271.420 ;
    END
  END sb_north_in[9]
  PIN sb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 267.420 159.070 271.420 ;
    END
  END sb_north_out[0]
  PIN sb_north_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 267.420 211.050 271.420 ;
    END
  END sb_north_out[10]
  PIN sb_north_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 267.420 216.110 271.420 ;
    END
  END sb_north_out[11]
  PIN sb_north_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 267.420 221.630 271.420 ;
    END
  END sb_north_out[12]
  PIN sb_north_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 267.420 226.690 271.420 ;
    END
  END sb_north_out[13]
  PIN sb_north_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 267.420 231.750 271.420 ;
    END
  END sb_north_out[14]
  PIN sb_north_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 267.420 237.270 271.420 ;
    END
  END sb_north_out[15]
  PIN sb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 267.420 164.130 271.420 ;
    END
  END sb_north_out[1]
  PIN sb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 267.420 169.190 271.420 ;
    END
  END sb_north_out[2]
  PIN sb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 267.420 174.710 271.420 ;
    END
  END sb_north_out[3]
  PIN sb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 267.420 179.770 271.420 ;
    END
  END sb_north_out[4]
  PIN sb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 267.420 184.830 271.420 ;
    END
  END sb_north_out[5]
  PIN sb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 267.420 190.350 271.420 ;
    END
  END sb_north_out[6]
  PIN sb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 267.420 195.410 271.420 ;
    END
  END sb_north_out[7]
  PIN sb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 267.420 200.470 271.420 ;
    END
  END sb_north_out[8]
  PIN sb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 267.420 205.990 271.420 ;
    END
  END sb_north_out[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 258.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 258.640 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 258.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 258.640 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 7.225 256.075 258.485 ;
      LAYER met1 ;
        RECT 2.370 213.820 260.700 262.100 ;
        RECT 2.370 213.560 260.750 213.820 ;
        RECT 2.370 6.500 260.700 213.560 ;
      LAYER met2 ;
        RECT 2.950 267.140 7.170 268.445 ;
        RECT 8.010 267.140 12.230 268.445 ;
        RECT 13.070 267.140 17.750 268.445 ;
        RECT 18.590 267.140 22.810 268.445 ;
        RECT 23.650 267.140 27.870 268.445 ;
        RECT 28.710 267.140 33.390 268.445 ;
        RECT 34.230 267.140 38.450 268.445 ;
        RECT 39.290 267.140 43.510 268.445 ;
        RECT 44.350 267.140 49.030 268.445 ;
        RECT 49.870 267.140 54.090 268.445 ;
        RECT 54.930 267.140 59.150 268.445 ;
        RECT 59.990 267.140 64.670 268.445 ;
        RECT 65.510 267.140 69.730 268.445 ;
        RECT 70.570 267.140 74.790 268.445 ;
        RECT 75.630 267.140 80.310 268.445 ;
        RECT 81.150 267.140 85.370 268.445 ;
        RECT 86.210 267.140 90.430 268.445 ;
        RECT 91.270 267.140 95.950 268.445 ;
        RECT 96.790 267.140 101.010 268.445 ;
        RECT 101.850 267.140 106.070 268.445 ;
        RECT 106.910 267.140 111.590 268.445 ;
        RECT 112.430 267.140 116.650 268.445 ;
        RECT 117.490 267.140 121.710 268.445 ;
        RECT 122.550 267.140 127.230 268.445 ;
        RECT 128.070 267.140 132.290 268.445 ;
        RECT 133.130 267.140 137.350 268.445 ;
        RECT 138.190 267.140 142.870 268.445 ;
        RECT 143.710 267.140 147.930 268.445 ;
        RECT 148.770 267.140 152.990 268.445 ;
        RECT 153.830 267.140 158.510 268.445 ;
        RECT 159.350 267.140 163.570 268.445 ;
        RECT 164.410 267.140 168.630 268.445 ;
        RECT 169.470 267.140 174.150 268.445 ;
        RECT 174.990 267.140 179.210 268.445 ;
        RECT 180.050 267.140 184.270 268.445 ;
        RECT 185.110 267.140 189.790 268.445 ;
        RECT 190.630 267.140 194.850 268.445 ;
        RECT 195.690 267.140 199.910 268.445 ;
        RECT 200.750 267.140 205.430 268.445 ;
        RECT 206.270 267.140 210.490 268.445 ;
        RECT 211.330 267.140 215.550 268.445 ;
        RECT 216.390 267.140 221.070 268.445 ;
        RECT 221.910 267.140 226.130 268.445 ;
        RECT 226.970 267.140 231.190 268.445 ;
        RECT 232.030 267.140 236.710 268.445 ;
        RECT 237.550 267.140 241.770 268.445 ;
        RECT 242.610 267.140 246.830 268.445 ;
        RECT 247.670 267.140 252.350 268.445 ;
        RECT 253.190 267.140 257.410 268.445 ;
        RECT 258.250 267.140 260.700 268.445 ;
        RECT 2.400 213.850 260.700 267.140 ;
        RECT 2.400 213.530 260.720 213.850 ;
        RECT 2.400 124.285 260.700 213.530 ;
        RECT 2.400 123.915 260.730 124.285 ;
        RECT 2.400 4.280 260.700 123.915 ;
        RECT 2.950 2.875 7.170 4.280 ;
        RECT 8.010 2.875 12.230 4.280 ;
        RECT 13.070 2.875 17.290 4.280 ;
        RECT 18.130 2.875 22.350 4.280 ;
        RECT 23.190 2.875 27.410 4.280 ;
        RECT 28.250 2.875 32.470 4.280 ;
        RECT 33.310 2.875 37.530 4.280 ;
        RECT 38.370 2.875 42.590 4.280 ;
        RECT 43.430 2.875 48.110 4.280 ;
        RECT 48.950 2.875 53.170 4.280 ;
        RECT 54.010 2.875 58.230 4.280 ;
        RECT 59.070 2.875 63.290 4.280 ;
        RECT 64.130 2.875 68.350 4.280 ;
        RECT 69.190 2.875 73.410 4.280 ;
        RECT 74.250 2.875 78.470 4.280 ;
        RECT 79.310 2.875 83.530 4.280 ;
        RECT 84.370 2.875 89.050 4.280 ;
        RECT 89.890 2.875 94.110 4.280 ;
        RECT 94.950 2.875 99.170 4.280 ;
        RECT 100.010 2.875 104.230 4.280 ;
        RECT 105.070 2.875 109.290 4.280 ;
        RECT 110.130 2.875 114.350 4.280 ;
        RECT 115.190 2.875 119.410 4.280 ;
        RECT 120.250 2.875 124.470 4.280 ;
        RECT 125.310 2.875 129.530 4.280 ;
        RECT 130.370 2.875 135.050 4.280 ;
        RECT 135.890 2.875 140.110 4.280 ;
        RECT 140.950 2.875 145.170 4.280 ;
        RECT 146.010 2.875 150.230 4.280 ;
        RECT 151.070 2.875 155.290 4.280 ;
        RECT 156.130 2.875 160.350 4.280 ;
        RECT 161.190 2.875 165.410 4.280 ;
        RECT 166.250 2.875 170.470 4.280 ;
        RECT 171.310 2.875 175.990 4.280 ;
        RECT 176.830 2.875 181.050 4.280 ;
        RECT 181.890 2.875 186.110 4.280 ;
        RECT 186.950 2.875 191.170 4.280 ;
        RECT 192.010 2.875 196.230 4.280 ;
        RECT 197.070 2.875 201.290 4.280 ;
        RECT 202.130 2.875 206.350 4.280 ;
        RECT 207.190 2.875 211.410 4.280 ;
        RECT 212.250 2.875 216.470 4.280 ;
        RECT 217.310 2.875 221.990 4.280 ;
        RECT 222.830 2.875 227.050 4.280 ;
        RECT 227.890 2.875 232.110 4.280 ;
        RECT 232.950 2.875 237.170 4.280 ;
        RECT 238.010 2.875 242.230 4.280 ;
        RECT 243.070 2.875 247.290 4.280 ;
        RECT 248.130 2.875 252.350 4.280 ;
        RECT 253.190 2.875 257.410 4.280 ;
        RECT 258.250 2.875 260.700 4.280 ;
      LAYER met3 ;
        RECT 4.400 267.560 256.300 268.425 ;
        RECT 4.000 263.520 260.700 267.560 ;
        RECT 4.400 262.840 260.700 263.520 ;
        RECT 4.400 262.120 256.300 262.840 ;
        RECT 4.000 261.440 256.300 262.120 ;
        RECT 4.000 257.400 260.700 261.440 ;
        RECT 4.400 256.720 260.700 257.400 ;
        RECT 4.400 256.000 256.300 256.720 ;
        RECT 4.000 255.320 256.300 256.000 ;
        RECT 4.000 251.960 260.700 255.320 ;
        RECT 4.400 251.280 260.700 251.960 ;
        RECT 4.400 250.560 256.300 251.280 ;
        RECT 4.000 249.880 256.300 250.560 ;
        RECT 4.000 245.840 260.700 249.880 ;
        RECT 4.400 245.160 260.700 245.840 ;
        RECT 4.400 244.440 256.300 245.160 ;
        RECT 4.000 243.760 256.300 244.440 ;
        RECT 4.000 240.400 260.700 243.760 ;
        RECT 4.400 239.040 260.700 240.400 ;
        RECT 4.400 239.000 256.300 239.040 ;
        RECT 4.000 237.640 256.300 239.000 ;
        RECT 4.000 234.280 260.700 237.640 ;
        RECT 4.400 233.600 260.700 234.280 ;
        RECT 4.400 232.880 256.300 233.600 ;
        RECT 4.000 232.200 256.300 232.880 ;
        RECT 4.000 228.840 260.700 232.200 ;
        RECT 4.400 227.480 260.700 228.840 ;
        RECT 4.400 227.440 256.300 227.480 ;
        RECT 4.000 226.080 256.300 227.440 ;
        RECT 4.000 222.720 260.700 226.080 ;
        RECT 4.400 221.360 260.700 222.720 ;
        RECT 4.400 221.320 256.300 221.360 ;
        RECT 4.000 219.960 256.300 221.320 ;
        RECT 4.000 217.280 260.700 219.960 ;
        RECT 4.400 215.920 260.700 217.280 ;
        RECT 4.400 215.880 256.300 215.920 ;
        RECT 4.000 214.520 256.300 215.880 ;
        RECT 4.000 211.160 260.700 214.520 ;
        RECT 4.400 209.800 260.700 211.160 ;
        RECT 4.400 209.760 256.300 209.800 ;
        RECT 4.000 208.400 256.300 209.760 ;
        RECT 4.000 205.720 260.700 208.400 ;
        RECT 4.400 204.320 260.700 205.720 ;
        RECT 4.000 203.680 260.700 204.320 ;
        RECT 4.000 202.280 256.300 203.680 ;
        RECT 4.000 199.600 260.700 202.280 ;
        RECT 4.400 198.240 260.700 199.600 ;
        RECT 4.400 198.200 256.300 198.240 ;
        RECT 4.000 196.840 256.300 198.200 ;
        RECT 4.000 194.160 260.700 196.840 ;
        RECT 4.400 192.760 260.700 194.160 ;
        RECT 4.000 192.120 260.700 192.760 ;
        RECT 4.000 190.720 256.300 192.120 ;
        RECT 4.000 188.040 260.700 190.720 ;
        RECT 4.400 186.640 260.700 188.040 ;
        RECT 4.000 186.000 260.700 186.640 ;
        RECT 4.000 184.600 256.300 186.000 ;
        RECT 4.000 182.600 260.700 184.600 ;
        RECT 4.400 181.200 260.700 182.600 ;
        RECT 4.000 180.560 260.700 181.200 ;
        RECT 4.000 179.160 256.300 180.560 ;
        RECT 4.000 176.480 260.700 179.160 ;
        RECT 4.400 175.080 260.700 176.480 ;
        RECT 4.000 174.440 260.700 175.080 ;
        RECT 4.000 173.040 256.300 174.440 ;
        RECT 4.000 171.040 260.700 173.040 ;
        RECT 4.400 169.640 260.700 171.040 ;
        RECT 4.000 168.320 260.700 169.640 ;
        RECT 4.000 166.920 256.300 168.320 ;
        RECT 4.000 164.920 260.700 166.920 ;
        RECT 4.400 163.520 260.700 164.920 ;
        RECT 4.000 162.880 260.700 163.520 ;
        RECT 4.000 161.480 256.300 162.880 ;
        RECT 4.000 159.480 260.700 161.480 ;
        RECT 4.400 158.080 260.700 159.480 ;
        RECT 4.000 156.760 260.700 158.080 ;
        RECT 4.000 155.360 256.300 156.760 ;
        RECT 4.000 153.360 260.700 155.360 ;
        RECT 4.400 151.960 260.700 153.360 ;
        RECT 4.000 150.640 260.700 151.960 ;
        RECT 4.000 149.240 256.300 150.640 ;
        RECT 4.000 147.920 260.700 149.240 ;
        RECT 4.400 146.520 260.700 147.920 ;
        RECT 4.000 145.200 260.700 146.520 ;
        RECT 4.000 143.800 256.300 145.200 ;
        RECT 4.000 141.800 260.700 143.800 ;
        RECT 4.400 140.400 260.700 141.800 ;
        RECT 4.000 139.080 260.700 140.400 ;
        RECT 4.000 137.680 256.300 139.080 ;
        RECT 4.000 136.360 260.700 137.680 ;
        RECT 4.400 134.960 260.700 136.360 ;
        RECT 4.000 132.960 260.700 134.960 ;
        RECT 4.000 131.560 256.300 132.960 ;
        RECT 4.000 130.240 260.700 131.560 ;
        RECT 4.400 128.840 260.700 130.240 ;
        RECT 4.000 127.520 260.700 128.840 ;
        RECT 4.000 126.120 256.300 127.520 ;
        RECT 4.000 124.800 260.700 126.120 ;
        RECT 4.400 124.265 260.700 124.800 ;
        RECT 4.400 123.935 260.755 124.265 ;
        RECT 4.400 123.400 260.700 123.935 ;
        RECT 4.000 121.400 260.700 123.400 ;
        RECT 4.000 120.000 256.300 121.400 ;
        RECT 4.000 118.680 260.700 120.000 ;
        RECT 4.400 117.280 260.700 118.680 ;
        RECT 4.000 115.280 260.700 117.280 ;
        RECT 4.000 113.880 256.300 115.280 ;
        RECT 4.000 113.240 260.700 113.880 ;
        RECT 4.400 111.840 260.700 113.240 ;
        RECT 4.000 109.840 260.700 111.840 ;
        RECT 4.000 108.440 256.300 109.840 ;
        RECT 4.000 107.120 260.700 108.440 ;
        RECT 4.400 105.720 260.700 107.120 ;
        RECT 4.000 103.720 260.700 105.720 ;
        RECT 4.000 102.320 256.300 103.720 ;
        RECT 4.000 101.680 260.700 102.320 ;
        RECT 4.400 100.280 260.700 101.680 ;
        RECT 4.000 97.600 260.700 100.280 ;
        RECT 4.000 96.200 256.300 97.600 ;
        RECT 4.000 95.560 260.700 96.200 ;
        RECT 4.400 94.160 260.700 95.560 ;
        RECT 4.000 92.160 260.700 94.160 ;
        RECT 4.000 90.760 256.300 92.160 ;
        RECT 4.000 90.120 260.700 90.760 ;
        RECT 4.400 88.720 260.700 90.120 ;
        RECT 4.000 86.040 260.700 88.720 ;
        RECT 4.000 84.640 256.300 86.040 ;
        RECT 4.000 84.000 260.700 84.640 ;
        RECT 4.400 82.600 260.700 84.000 ;
        RECT 4.000 79.920 260.700 82.600 ;
        RECT 4.000 78.560 256.300 79.920 ;
        RECT 4.400 78.520 256.300 78.560 ;
        RECT 4.400 77.160 260.700 78.520 ;
        RECT 4.000 74.480 260.700 77.160 ;
        RECT 4.000 73.080 256.300 74.480 ;
        RECT 4.000 72.440 260.700 73.080 ;
        RECT 4.400 71.040 260.700 72.440 ;
        RECT 4.000 68.360 260.700 71.040 ;
        RECT 4.000 67.000 256.300 68.360 ;
        RECT 4.400 66.960 256.300 67.000 ;
        RECT 4.400 65.600 260.700 66.960 ;
        RECT 4.000 62.240 260.700 65.600 ;
        RECT 4.000 60.880 256.300 62.240 ;
        RECT 4.400 60.840 256.300 60.880 ;
        RECT 4.400 59.480 260.700 60.840 ;
        RECT 4.000 56.800 260.700 59.480 ;
        RECT 4.000 55.440 256.300 56.800 ;
        RECT 4.400 55.400 256.300 55.440 ;
        RECT 4.400 54.040 260.700 55.400 ;
        RECT 4.000 50.680 260.700 54.040 ;
        RECT 4.000 49.320 256.300 50.680 ;
        RECT 4.400 49.280 256.300 49.320 ;
        RECT 4.400 47.920 260.700 49.280 ;
        RECT 4.000 44.560 260.700 47.920 ;
        RECT 4.000 43.880 256.300 44.560 ;
        RECT 4.400 43.160 256.300 43.880 ;
        RECT 4.400 42.480 260.700 43.160 ;
        RECT 4.000 39.120 260.700 42.480 ;
        RECT 4.000 37.760 256.300 39.120 ;
        RECT 4.400 37.720 256.300 37.760 ;
        RECT 4.400 36.360 260.700 37.720 ;
        RECT 4.000 33.000 260.700 36.360 ;
        RECT 4.000 32.320 256.300 33.000 ;
        RECT 4.400 31.600 256.300 32.320 ;
        RECT 4.400 30.920 260.700 31.600 ;
        RECT 4.000 26.880 260.700 30.920 ;
        RECT 4.000 26.200 256.300 26.880 ;
        RECT 4.400 25.480 256.300 26.200 ;
        RECT 4.400 24.800 260.700 25.480 ;
        RECT 4.000 21.440 260.700 24.800 ;
        RECT 4.000 20.760 256.300 21.440 ;
        RECT 4.400 20.040 256.300 20.760 ;
        RECT 4.400 19.360 260.700 20.040 ;
        RECT 4.000 15.320 260.700 19.360 ;
        RECT 4.000 14.640 256.300 15.320 ;
        RECT 4.400 13.920 256.300 14.640 ;
        RECT 4.400 13.240 260.700 13.920 ;
        RECT 4.000 9.200 260.700 13.240 ;
        RECT 4.400 7.800 256.300 9.200 ;
        RECT 4.000 3.760 260.700 7.800 ;
        RECT 4.400 2.895 256.300 3.760 ;
      LAYER met4 ;
        RECT 9.495 12.415 20.640 254.145 ;
        RECT 23.040 12.415 97.440 254.145 ;
        RECT 99.840 12.415 174.240 254.145 ;
        RECT 176.640 12.415 250.865 254.145 ;
      LAYER met5 ;
        RECT 154.220 79.100 190.780 87.500 ;
  END
END clb_tile
END LIBRARY

