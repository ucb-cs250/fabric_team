VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block_north
  CLASS BLOCK ;
  FOREIGN baked_connection_block_north ;
  ORIGIN 0.000 0.000 ;
  SIZE 305.645 BY 316.365 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.910 312.365 8.190 316.365 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 312.365 23.830 316.365 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 312.365 39.930 316.365 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 312.365 56.030 316.365 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 312.365 72.130 316.365 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 312.365 88.230 316.365 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 312.365 104.330 316.365 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 312.365 120.430 316.365 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 312.365 136.530 316.365 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.350 312.365 152.630 316.365 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.450 312.365 168.730 316.365 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.550 312.365 184.830 316.365 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.650 312.365 200.930 316.365 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.750 312.365 217.030 316.365 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 312.365 233.130 316.365 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.950 312.365 249.230 316.365 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.050 312.365 265.330 316.365 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.150 312.365 281.430 316.365 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 118.360 305.645 118.960 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 144.200 305.645 144.800 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 170.720 305.645 171.320 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 197.240 305.645 197.840 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 223.760 305.645 224.360 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 249.600 305.645 250.200 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 276.120 305.645 276.720 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 302.640 305.645 303.240 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END double1[7]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.250 312.365 297.530 316.365 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 12.960 305.645 13.560 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 38.800 305.645 39.400 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 65.320 305.645 65.920 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 301.645 91.840 305.645 92.440 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 304.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 304.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 6.545 299.920 304.725 ;
      LAYER met1 ;
        RECT 4.685 6.515 299.920 312.080 ;
      LAYER met2 ;
        RECT 5.620 312.085 7.630 312.365 ;
        RECT 8.470 312.085 23.270 312.365 ;
        RECT 24.110 312.085 39.370 312.365 ;
        RECT 40.210 312.085 55.470 312.365 ;
        RECT 56.310 312.085 71.570 312.365 ;
        RECT 72.410 312.085 87.670 312.365 ;
        RECT 88.510 312.085 103.770 312.365 ;
        RECT 104.610 312.085 119.870 312.365 ;
        RECT 120.710 312.085 135.970 312.365 ;
        RECT 136.810 312.085 152.070 312.365 ;
        RECT 152.910 312.085 168.170 312.365 ;
        RECT 169.010 312.085 184.270 312.365 ;
        RECT 185.110 312.085 200.370 312.365 ;
        RECT 201.210 312.085 216.470 312.365 ;
        RECT 217.310 312.085 232.570 312.365 ;
        RECT 233.410 312.085 248.670 312.365 ;
        RECT 249.510 312.085 264.770 312.365 ;
        RECT 265.610 312.085 280.870 312.365 ;
        RECT 281.710 312.085 296.970 312.365 ;
        RECT 297.810 312.085 298.440 312.365 ;
        RECT 5.620 4.280 298.440 312.085 ;
        RECT 5.620 4.000 7.170 4.280 ;
        RECT 8.010 4.000 22.350 4.280 ;
        RECT 23.190 4.000 37.530 4.280 ;
        RECT 38.370 4.000 52.710 4.280 ;
        RECT 53.550 4.000 67.890 4.280 ;
        RECT 68.730 4.000 83.530 4.280 ;
        RECT 84.370 4.000 98.710 4.280 ;
        RECT 99.550 4.000 113.890 4.280 ;
        RECT 114.730 4.000 129.070 4.280 ;
        RECT 129.910 4.000 144.250 4.280 ;
        RECT 145.090 4.000 159.890 4.280 ;
        RECT 160.730 4.000 175.070 4.280 ;
        RECT 175.910 4.000 190.250 4.280 ;
        RECT 191.090 4.000 205.430 4.280 ;
        RECT 206.270 4.000 220.610 4.280 ;
        RECT 221.450 4.000 236.250 4.280 ;
        RECT 237.090 4.000 251.430 4.280 ;
        RECT 252.270 4.000 266.610 4.280 ;
        RECT 267.450 4.000 281.790 4.280 ;
        RECT 282.630 4.000 296.970 4.280 ;
        RECT 297.810 4.000 298.440 4.280 ;
      LAYER met3 ;
        RECT 4.000 304.320 301.645 304.805 ;
        RECT 4.400 303.640 301.645 304.320 ;
        RECT 4.400 302.920 301.245 303.640 ;
        RECT 4.000 302.240 301.245 302.920 ;
        RECT 4.000 279.840 301.645 302.240 ;
        RECT 4.400 278.440 301.645 279.840 ;
        RECT 4.000 277.120 301.645 278.440 ;
        RECT 4.000 275.720 301.245 277.120 ;
        RECT 4.000 255.360 301.645 275.720 ;
        RECT 4.400 253.960 301.645 255.360 ;
        RECT 4.000 250.600 301.645 253.960 ;
        RECT 4.000 249.200 301.245 250.600 ;
        RECT 4.000 230.880 301.645 249.200 ;
        RECT 4.400 229.480 301.645 230.880 ;
        RECT 4.000 224.760 301.645 229.480 ;
        RECT 4.000 223.360 301.245 224.760 ;
        RECT 4.000 207.080 301.645 223.360 ;
        RECT 4.400 205.680 301.645 207.080 ;
        RECT 4.000 198.240 301.645 205.680 ;
        RECT 4.000 196.840 301.245 198.240 ;
        RECT 4.000 182.600 301.645 196.840 ;
        RECT 4.400 181.200 301.645 182.600 ;
        RECT 4.000 171.720 301.645 181.200 ;
        RECT 4.000 170.320 301.245 171.720 ;
        RECT 4.000 158.120 301.645 170.320 ;
        RECT 4.400 156.720 301.645 158.120 ;
        RECT 4.000 145.200 301.645 156.720 ;
        RECT 4.000 143.800 301.245 145.200 ;
        RECT 4.000 133.640 301.645 143.800 ;
        RECT 4.400 132.240 301.645 133.640 ;
        RECT 4.000 119.360 301.645 132.240 ;
        RECT 4.000 117.960 301.245 119.360 ;
        RECT 4.000 109.840 301.645 117.960 ;
        RECT 4.400 108.440 301.645 109.840 ;
        RECT 4.000 92.840 301.645 108.440 ;
        RECT 4.000 91.440 301.245 92.840 ;
        RECT 4.000 85.360 301.645 91.440 ;
        RECT 4.400 83.960 301.645 85.360 ;
        RECT 4.000 66.320 301.645 83.960 ;
        RECT 4.000 64.920 301.245 66.320 ;
        RECT 4.000 60.880 301.645 64.920 ;
        RECT 4.400 59.480 301.645 60.880 ;
        RECT 4.000 39.800 301.645 59.480 ;
        RECT 4.000 38.400 301.245 39.800 ;
        RECT 4.000 36.400 301.645 38.400 ;
        RECT 4.400 35.000 301.645 36.400 ;
        RECT 4.000 13.960 301.645 35.000 ;
        RECT 4.000 12.600 301.245 13.960 ;
        RECT 4.400 12.560 301.245 12.600 ;
        RECT 4.400 11.200 301.645 12.560 ;
        RECT 4.000 10.715 301.645 11.200 ;
      LAYER met4 ;
        RECT 7.655 10.640 20.640 304.880 ;
        RECT 23.040 10.640 97.440 304.880 ;
        RECT 99.840 10.640 253.040 304.880 ;
  END
END baked_connection_block_north
END LIBRARY

