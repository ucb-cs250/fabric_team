VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block_north
  CLASS BLOCK ;
  FOREIGN baked_connection_block_north ;
  ORIGIN 0.000 0.000 ;
  SIZE 254.225 BY 264.945 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 236.000 254.225 236.600 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 260.945 7.270 264.945 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 260.945 21.070 264.945 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 260.945 35.330 264.945 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.310 260.945 49.590 264.945 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 260.945 63.390 264.945 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 260.945 77.650 264.945 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 260.945 91.910 264.945 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 260.945 106.170 264.945 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 260.945 119.970 264.945 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.950 260.945 134.230 264.945 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 260.945 148.490 264.945 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 260.945 162.290 264.945 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.270 260.945 176.550 264.945 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 260.945 190.810 264.945 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.790 260.945 205.070 264.945 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 260.945 218.870 264.945 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 260.945 233.130 264.945 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 84.360 254.225 84.960 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 103.400 254.225 104.000 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 122.440 254.225 123.040 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 141.480 254.225 142.080 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 159.840 254.225 160.440 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 178.880 254.225 179.480 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 197.920 254.225 198.520 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 216.960 254.225 217.560 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END double1[7]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 260.945 247.390 264.945 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 255.040 254.225 255.640 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 8.880 254.225 9.480 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 27.240 254.225 27.840 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 46.280 254.225 46.880 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 65.320 254.225 65.920 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 253.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 253.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 249.175 253.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 249.250 253.200 ;
      LAYER met2 ;
        RECT 7.550 260.665 20.510 260.945 ;
        RECT 21.350 260.665 34.770 260.945 ;
        RECT 35.610 260.665 49.030 260.945 ;
        RECT 49.870 260.665 62.830 260.945 ;
        RECT 63.670 260.665 77.090 260.945 ;
        RECT 77.930 260.665 91.350 260.945 ;
        RECT 92.190 260.665 105.610 260.945 ;
        RECT 106.450 260.665 119.410 260.945 ;
        RECT 120.250 260.665 133.670 260.945 ;
        RECT 134.510 260.665 147.930 260.945 ;
        RECT 148.770 260.665 161.730 260.945 ;
        RECT 162.570 260.665 175.990 260.945 ;
        RECT 176.830 260.665 190.250 260.945 ;
        RECT 191.090 260.665 204.510 260.945 ;
        RECT 205.350 260.665 218.310 260.945 ;
        RECT 219.150 260.665 232.570 260.945 ;
        RECT 233.410 260.665 246.830 260.945 ;
        RECT 247.670 260.665 249.230 260.945 ;
        RECT 7.000 4.280 249.230 260.665 ;
        RECT 7.550 4.000 20.510 4.280 ;
        RECT 21.350 4.000 34.770 4.280 ;
        RECT 35.610 4.000 49.030 4.280 ;
        RECT 49.870 4.000 62.830 4.280 ;
        RECT 63.670 4.000 77.090 4.280 ;
        RECT 77.930 4.000 91.350 4.280 ;
        RECT 92.190 4.000 105.610 4.280 ;
        RECT 106.450 4.000 119.410 4.280 ;
        RECT 120.250 4.000 133.670 4.280 ;
        RECT 134.510 4.000 147.930 4.280 ;
        RECT 148.770 4.000 161.730 4.280 ;
        RECT 162.570 4.000 175.990 4.280 ;
        RECT 176.830 4.000 190.250 4.280 ;
        RECT 191.090 4.000 204.510 4.280 ;
        RECT 205.350 4.000 218.310 4.280 ;
        RECT 219.150 4.000 232.570 4.280 ;
        RECT 233.410 4.000 246.830 4.280 ;
        RECT 247.670 4.000 249.230 4.280 ;
      LAYER met3 ;
        RECT 4.400 254.640 249.825 255.505 ;
        RECT 4.000 237.000 250.225 254.640 ;
        RECT 4.400 235.600 249.825 237.000 ;
        RECT 4.000 217.960 250.225 235.600 ;
        RECT 4.400 216.560 249.825 217.960 ;
        RECT 4.000 198.920 250.225 216.560 ;
        RECT 4.400 197.520 249.825 198.920 ;
        RECT 4.000 179.880 250.225 197.520 ;
        RECT 4.400 178.480 249.825 179.880 ;
        RECT 4.000 160.840 250.225 178.480 ;
        RECT 4.400 159.440 249.825 160.840 ;
        RECT 4.000 142.480 250.225 159.440 ;
        RECT 4.400 141.080 249.825 142.480 ;
        RECT 4.000 123.440 250.225 141.080 ;
        RECT 4.400 122.040 249.825 123.440 ;
        RECT 4.000 104.400 250.225 122.040 ;
        RECT 4.400 103.000 249.825 104.400 ;
        RECT 4.000 85.360 250.225 103.000 ;
        RECT 4.400 83.960 249.825 85.360 ;
        RECT 4.000 66.320 250.225 83.960 ;
        RECT 4.400 64.920 249.825 66.320 ;
        RECT 4.000 47.280 250.225 64.920 ;
        RECT 4.400 45.880 249.825 47.280 ;
        RECT 4.000 28.240 250.225 45.880 ;
        RECT 4.400 26.840 249.825 28.240 ;
        RECT 4.000 9.880 250.225 26.840 ;
        RECT 4.400 9.015 249.825 9.880 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 253.200 ;
  END
END baked_connection_block_north
END LIBRARY

