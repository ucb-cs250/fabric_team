VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 258.155 BY 268.875 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 264.875 240.030 268.875 ;
    END
  END COUT
  PIN cb_e_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 2.760 258.155 3.360 ;
    END
  END cb_e_clb1_input[0]
  PIN cb_e_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 8.200 258.155 8.800 ;
    END
  END cb_e_clb1_input[1]
  PIN cb_e_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 14.320 258.155 14.920 ;
    END
  END cb_e_clb1_input[2]
  PIN cb_e_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 19.760 258.155 20.360 ;
    END
  END cb_e_clb1_input[3]
  PIN cb_e_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 25.880 258.155 26.480 ;
    END
  END cb_e_clb1_input[4]
  PIN cb_e_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 31.320 258.155 31.920 ;
    END
  END cb_e_clb1_input[5]
  PIN cb_e_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 37.440 258.155 38.040 ;
    END
  END cb_e_clb1_input[6]
  PIN cb_e_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 43.560 258.155 44.160 ;
    END
  END cb_e_clb1_input[7]
  PIN cb_e_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 49.000 258.155 49.600 ;
    END
  END cb_e_clb1_input[8]
  PIN cb_e_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 55.120 258.155 55.720 ;
    END
  END cb_e_clb1_input[9]
  PIN cb_e_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 60.560 258.155 61.160 ;
    END
  END cb_e_clb1_output[0]
  PIN cb_e_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 66.680 258.155 67.280 ;
    END
  END cb_e_clb1_output[1]
  PIN cb_e_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 72.800 258.155 73.400 ;
    END
  END cb_e_clb1_output[2]
  PIN cb_e_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 78.240 258.155 78.840 ;
    END
  END cb_e_clb1_output[3]
  PIN cb_e_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END cb_e_single1_in[0]
  PIN cb_e_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END cb_e_single1_in[10]
  PIN cb_e_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END cb_e_single1_in[11]
  PIN cb_e_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END cb_e_single1_in[12]
  PIN cb_e_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END cb_e_single1_in[13]
  PIN cb_e_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END cb_e_single1_in[14]
  PIN cb_e_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END cb_e_single1_in[15]
  PIN cb_e_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END cb_e_single1_in[1]
  PIN cb_e_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END cb_e_single1_in[2]
  PIN cb_e_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END cb_e_single1_in[3]
  PIN cb_e_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END cb_e_single1_in[4]
  PIN cb_e_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END cb_e_single1_in[5]
  PIN cb_e_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END cb_e_single1_in[6]
  PIN cb_e_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END cb_e_single1_in[7]
  PIN cb_e_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END cb_e_single1_in[8]
  PIN cb_e_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END cb_e_single1_in[9]
  PIN cb_e_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END cb_e_single1_out[0]
  PIN cb_e_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END cb_e_single1_out[10]
  PIN cb_e_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END cb_e_single1_out[11]
  PIN cb_e_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END cb_e_single1_out[12]
  PIN cb_e_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END cb_e_single1_out[13]
  PIN cb_e_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END cb_e_single1_out[14]
  PIN cb_e_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END cb_e_single1_out[15]
  PIN cb_e_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END cb_e_single1_out[1]
  PIN cb_e_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END cb_e_single1_out[2]
  PIN cb_e_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END cb_e_single1_out[3]
  PIN cb_e_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END cb_e_single1_out[4]
  PIN cb_e_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END cb_e_single1_out[5]
  PIN cb_e_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END cb_e_single1_out[6]
  PIN cb_e_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END cb_e_single1_out[7]
  PIN cb_e_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END cb_e_single1_out[8]
  PIN cb_e_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END cb_e_single1_out[9]
  PIN cb_n_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 264.875 2.670 268.875 ;
    END
  END cb_n_clb1_input[0]
  PIN cb_n_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 264.875 7.730 268.875 ;
    END
  END cb_n_clb1_input[1]
  PIN cb_n_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 264.875 12.790 268.875 ;
    END
  END cb_n_clb1_input[2]
  PIN cb_n_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 264.875 17.850 268.875 ;
    END
  END cb_n_clb1_input[3]
  PIN cb_n_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 264.875 22.910 268.875 ;
    END
  END cb_n_clb1_input[4]
  PIN cb_n_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 264.875 28.430 268.875 ;
    END
  END cb_n_clb1_input[5]
  PIN cb_n_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 264.875 33.490 268.875 ;
    END
  END cb_n_clb1_input[6]
  PIN cb_n_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 264.875 38.550 268.875 ;
    END
  END cb_n_clb1_input[7]
  PIN cb_n_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 264.875 43.610 268.875 ;
    END
  END cb_n_clb1_input[8]
  PIN cb_n_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 264.875 48.670 268.875 ;
    END
  END cb_n_clb1_input[9]
  PIN cb_n_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 264.875 54.190 268.875 ;
    END
  END cb_n_clb1_output[0]
  PIN cb_n_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 264.875 59.250 268.875 ;
    END
  END cb_n_clb1_output[1]
  PIN cb_n_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 264.875 64.310 268.875 ;
    END
  END cb_n_clb1_output[2]
  PIN cb_n_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 264.875 69.370 268.875 ;
    END
  END cb_n_clb1_output[3]
  PIN cb_n_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END cb_n_single1_in[0]
  PIN cb_n_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END cb_n_single1_in[10]
  PIN cb_n_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END cb_n_single1_in[11]
  PIN cb_n_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END cb_n_single1_in[12]
  PIN cb_n_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END cb_n_single1_in[13]
  PIN cb_n_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END cb_n_single1_in[14]
  PIN cb_n_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END cb_n_single1_in[15]
  PIN cb_n_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END cb_n_single1_in[1]
  PIN cb_n_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END cb_n_single1_in[2]
  PIN cb_n_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END cb_n_single1_in[3]
  PIN cb_n_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END cb_n_single1_in[4]
  PIN cb_n_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END cb_n_single1_in[5]
  PIN cb_n_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END cb_n_single1_in[6]
  PIN cb_n_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END cb_n_single1_in[7]
  PIN cb_n_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END cb_n_single1_in[8]
  PIN cb_n_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END cb_n_single1_in[9]
  PIN cb_n_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END cb_n_single1_out[0]
  PIN cb_n_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END cb_n_single1_out[10]
  PIN cb_n_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END cb_n_single1_out[11]
  PIN cb_n_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END cb_n_single1_out[12]
  PIN cb_n_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END cb_n_single1_out[13]
  PIN cb_n_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END cb_n_single1_out[14]
  PIN cb_n_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END cb_n_single1_out[15]
  PIN cb_n_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END cb_n_single1_out[1]
  PIN cb_n_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END cb_n_single1_out[2]
  PIN cb_n_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END cb_n_single1_out[3]
  PIN cb_n_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END cb_n_single1_out[4]
  PIN cb_n_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END cb_n_single1_out[5]
  PIN cb_n_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END cb_n_single1_out[6]
  PIN cb_n_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END cb_n_single1_out[7]
  PIN cb_n_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END cb_n_single1_out[8]
  PIN cb_n_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END cb_n_single1_out[9]
  PIN cfg_bit_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END cfg_bit_in
  PIN cfg_bit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 264.875 250.150 268.875 ;
    END
  END cfg_bit_out
  PIN cfg_in_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END cfg_in_start
  PIN cfg_out_start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 264.875 245.090 268.875 ;
    END
  END cfg_out_start
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END clb_south_out[3]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END clb_west_out[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END clk
  PIN crst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 264.875 255.210 268.875 ;
    END
  END crst
  PIN sb_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 84.360 258.155 84.960 ;
    END
  END sb_east_in[0]
  PIN sb_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 142.840 258.155 143.440 ;
    END
  END sb_east_in[10]
  PIN sb_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 148.280 258.155 148.880 ;
    END
  END sb_east_in[11]
  PIN sb_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 154.400 258.155 155.000 ;
    END
  END sb_east_in[12]
  PIN sb_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 159.840 258.155 160.440 ;
    END
  END sb_east_in[13]
  PIN sb_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 165.960 258.155 166.560 ;
    END
  END sb_east_in[14]
  PIN sb_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 172.080 258.155 172.680 ;
    END
  END sb_east_in[15]
  PIN sb_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 89.800 258.155 90.400 ;
    END
  END sb_east_in[1]
  PIN sb_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 95.920 258.155 96.520 ;
    END
  END sb_east_in[2]
  PIN sb_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 101.360 258.155 101.960 ;
    END
  END sb_east_in[3]
  PIN sb_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 107.480 258.155 108.080 ;
    END
  END sb_east_in[4]
  PIN sb_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 113.600 258.155 114.200 ;
    END
  END sb_east_in[5]
  PIN sb_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 119.040 258.155 119.640 ;
    END
  END sb_east_in[6]
  PIN sb_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 125.160 258.155 125.760 ;
    END
  END sb_east_in[7]
  PIN sb_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 130.600 258.155 131.200 ;
    END
  END sb_east_in[8]
  PIN sb_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 136.720 258.155 137.320 ;
    END
  END sb_east_in[9]
  PIN sb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 177.520 258.155 178.120 ;
    END
  END sb_east_out[0]
  PIN sb_east_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 236.000 258.155 236.600 ;
    END
  END sb_east_out[10]
  PIN sb_east_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 242.120 258.155 242.720 ;
    END
  END sb_east_out[11]
  PIN sb_east_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 247.560 258.155 248.160 ;
    END
  END sb_east_out[12]
  PIN sb_east_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 253.680 258.155 254.280 ;
    END
  END sb_east_out[13]
  PIN sb_east_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 259.120 258.155 259.720 ;
    END
  END sb_east_out[14]
  PIN sb_east_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 265.240 258.155 265.840 ;
    END
  END sb_east_out[15]
  PIN sb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 183.640 258.155 184.240 ;
    END
  END sb_east_out[1]
  PIN sb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 189.080 258.155 189.680 ;
    END
  END sb_east_out[2]
  PIN sb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 195.200 258.155 195.800 ;
    END
  END sb_east_out[3]
  PIN sb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 200.640 258.155 201.240 ;
    END
  END sb_east_out[4]
  PIN sb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 206.760 258.155 207.360 ;
    END
  END sb_east_out[5]
  PIN sb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 212.880 258.155 213.480 ;
    END
  END sb_east_out[6]
  PIN sb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 218.320 258.155 218.920 ;
    END
  END sb_east_out[7]
  PIN sb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 224.440 258.155 225.040 ;
    END
  END sb_east_out[8]
  PIN sb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.155 229.880 258.155 230.480 ;
    END
  END sb_east_out[9]
  PIN sb_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 264.875 74.890 268.875 ;
    END
  END sb_north_in[0]
  PIN sb_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 264.875 126.410 268.875 ;
    END
  END sb_north_in[10]
  PIN sb_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 264.875 131.470 268.875 ;
    END
  END sb_north_in[11]
  PIN sb_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 264.875 136.530 268.875 ;
    END
  END sb_north_in[12]
  PIN sb_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 264.875 141.590 268.875 ;
    END
  END sb_north_in[13]
  PIN sb_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 264.875 147.110 268.875 ;
    END
  END sb_north_in[14]
  PIN sb_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 264.875 152.170 268.875 ;
    END
  END sb_north_in[15]
  PIN sb_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 264.875 79.950 268.875 ;
    END
  END sb_north_in[1]
  PIN sb_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 264.875 85.010 268.875 ;
    END
  END sb_north_in[2]
  PIN sb_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 264.875 90.070 268.875 ;
    END
  END sb_north_in[3]
  PIN sb_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 264.875 95.130 268.875 ;
    END
  END sb_north_in[4]
  PIN sb_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 264.875 100.650 268.875 ;
    END
  END sb_north_in[5]
  PIN sb_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 264.875 105.710 268.875 ;
    END
  END sb_north_in[6]
  PIN sb_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 264.875 110.770 268.875 ;
    END
  END sb_north_in[7]
  PIN sb_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 264.875 115.830 268.875 ;
    END
  END sb_north_in[8]
  PIN sb_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 264.875 121.350 268.875 ;
    END
  END sb_north_in[9]
  PIN sb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 264.875 157.230 268.875 ;
    END
  END sb_north_out[0]
  PIN sb_north_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 264.875 208.750 268.875 ;
    END
  END sb_north_out[10]
  PIN sb_north_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 264.875 214.270 268.875 ;
    END
  END sb_north_out[11]
  PIN sb_north_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 264.875 219.330 268.875 ;
    END
  END sb_north_out[12]
  PIN sb_north_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 264.875 224.390 268.875 ;
    END
  END sb_north_out[13]
  PIN sb_north_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 264.875 229.450 268.875 ;
    END
  END sb_north_out[14]
  PIN sb_north_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 264.875 234.510 268.875 ;
    END
  END sb_north_out[15]
  PIN sb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 264.875 162.290 268.875 ;
    END
  END sb_north_out[1]
  PIN sb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 264.875 167.810 268.875 ;
    END
  END sb_north_out[2]
  PIN sb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 264.875 172.870 268.875 ;
    END
  END sb_north_out[3]
  PIN sb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 264.875 177.930 268.875 ;
    END
  END sb_north_out[4]
  PIN sb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 264.875 182.990 268.875 ;
    END
  END sb_north_out[5]
  PIN sb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 264.875 188.050 268.875 ;
    END
  END sb_north_out[6]
  PIN sb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 264.875 193.570 268.875 ;
    END
  END sb_north_out[7]
  PIN sb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 264.875 198.630 268.875 ;
    END
  END sb_north_out[8]
  PIN sb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 264.875 203.690 268.875 ;
    END
  END sb_north_out[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 255.920 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 255.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 255.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 7.565 253.315 255.765 ;
      LAYER met1 ;
        RECT 2.370 6.160 255.230 260.060 ;
      LAYER met2 ;
        RECT 2.950 264.595 7.170 265.725 ;
        RECT 8.010 264.595 12.230 265.725 ;
        RECT 13.070 264.595 17.290 265.725 ;
        RECT 18.130 264.595 22.350 265.725 ;
        RECT 23.190 264.595 27.870 265.725 ;
        RECT 28.710 264.595 32.930 265.725 ;
        RECT 33.770 264.595 37.990 265.725 ;
        RECT 38.830 264.595 43.050 265.725 ;
        RECT 43.890 264.595 48.110 265.725 ;
        RECT 48.950 264.595 53.630 265.725 ;
        RECT 54.470 264.595 58.690 265.725 ;
        RECT 59.530 264.595 63.750 265.725 ;
        RECT 64.590 264.595 68.810 265.725 ;
        RECT 69.650 264.595 74.330 265.725 ;
        RECT 75.170 264.595 79.390 265.725 ;
        RECT 80.230 264.595 84.450 265.725 ;
        RECT 85.290 264.595 89.510 265.725 ;
        RECT 90.350 264.595 94.570 265.725 ;
        RECT 95.410 264.595 100.090 265.725 ;
        RECT 100.930 264.595 105.150 265.725 ;
        RECT 105.990 264.595 110.210 265.725 ;
        RECT 111.050 264.595 115.270 265.725 ;
        RECT 116.110 264.595 120.790 265.725 ;
        RECT 121.630 264.595 125.850 265.725 ;
        RECT 126.690 264.595 130.910 265.725 ;
        RECT 131.750 264.595 135.970 265.725 ;
        RECT 136.810 264.595 141.030 265.725 ;
        RECT 141.870 264.595 146.550 265.725 ;
        RECT 147.390 264.595 151.610 265.725 ;
        RECT 152.450 264.595 156.670 265.725 ;
        RECT 157.510 264.595 161.730 265.725 ;
        RECT 162.570 264.595 167.250 265.725 ;
        RECT 168.090 264.595 172.310 265.725 ;
        RECT 173.150 264.595 177.370 265.725 ;
        RECT 178.210 264.595 182.430 265.725 ;
        RECT 183.270 264.595 187.490 265.725 ;
        RECT 188.330 264.595 193.010 265.725 ;
        RECT 193.850 264.595 198.070 265.725 ;
        RECT 198.910 264.595 203.130 265.725 ;
        RECT 203.970 264.595 208.190 265.725 ;
        RECT 209.030 264.595 213.710 265.725 ;
        RECT 214.550 264.595 218.770 265.725 ;
        RECT 219.610 264.595 223.830 265.725 ;
        RECT 224.670 264.595 228.890 265.725 ;
        RECT 229.730 264.595 233.950 265.725 ;
        RECT 234.790 264.595 239.470 265.725 ;
        RECT 240.310 264.595 244.530 265.725 ;
        RECT 245.370 264.595 249.590 265.725 ;
        RECT 250.430 264.595 254.650 265.725 ;
        RECT 2.400 4.280 255.200 264.595 ;
        RECT 2.950 2.875 7.170 4.280 ;
        RECT 8.010 2.875 12.230 4.280 ;
        RECT 13.070 2.875 17.750 4.280 ;
        RECT 18.590 2.875 22.810 4.280 ;
        RECT 23.650 2.875 28.330 4.280 ;
        RECT 29.170 2.875 33.390 4.280 ;
        RECT 34.230 2.875 38.910 4.280 ;
        RECT 39.750 2.875 43.970 4.280 ;
        RECT 44.810 2.875 49.490 4.280 ;
        RECT 50.330 2.875 54.550 4.280 ;
        RECT 55.390 2.875 59.610 4.280 ;
        RECT 60.450 2.875 65.130 4.280 ;
        RECT 65.970 2.875 70.190 4.280 ;
        RECT 71.030 2.875 75.710 4.280 ;
        RECT 76.550 2.875 80.770 4.280 ;
        RECT 81.610 2.875 86.290 4.280 ;
        RECT 87.130 2.875 91.350 4.280 ;
        RECT 92.190 2.875 96.870 4.280 ;
        RECT 97.710 2.875 101.930 4.280 ;
        RECT 102.770 2.875 106.990 4.280 ;
        RECT 107.830 2.875 112.510 4.280 ;
        RECT 113.350 2.875 117.570 4.280 ;
        RECT 118.410 2.875 123.090 4.280 ;
        RECT 123.930 2.875 128.150 4.280 ;
        RECT 128.990 2.875 133.670 4.280 ;
        RECT 134.510 2.875 138.730 4.280 ;
        RECT 139.570 2.875 144.250 4.280 ;
        RECT 145.090 2.875 149.310 4.280 ;
        RECT 150.150 2.875 154.830 4.280 ;
        RECT 155.670 2.875 159.890 4.280 ;
        RECT 160.730 2.875 164.950 4.280 ;
        RECT 165.790 2.875 170.470 4.280 ;
        RECT 171.310 2.875 175.530 4.280 ;
        RECT 176.370 2.875 181.050 4.280 ;
        RECT 181.890 2.875 186.110 4.280 ;
        RECT 186.950 2.875 191.630 4.280 ;
        RECT 192.470 2.875 196.690 4.280 ;
        RECT 197.530 2.875 202.210 4.280 ;
        RECT 203.050 2.875 207.270 4.280 ;
        RECT 208.110 2.875 212.330 4.280 ;
        RECT 213.170 2.875 217.850 4.280 ;
        RECT 218.690 2.875 222.910 4.280 ;
        RECT 223.750 2.875 228.430 4.280 ;
        RECT 229.270 2.875 233.490 4.280 ;
        RECT 234.330 2.875 239.010 4.280 ;
        RECT 239.850 2.875 244.070 4.280 ;
        RECT 244.910 2.875 249.590 4.280 ;
        RECT 250.430 2.875 254.650 4.280 ;
      LAYER met3 ;
        RECT 4.400 264.840 253.755 265.705 ;
        RECT 3.990 260.800 254.155 264.840 ;
        RECT 4.400 260.120 254.155 260.800 ;
        RECT 4.400 259.400 253.755 260.120 ;
        RECT 3.990 258.720 253.755 259.400 ;
        RECT 3.990 254.680 254.155 258.720 ;
        RECT 4.400 253.280 253.755 254.680 ;
        RECT 3.990 249.240 254.155 253.280 ;
        RECT 4.400 248.560 254.155 249.240 ;
        RECT 4.400 247.840 253.755 248.560 ;
        RECT 3.990 247.160 253.755 247.840 ;
        RECT 3.990 243.120 254.155 247.160 ;
        RECT 4.400 241.720 253.755 243.120 ;
        RECT 3.990 237.680 254.155 241.720 ;
        RECT 4.400 237.000 254.155 237.680 ;
        RECT 4.400 236.280 253.755 237.000 ;
        RECT 3.990 235.600 253.755 236.280 ;
        RECT 3.990 232.240 254.155 235.600 ;
        RECT 4.400 230.880 254.155 232.240 ;
        RECT 4.400 230.840 253.755 230.880 ;
        RECT 3.990 229.480 253.755 230.840 ;
        RECT 3.990 226.120 254.155 229.480 ;
        RECT 4.400 225.440 254.155 226.120 ;
        RECT 4.400 224.720 253.755 225.440 ;
        RECT 3.990 224.040 253.755 224.720 ;
        RECT 3.990 220.680 254.155 224.040 ;
        RECT 4.400 219.320 254.155 220.680 ;
        RECT 4.400 219.280 253.755 219.320 ;
        RECT 3.990 217.920 253.755 219.280 ;
        RECT 3.990 214.560 254.155 217.920 ;
        RECT 4.400 213.880 254.155 214.560 ;
        RECT 4.400 213.160 253.755 213.880 ;
        RECT 3.990 212.480 253.755 213.160 ;
        RECT 3.990 209.120 254.155 212.480 ;
        RECT 4.400 207.760 254.155 209.120 ;
        RECT 4.400 207.720 253.755 207.760 ;
        RECT 3.990 206.360 253.755 207.720 ;
        RECT 3.990 203.680 254.155 206.360 ;
        RECT 4.400 202.280 254.155 203.680 ;
        RECT 3.990 201.640 254.155 202.280 ;
        RECT 3.990 200.240 253.755 201.640 ;
        RECT 3.990 197.560 254.155 200.240 ;
        RECT 4.400 196.200 254.155 197.560 ;
        RECT 4.400 196.160 253.755 196.200 ;
        RECT 3.990 194.800 253.755 196.160 ;
        RECT 3.990 192.120 254.155 194.800 ;
        RECT 4.400 190.720 254.155 192.120 ;
        RECT 3.990 190.080 254.155 190.720 ;
        RECT 3.990 188.680 253.755 190.080 ;
        RECT 3.990 186.000 254.155 188.680 ;
        RECT 4.400 184.640 254.155 186.000 ;
        RECT 4.400 184.600 253.755 184.640 ;
        RECT 3.990 183.240 253.755 184.600 ;
        RECT 3.990 180.560 254.155 183.240 ;
        RECT 4.400 179.160 254.155 180.560 ;
        RECT 3.990 178.520 254.155 179.160 ;
        RECT 3.990 177.120 253.755 178.520 ;
        RECT 3.990 175.120 254.155 177.120 ;
        RECT 4.400 173.720 254.155 175.120 ;
        RECT 3.990 173.080 254.155 173.720 ;
        RECT 3.990 171.680 253.755 173.080 ;
        RECT 3.990 169.000 254.155 171.680 ;
        RECT 4.400 167.600 254.155 169.000 ;
        RECT 3.990 166.960 254.155 167.600 ;
        RECT 3.990 165.560 253.755 166.960 ;
        RECT 3.990 163.560 254.155 165.560 ;
        RECT 4.400 162.160 254.155 163.560 ;
        RECT 3.990 160.840 254.155 162.160 ;
        RECT 3.990 159.440 253.755 160.840 ;
        RECT 3.990 157.440 254.155 159.440 ;
        RECT 4.400 156.040 254.155 157.440 ;
        RECT 3.990 155.400 254.155 156.040 ;
        RECT 3.990 154.000 253.755 155.400 ;
        RECT 3.990 152.000 254.155 154.000 ;
        RECT 4.400 150.600 254.155 152.000 ;
        RECT 3.990 149.280 254.155 150.600 ;
        RECT 3.990 147.880 253.755 149.280 ;
        RECT 3.990 146.560 254.155 147.880 ;
        RECT 4.400 145.160 254.155 146.560 ;
        RECT 3.990 143.840 254.155 145.160 ;
        RECT 3.990 142.440 253.755 143.840 ;
        RECT 3.990 140.440 254.155 142.440 ;
        RECT 4.400 139.040 254.155 140.440 ;
        RECT 3.990 137.720 254.155 139.040 ;
        RECT 3.990 136.320 253.755 137.720 ;
        RECT 3.990 135.000 254.155 136.320 ;
        RECT 4.400 133.600 254.155 135.000 ;
        RECT 3.990 131.600 254.155 133.600 ;
        RECT 3.990 130.200 253.755 131.600 ;
        RECT 3.990 128.880 254.155 130.200 ;
        RECT 4.400 127.480 254.155 128.880 ;
        RECT 3.990 126.160 254.155 127.480 ;
        RECT 3.990 124.760 253.755 126.160 ;
        RECT 3.990 123.440 254.155 124.760 ;
        RECT 4.400 122.040 254.155 123.440 ;
        RECT 3.990 120.040 254.155 122.040 ;
        RECT 3.990 118.640 253.755 120.040 ;
        RECT 3.990 118.000 254.155 118.640 ;
        RECT 4.400 116.600 254.155 118.000 ;
        RECT 3.990 114.600 254.155 116.600 ;
        RECT 3.990 113.200 253.755 114.600 ;
        RECT 3.990 111.880 254.155 113.200 ;
        RECT 4.400 110.480 254.155 111.880 ;
        RECT 3.990 108.480 254.155 110.480 ;
        RECT 3.990 107.080 253.755 108.480 ;
        RECT 3.990 106.440 254.155 107.080 ;
        RECT 4.400 105.040 254.155 106.440 ;
        RECT 3.990 102.360 254.155 105.040 ;
        RECT 3.990 100.960 253.755 102.360 ;
        RECT 3.990 100.320 254.155 100.960 ;
        RECT 4.400 98.920 254.155 100.320 ;
        RECT 3.990 96.920 254.155 98.920 ;
        RECT 3.990 95.520 253.755 96.920 ;
        RECT 3.990 94.880 254.155 95.520 ;
        RECT 4.400 93.480 254.155 94.880 ;
        RECT 3.990 90.800 254.155 93.480 ;
        RECT 3.990 89.440 253.755 90.800 ;
        RECT 4.400 89.400 253.755 89.440 ;
        RECT 4.400 88.040 254.155 89.400 ;
        RECT 3.990 85.360 254.155 88.040 ;
        RECT 3.990 83.960 253.755 85.360 ;
        RECT 3.990 83.320 254.155 83.960 ;
        RECT 4.400 81.920 254.155 83.320 ;
        RECT 3.990 79.240 254.155 81.920 ;
        RECT 3.990 77.880 253.755 79.240 ;
        RECT 4.400 77.840 253.755 77.880 ;
        RECT 4.400 76.480 254.155 77.840 ;
        RECT 3.990 73.800 254.155 76.480 ;
        RECT 3.990 72.400 253.755 73.800 ;
        RECT 3.990 71.760 254.155 72.400 ;
        RECT 4.400 70.360 254.155 71.760 ;
        RECT 3.990 67.680 254.155 70.360 ;
        RECT 3.990 66.320 253.755 67.680 ;
        RECT 4.400 66.280 253.755 66.320 ;
        RECT 4.400 64.920 254.155 66.280 ;
        RECT 3.990 61.560 254.155 64.920 ;
        RECT 3.990 60.880 253.755 61.560 ;
        RECT 4.400 60.160 253.755 60.880 ;
        RECT 4.400 59.480 254.155 60.160 ;
        RECT 3.990 56.120 254.155 59.480 ;
        RECT 3.990 54.760 253.755 56.120 ;
        RECT 4.400 54.720 253.755 54.760 ;
        RECT 4.400 53.360 254.155 54.720 ;
        RECT 3.990 50.000 254.155 53.360 ;
        RECT 3.990 49.320 253.755 50.000 ;
        RECT 4.400 48.600 253.755 49.320 ;
        RECT 4.400 47.920 254.155 48.600 ;
        RECT 3.990 44.560 254.155 47.920 ;
        RECT 3.990 43.200 253.755 44.560 ;
        RECT 4.400 43.160 253.755 43.200 ;
        RECT 4.400 41.800 254.155 43.160 ;
        RECT 3.990 38.440 254.155 41.800 ;
        RECT 3.990 37.760 253.755 38.440 ;
        RECT 4.400 37.040 253.755 37.760 ;
        RECT 4.400 36.360 254.155 37.040 ;
        RECT 3.990 32.320 254.155 36.360 ;
        RECT 4.400 30.920 253.755 32.320 ;
        RECT 3.990 26.880 254.155 30.920 ;
        RECT 3.990 26.200 253.755 26.880 ;
        RECT 4.400 25.480 253.755 26.200 ;
        RECT 4.400 24.800 254.155 25.480 ;
        RECT 3.990 20.760 254.155 24.800 ;
        RECT 4.400 19.360 253.755 20.760 ;
        RECT 3.990 15.320 254.155 19.360 ;
        RECT 3.990 14.640 253.755 15.320 ;
        RECT 4.400 13.920 253.755 14.640 ;
        RECT 4.400 13.240 254.155 13.920 ;
        RECT 3.990 9.200 254.155 13.240 ;
        RECT 4.400 7.800 253.755 9.200 ;
        RECT 3.990 3.760 254.155 7.800 ;
        RECT 4.400 2.895 253.755 3.760 ;
      LAYER met4 ;
        RECT 9.495 256.320 243.505 265.705 ;
        RECT 9.495 11.055 20.640 256.320 ;
        RECT 23.040 11.055 97.440 256.320 ;
        RECT 99.840 11.055 174.240 256.320 ;
        RECT 176.640 11.055 243.505 256.320 ;
      LAYER met5 ;
        RECT 190.100 38.300 210.100 39.900 ;
  END
END clb_tile
END LIBRARY

