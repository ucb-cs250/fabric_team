module wishbone_configuratorinator_10 (cen,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    VPWR,
    VGND,
    set_out,
    shift_out,
    wbs_addr_i,
    wbs_data_i,
    wbs_data_o,
    wbs_sel_i);
 output cen;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input VPWR;
 input VGND;
 output [3:0] set_out;
 output [3:0] shift_out;
 input [31:0] wbs_addr_i;
 input [31:0] wbs_data_i;
 output [31:0] wbs_data_o;
 input [3:0] wbs_sel_i;

 sky130_fd_sc_hd__nor2_4 _0671_ (.A(wb_rst_i),
    .B(wbs_ack_o),
    .Y(_0108_));
 sky130_fd_sc_hd__buf_2 _0672_ (.A(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_2 _0673_ (.A(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(wbs_addr_i[4]),
    .Y(_0111_));
 sky130_fd_sc_hd__or4_4 _0675_ (.A(wbs_addr_i[5]),
    .B(_0111_),
    .C(wbs_addr_i[7]),
    .D(wbs_addr_i[6]),
    .X(_0112_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(wbs_cyc_i),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(wbs_stb_i),
    .Y(_0114_));
 sky130_fd_sc_hd__or4_4 _0678_ (.A(\configy.read_transaction_in_progress ),
    .B(wbs_ack_o),
    .C(_0113_),
    .D(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__or4_4 _0679_ (.A(wbs_addr_i[16]),
    .B(wbs_addr_i[19]),
    .C(wbs_addr_i[21]),
    .D(wbs_addr_i[22]),
    .X(_0116_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(wbs_addr_i[28]),
    .Y(_0117_));
 sky130_fd_sc_hd__or4_4 _0681_ (.A(wbs_addr_i[25]),
    .B(wbs_addr_i[26]),
    .C(_0117_),
    .D(wbs_addr_i[31]),
    .X(_0118_));
 sky130_fd_sc_hd__nor4_4 _0682_ (.A(_0112_),
    .B(_0115_),
    .C(_0116_),
    .D(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__buf_2 _0683_ (.A(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_2 _0684_ (.A(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or4_4 _0685_ (.A(wbs_addr_i[13]),
    .B(wbs_addr_i[12]),
    .C(wbs_addr_i[15]),
    .D(wbs_addr_i[14]),
    .X(_0122_));
 sky130_fd_sc_hd__or4_4 _0686_ (.A(wbs_addr_i[9]),
    .B(wbs_addr_i[8]),
    .C(wbs_addr_i[11]),
    .D(wbs_addr_i[10]),
    .X(_0123_));
 sky130_fd_sc_hd__or2_4 _0687_ (.A(_0122_),
    .B(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__or4_4 _0688_ (.A(wbs_addr_i[17]),
    .B(wbs_addr_i[18]),
    .C(wbs_addr_i[20]),
    .D(wbs_addr_i[23]),
    .X(_0125_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(wbs_addr_i[29]),
    .Y(_0126_));
 sky130_fd_sc_hd__or4_4 _0690_ (.A(wbs_addr_i[24]),
    .B(wbs_addr_i[27]),
    .C(_0126_),
    .D(wbs_addr_i[30]),
    .X(_0127_));
 sky130_fd_sc_hd__nor3_4 _0691_ (.A(_0124_),
    .B(_0125_),
    .C(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__buf_2 _0692_ (.A(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__buf_2 _0693_ (.A(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__a21o_4 _0694_ (.A1(_0121_),
    .A2(_0130_),
    .B1(wbs_data_o[30]),
    .X(_0131_));
 sky130_fd_sc_hd__nor3_4 _0695_ (.A(wbs_addr_i[1]),
    .B(wbs_addr_i[0]),
    .C(wbs_addr_i[2]),
    .Y(_0132_));
 sky130_fd_sc_hd__and2_4 _0696_ (.A(wbs_addr_i[3]),
    .B(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_2 _0697_ (.A(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_4 _0698_ (.A(\configy.counter_d[6] ),
    .B(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(wbs_addr_i[1]),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(wbs_addr_i[0]),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(wbs_addr_i[3]),
    .Y(_0138_));
 sky130_fd_sc_hd__and4_4 _0702_ (.A(_0136_),
    .B(_0137_),
    .C(_0138_),
    .D(wbs_addr_i[2]),
    .X(_0139_));
 sky130_fd_sc_hd__buf_2 _0703_ (.A(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__and2_4 _0704_ (.A(\configy.bits_d[6] ),
    .B(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__or4_4 _0705_ (.A(_0112_),
    .B(_0115_),
    .C(_0116_),
    .D(_0118_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_2 _0706_ (.A(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__or3_4 _0707_ (.A(_0124_),
    .B(_0125_),
    .C(_0127_),
    .X(_0144_));
 sky130_fd_sc_hd__buf_2 _0708_ (.A(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__buf_2 _0709_ (.A(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__or4_4 _0710_ (.A(_0135_),
    .B(_0141_),
    .C(_0143_),
    .D(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__and3_4 _0711_ (.A(_0110_),
    .B(_0131_),
    .C(_0147_),
    .X(_0106_));
 sky130_fd_sc_hd__a21o_4 _0712_ (.A1(_0121_),
    .A2(_0130_),
    .B1(wbs_data_o[29]),
    .X(_0148_));
 sky130_fd_sc_hd__buf_2 _0713_ (.A(\configy.counter_d[5] ),
    .X(_0149_));
 sky130_fd_sc_hd__buf_2 _0714_ (.A(_0134_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_4 _0715_ (.A(_0149_),
    .B(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__buf_2 _0716_ (.A(_0140_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_4 _0717_ (.A(\configy.bits_d[5] ),
    .B(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__or4_4 _0718_ (.A(_0143_),
    .B(_0146_),
    .C(_0151_),
    .D(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__and3_4 _0719_ (.A(_0110_),
    .B(_0148_),
    .C(_0154_),
    .X(_0105_));
 sky130_fd_sc_hd__a21o_4 _0720_ (.A1(_0121_),
    .A2(_0130_),
    .B1(wbs_data_o[28]),
    .X(_0155_));
 sky130_fd_sc_hd__and2_4 _0721_ (.A(\configy.counter_d[4] ),
    .B(_0150_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_4 _0722_ (.A(\configy.bits_d[4] ),
    .B(_0152_),
    .X(_0157_));
 sky130_fd_sc_hd__or4_4 _0723_ (.A(_0143_),
    .B(_0146_),
    .C(_0156_),
    .D(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__and3_4 _0724_ (.A(_0110_),
    .B(_0155_),
    .C(_0158_),
    .X(_0104_));
 sky130_fd_sc_hd__a21o_4 _0725_ (.A1(_0121_),
    .A2(_0130_),
    .B1(wbs_data_o[27]),
    .X(_0159_));
 sky130_fd_sc_hd__and2_4 _0726_ (.A(\configy.counter_d[3] ),
    .B(_0150_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_4 _0727_ (.A(\configy.bits_d[3] ),
    .B(_0152_),
    .X(_0161_));
 sky130_fd_sc_hd__or4_4 _0728_ (.A(_0143_),
    .B(_0146_),
    .C(_0160_),
    .D(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__and3_4 _0729_ (.A(_0110_),
    .B(_0159_),
    .C(_0162_),
    .X(_0103_));
 sky130_fd_sc_hd__buf_2 _0730_ (.A(_0109_),
    .X(_0163_));
 sky130_fd_sc_hd__buf_2 _0731_ (.A(_0119_),
    .X(_0164_));
 sky130_fd_sc_hd__buf_2 _0732_ (.A(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _0733_ (.A(_0128_),
    .X(_0166_));
 sky130_fd_sc_hd__buf_2 _0734_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__a21o_4 _0735_ (.A1(_0165_),
    .A2(_0167_),
    .B1(wbs_data_o[26]),
    .X(_0168_));
 sky130_fd_sc_hd__and2_4 _0736_ (.A(\configy.counter_d[2] ),
    .B(_0150_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_4 _0737_ (.A(\configy.bits_d[2] ),
    .B(_0152_),
    .X(_0170_));
 sky130_fd_sc_hd__or4_4 _0738_ (.A(_0143_),
    .B(_0146_),
    .C(_0169_),
    .D(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__and3_4 _0739_ (.A(_0163_),
    .B(_0168_),
    .C(_0171_),
    .X(_0102_));
 sky130_fd_sc_hd__a21o_4 _0740_ (.A1(_0165_),
    .A2(_0167_),
    .B1(wbs_data_o[25]),
    .X(_0172_));
 sky130_fd_sc_hd__buf_2 _0741_ (.A(_0142_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_2 _0742_ (.A(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__buf_2 _0743_ (.A(_0145_),
    .X(_0175_));
 sky130_fd_sc_hd__buf_2 _0744_ (.A(\configy.counter_d[1] ),
    .X(_0176_));
 sky130_fd_sc_hd__and2_4 _0745_ (.A(_0176_),
    .B(_0150_),
    .X(_0177_));
 sky130_fd_sc_hd__and2_4 _0746_ (.A(\configy.bits_d[1] ),
    .B(_0152_),
    .X(_0178_));
 sky130_fd_sc_hd__or4_4 _0747_ (.A(_0174_),
    .B(_0175_),
    .C(_0177_),
    .D(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__and3_4 _0748_ (.A(_0163_),
    .B(_0172_),
    .C(_0179_),
    .X(_0101_));
 sky130_fd_sc_hd__a21o_4 _0749_ (.A1(_0165_),
    .A2(_0167_),
    .B1(wbs_data_o[24]),
    .X(_0180_));
 sky130_fd_sc_hd__buf_2 _0750_ (.A(\configy.counter_d[0] ),
    .X(_0181_));
 sky130_fd_sc_hd__buf_2 _0751_ (.A(_0134_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_4 _0752_ (.A(_0181_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__buf_2 _0753_ (.A(_0140_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_4 _0754_ (.A(\configy.bits_d[0] ),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or4_4 _0755_ (.A(_0174_),
    .B(_0175_),
    .C(_0183_),
    .D(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_4 _0756_ (.A(_0163_),
    .B(_0180_),
    .C(_0186_),
    .X(_0100_));
 sky130_fd_sc_hd__a21o_4 _0757_ (.A1(_0165_),
    .A2(_0167_),
    .B1(wbs_data_o[23]),
    .X(_0187_));
 sky130_fd_sc_hd__and2_4 _0758_ (.A(\configy.counter_c[7] ),
    .B(_0182_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_4 _0759_ (.A(\configy.bits_c[7] ),
    .B(_0184_),
    .X(_0189_));
 sky130_fd_sc_hd__or4_4 _0760_ (.A(_0174_),
    .B(_0175_),
    .C(_0188_),
    .D(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__and3_4 _0761_ (.A(_0163_),
    .B(_0187_),
    .C(_0190_),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_4 _0762_ (.A1(_0165_),
    .A2(_0167_),
    .B1(wbs_data_o[22]),
    .X(_0191_));
 sky130_fd_sc_hd__and2_4 _0763_ (.A(\configy.counter_c[6] ),
    .B(_0182_),
    .X(_0192_));
 sky130_fd_sc_hd__and2_4 _0764_ (.A(\configy.bits_c[6] ),
    .B(_0184_),
    .X(_0193_));
 sky130_fd_sc_hd__or4_4 _0765_ (.A(_0174_),
    .B(_0175_),
    .C(_0192_),
    .D(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__and3_4 _0766_ (.A(_0163_),
    .B(_0191_),
    .C(_0194_),
    .X(_0098_));
 sky130_fd_sc_hd__buf_2 _0767_ (.A(_0108_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _0768_ (.A(_0120_),
    .X(_0196_));
 sky130_fd_sc_hd__buf_2 _0769_ (.A(_0129_),
    .X(_0197_));
 sky130_fd_sc_hd__a21o_4 _0770_ (.A1(_0196_),
    .A2(_0197_),
    .B1(wbs_data_o[21]),
    .X(_0198_));
 sky130_fd_sc_hd__buf_2 _0771_ (.A(\configy.counter_c[5] ),
    .X(_0199_));
 sky130_fd_sc_hd__and2_4 _0772_ (.A(_0199_),
    .B(_0182_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_4 _0773_ (.A(\configy.bits_c[5] ),
    .B(_0184_),
    .X(_0201_));
 sky130_fd_sc_hd__or4_4 _0774_ (.A(_0174_),
    .B(_0175_),
    .C(_0200_),
    .D(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__and3_4 _0775_ (.A(_0195_),
    .B(_0198_),
    .C(_0202_),
    .X(_0097_));
 sky130_fd_sc_hd__a21o_4 _0776_ (.A1(_0196_),
    .A2(_0197_),
    .B1(wbs_data_o[20]),
    .X(_0203_));
 sky130_fd_sc_hd__buf_2 _0777_ (.A(_0173_),
    .X(_0204_));
 sky130_fd_sc_hd__buf_2 _0778_ (.A(_0145_),
    .X(_0205_));
 sky130_fd_sc_hd__and2_4 _0779_ (.A(\configy.counter_c[4] ),
    .B(_0182_),
    .X(_0206_));
 sky130_fd_sc_hd__and2_4 _0780_ (.A(\configy.bits_c[4] ),
    .B(_0184_),
    .X(_0207_));
 sky130_fd_sc_hd__or4_4 _0781_ (.A(_0204_),
    .B(_0205_),
    .C(_0206_),
    .D(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__and3_4 _0782_ (.A(_0195_),
    .B(_0203_),
    .C(_0208_),
    .X(_0096_));
 sky130_fd_sc_hd__a21o_4 _0783_ (.A1(_0196_),
    .A2(_0197_),
    .B1(wbs_data_o[19]),
    .X(_0209_));
 sky130_fd_sc_hd__buf_2 _0784_ (.A(_0134_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_4 _0785_ (.A(\configy.counter_c[3] ),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__buf_2 _0786_ (.A(_0140_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_4 _0787_ (.A(\configy.bits_c[3] ),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__or4_4 _0788_ (.A(_0204_),
    .B(_0205_),
    .C(_0211_),
    .D(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_4 _0789_ (.A(_0195_),
    .B(_0209_),
    .C(_0214_),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_4 _0790_ (.A1(_0196_),
    .A2(_0197_),
    .B1(wbs_data_o[18]),
    .X(_0215_));
 sky130_fd_sc_hd__and2_4 _0791_ (.A(\configy.counter_c[2] ),
    .B(_0210_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_4 _0792_ (.A(\configy.bits_c[2] ),
    .B(_0212_),
    .X(_0217_));
 sky130_fd_sc_hd__or4_4 _0793_ (.A(_0204_),
    .B(_0205_),
    .C(_0216_),
    .D(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_4 _0794_ (.A(_0195_),
    .B(_0215_),
    .C(_0218_),
    .X(_0094_));
 sky130_fd_sc_hd__a21o_4 _0795_ (.A1(_0196_),
    .A2(_0197_),
    .B1(wbs_data_o[17]),
    .X(_0219_));
 sky130_fd_sc_hd__buf_2 _0796_ (.A(\configy.counter_c[1] ),
    .X(_0220_));
 sky130_fd_sc_hd__and2_4 _0797_ (.A(_0220_),
    .B(_0210_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_4 _0798_ (.A(\configy.bits_c[1] ),
    .B(_0212_),
    .X(_0222_));
 sky130_fd_sc_hd__or4_4 _0799_ (.A(_0204_),
    .B(_0205_),
    .C(_0221_),
    .D(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_4 _0800_ (.A(_0195_),
    .B(_0219_),
    .C(_0223_),
    .X(_0093_));
 sky130_fd_sc_hd__buf_2 _0801_ (.A(_0108_),
    .X(_0224_));
 sky130_fd_sc_hd__buf_2 _0802_ (.A(_0120_),
    .X(_0225_));
 sky130_fd_sc_hd__buf_2 _0803_ (.A(_0129_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_4 _0804_ (.A1(_0225_),
    .A2(_0226_),
    .B1(wbs_data_o[16]),
    .X(_0227_));
 sky130_fd_sc_hd__buf_2 _0805_ (.A(\configy.counter_c[0] ),
    .X(_0228_));
 sky130_fd_sc_hd__and2_4 _0806_ (.A(_0228_),
    .B(_0210_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_4 _0807_ (.A(\configy.bits_c[0] ),
    .B(_0212_),
    .X(_0230_));
 sky130_fd_sc_hd__or4_4 _0808_ (.A(_0204_),
    .B(_0205_),
    .C(_0229_),
    .D(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_4 _0809_ (.A(_0224_),
    .B(_0227_),
    .C(_0231_),
    .X(_0092_));
 sky130_fd_sc_hd__a21o_4 _0810_ (.A1(_0225_),
    .A2(_0226_),
    .B1(wbs_data_o[15]),
    .X(_0232_));
 sky130_fd_sc_hd__buf_2 _0811_ (.A(_0173_),
    .X(_0233_));
 sky130_fd_sc_hd__buf_2 _0812_ (.A(_0144_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_4 _0813_ (.A(\configy.counter_b[7] ),
    .B(_0210_),
    .X(_0235_));
 sky130_fd_sc_hd__and2_4 _0814_ (.A(\configy.bits_b[7] ),
    .B(_0212_),
    .X(_0236_));
 sky130_fd_sc_hd__or4_4 _0815_ (.A(_0233_),
    .B(_0234_),
    .C(_0235_),
    .D(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__and3_4 _0816_ (.A(_0224_),
    .B(_0232_),
    .C(_0237_),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_4 _0817_ (.A1(_0225_),
    .A2(_0226_),
    .B1(wbs_data_o[14]),
    .X(_0238_));
 sky130_fd_sc_hd__buf_2 _0818_ (.A(_0134_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_4 _0819_ (.A(\configy.counter_b[6] ),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__buf_2 _0820_ (.A(_0139_),
    .X(_0241_));
 sky130_fd_sc_hd__buf_2 _0821_ (.A(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_4 _0822_ (.A(\configy.bits_b[6] ),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__or4_4 _0823_ (.A(_0233_),
    .B(_0234_),
    .C(_0240_),
    .D(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__and3_4 _0824_ (.A(_0224_),
    .B(_0238_),
    .C(_0244_),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_4 _0825_ (.A1(_0225_),
    .A2(_0226_),
    .B1(wbs_data_o[13]),
    .X(_0245_));
 sky130_fd_sc_hd__buf_2 _0826_ (.A(\configy.counter_b[5] ),
    .X(_0246_));
 sky130_fd_sc_hd__and2_4 _0827_ (.A(_0246_),
    .B(_0239_),
    .X(_0247_));
 sky130_fd_sc_hd__and2_4 _0828_ (.A(\configy.bits_b[5] ),
    .B(_0242_),
    .X(_0248_));
 sky130_fd_sc_hd__or4_4 _0829_ (.A(_0233_),
    .B(_0234_),
    .C(_0247_),
    .D(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_4 _0830_ (.A(_0224_),
    .B(_0245_),
    .C(_0249_),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_4 _0831_ (.A1(_0225_),
    .A2(_0226_),
    .B1(wbs_data_o[12]),
    .X(_0250_));
 sky130_fd_sc_hd__and2_4 _0832_ (.A(\configy.counter_b[4] ),
    .B(_0239_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_4 _0833_ (.A(\configy.bits_b[4] ),
    .B(_0242_),
    .X(_0252_));
 sky130_fd_sc_hd__or4_4 _0834_ (.A(_0233_),
    .B(_0234_),
    .C(_0251_),
    .D(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_4 _0835_ (.A(_0224_),
    .B(_0250_),
    .C(_0253_),
    .X(_0088_));
 sky130_fd_sc_hd__buf_2 _0836_ (.A(_0108_),
    .X(_0254_));
 sky130_fd_sc_hd__buf_2 _0837_ (.A(_0120_),
    .X(_0255_));
 sky130_fd_sc_hd__buf_2 _0838_ (.A(_0129_),
    .X(_0256_));
 sky130_fd_sc_hd__a21o_4 _0839_ (.A1(_0255_),
    .A2(_0256_),
    .B1(wbs_data_o[11]),
    .X(_0257_));
 sky130_fd_sc_hd__and2_4 _0840_ (.A(\configy.counter_b[3] ),
    .B(_0239_),
    .X(_0258_));
 sky130_fd_sc_hd__and2_4 _0841_ (.A(\configy.bits_b[3] ),
    .B(_0242_),
    .X(_0259_));
 sky130_fd_sc_hd__or4_4 _0842_ (.A(_0233_),
    .B(_0234_),
    .C(_0258_),
    .D(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__and3_4 _0843_ (.A(_0254_),
    .B(_0257_),
    .C(_0260_),
    .X(_0087_));
 sky130_fd_sc_hd__a21o_4 _0844_ (.A1(_0255_),
    .A2(_0256_),
    .B1(wbs_data_o[10]),
    .X(_0261_));
 sky130_fd_sc_hd__buf_2 _0845_ (.A(_0142_),
    .X(_0262_));
 sky130_fd_sc_hd__buf_2 _0846_ (.A(_0144_),
    .X(_0263_));
 sky130_fd_sc_hd__and2_4 _0847_ (.A(\configy.counter_b[2] ),
    .B(_0239_),
    .X(_0264_));
 sky130_fd_sc_hd__and2_4 _0848_ (.A(\configy.bits_b[2] ),
    .B(_0242_),
    .X(_0265_));
 sky130_fd_sc_hd__or4_4 _0849_ (.A(_0262_),
    .B(_0263_),
    .C(_0264_),
    .D(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__and3_4 _0850_ (.A(_0254_),
    .B(_0261_),
    .C(_0266_),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_4 _0851_ (.A1(_0255_),
    .A2(_0256_),
    .B1(wbs_data_o[9]),
    .X(_0267_));
 sky130_fd_sc_hd__buf_2 _0852_ (.A(\configy.counter_b[1] ),
    .X(_0268_));
 sky130_fd_sc_hd__buf_2 _0853_ (.A(_0133_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_4 _0854_ (.A(_0268_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__buf_2 _0855_ (.A(_0241_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_4 _0856_ (.A(\configy.bits_b[1] ),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or4_4 _0857_ (.A(_0262_),
    .B(_0263_),
    .C(_0270_),
    .D(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__and3_4 _0858_ (.A(_0254_),
    .B(_0267_),
    .C(_0273_),
    .X(_0085_));
 sky130_fd_sc_hd__a21o_4 _0859_ (.A1(_0255_),
    .A2(_0256_),
    .B1(wbs_data_o[8]),
    .X(_0274_));
 sky130_fd_sc_hd__buf_2 _0860_ (.A(\configy.counter_b[0] ),
    .X(_0275_));
 sky130_fd_sc_hd__and2_4 _0861_ (.A(_0275_),
    .B(_0269_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_4 _0862_ (.A(\configy.bits_b[0] ),
    .B(_0271_),
    .X(_0277_));
 sky130_fd_sc_hd__or4_4 _0863_ (.A(_0262_),
    .B(_0263_),
    .C(_0276_),
    .D(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__and3_4 _0864_ (.A(_0254_),
    .B(_0274_),
    .C(_0278_),
    .X(_0084_));
 sky130_fd_sc_hd__a21o_4 _0865_ (.A1(_0255_),
    .A2(_0256_),
    .B1(wbs_data_o[7]),
    .X(_0279_));
 sky130_fd_sc_hd__and2_4 _0866_ (.A(\configy.counter_a[7] ),
    .B(_0269_),
    .X(_0280_));
 sky130_fd_sc_hd__and2_4 _0867_ (.A(\configy.bits_a[7] ),
    .B(_0271_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_4 _0868_ (.A(_0262_),
    .B(_0263_),
    .C(_0280_),
    .D(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__and3_4 _0869_ (.A(_0254_),
    .B(_0279_),
    .C(_0282_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_2 _0870_ (.A(_0108_),
    .X(_0283_));
 sky130_fd_sc_hd__buf_2 _0871_ (.A(_0120_),
    .X(_0284_));
 sky130_fd_sc_hd__buf_2 _0872_ (.A(_0129_),
    .X(_0285_));
 sky130_fd_sc_hd__a21o_4 _0873_ (.A1(_0284_),
    .A2(_0285_),
    .B1(wbs_data_o[6]),
    .X(_0286_));
 sky130_fd_sc_hd__and2_4 _0874_ (.A(\configy.counter_a[6] ),
    .B(_0269_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_4 _0875_ (.A(\configy.bits_a[6] ),
    .B(_0271_),
    .X(_0288_));
 sky130_fd_sc_hd__or4_4 _0876_ (.A(_0262_),
    .B(_0263_),
    .C(_0287_),
    .D(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__and3_4 _0877_ (.A(_0283_),
    .B(_0286_),
    .C(_0289_),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_4 _0878_ (.A1(_0284_),
    .A2(_0285_),
    .B1(wbs_data_o[5]),
    .X(_0290_));
 sky130_fd_sc_hd__buf_2 _0879_ (.A(_0142_),
    .X(_0291_));
 sky130_fd_sc_hd__buf_2 _0880_ (.A(_0144_),
    .X(_0292_));
 sky130_fd_sc_hd__buf_2 _0881_ (.A(\configy.counter_a[5] ),
    .X(_0293_));
 sky130_fd_sc_hd__and2_4 _0882_ (.A(_0293_),
    .B(_0269_),
    .X(_0294_));
 sky130_fd_sc_hd__and2_4 _0883_ (.A(\configy.bits_a[5] ),
    .B(_0271_),
    .X(_0295_));
 sky130_fd_sc_hd__or4_4 _0884_ (.A(_0291_),
    .B(_0292_),
    .C(_0294_),
    .D(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__and3_4 _0885_ (.A(_0283_),
    .B(_0290_),
    .C(_0296_),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_4 _0886_ (.A1(_0284_),
    .A2(_0285_),
    .B1(wbs_data_o[4]),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _0887_ (.A(_0133_),
    .X(_0298_));
 sky130_fd_sc_hd__and2_4 _0888_ (.A(\configy.counter_a[4] ),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _0889_ (.A(_0241_),
    .X(_0300_));
 sky130_fd_sc_hd__and2_4 _0890_ (.A(\configy.bits_a[4] ),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or4_4 _0891_ (.A(_0291_),
    .B(_0292_),
    .C(_0299_),
    .D(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__and3_4 _0892_ (.A(_0283_),
    .B(_0297_),
    .C(_0302_),
    .X(_0080_));
 sky130_fd_sc_hd__a21o_4 _0893_ (.A1(_0284_),
    .A2(_0285_),
    .B1(wbs_data_o[3]),
    .X(_0303_));
 sky130_fd_sc_hd__and2_4 _0894_ (.A(\configy.counter_a[3] ),
    .B(_0298_),
    .X(_0304_));
 sky130_fd_sc_hd__and2_4 _0895_ (.A(\configy.bits_a[3] ),
    .B(_0300_),
    .X(_0305_));
 sky130_fd_sc_hd__or4_4 _0896_ (.A(_0291_),
    .B(_0292_),
    .C(_0304_),
    .D(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__and3_4 _0897_ (.A(_0283_),
    .B(_0303_),
    .C(_0306_),
    .X(_0079_));
 sky130_fd_sc_hd__a21o_4 _0898_ (.A1(_0284_),
    .A2(_0285_),
    .B1(wbs_data_o[2]),
    .X(_0307_));
 sky130_fd_sc_hd__and2_4 _0899_ (.A(\configy.counter_a[2] ),
    .B(_0298_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_4 _0900_ (.A(\configy.bits_a[2] ),
    .B(_0300_),
    .X(_0309_));
 sky130_fd_sc_hd__or4_4 _0901_ (.A(_0291_),
    .B(_0292_),
    .C(_0308_),
    .D(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and3_4 _0902_ (.A(_0283_),
    .B(_0307_),
    .C(_0310_),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_4 _0903_ (.A1(_0164_),
    .A2(_0166_),
    .B1(wbs_data_o[1]),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _0904_ (.A(\configy.counter_a[1] ),
    .X(_0312_));
 sky130_fd_sc_hd__and2_4 _0905_ (.A(_0312_),
    .B(_0298_),
    .X(_0313_));
 sky130_fd_sc_hd__and2_4 _0906_ (.A(\configy.bits_a[1] ),
    .B(_0300_),
    .X(_0314_));
 sky130_fd_sc_hd__or4_4 _0907_ (.A(_0291_),
    .B(_0292_),
    .C(_0313_),
    .D(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__and3_4 _0908_ (.A(_0109_),
    .B(_0311_),
    .C(_0315_),
    .X(_0077_));
 sky130_fd_sc_hd__a21o_4 _0909_ (.A1(_0164_),
    .A2(_0166_),
    .B1(wbs_data_o[0]),
    .X(_0316_));
 sky130_fd_sc_hd__and2_4 _0910_ (.A(\configy.bits_a[0] ),
    .B(_0140_),
    .X(_0317_));
 sky130_fd_sc_hd__and2_4 _0911_ (.A(_0138_),
    .B(_0132_),
    .X(_0318_));
 sky130_fd_sc_hd__buf_2 _0912_ (.A(\configy.counter_a[0] ),
    .X(_0319_));
 sky130_fd_sc_hd__and3_4 _0913_ (.A(_0319_),
    .B(wbs_addr_i[3]),
    .C(_0132_),
    .X(_0320_));
 sky130_fd_sc_hd__a21o_4 _0914_ (.A1(\configy.free_run ),
    .A2(_0318_),
    .B1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__or4_4 _0915_ (.A(_0173_),
    .B(_0145_),
    .C(_0317_),
    .D(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__and3_4 _0916_ (.A(_0109_),
    .B(_0316_),
    .C(_0322_),
    .X(_0076_));
 sky130_fd_sc_hd__buf_2 _0917_ (.A(wb_rst_i),
    .X(_0323_));
 sky130_fd_sc_hd__buf_2 _0918_ (.A(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a21oi_4 _0919_ (.A1(_0121_),
    .A2(_0130_),
    .B1(\configy.read_transaction_in_progress ),
    .Y(_0325_));
 sky130_fd_sc_hd__buf_2 _0920_ (.A(\configy.write_transaction_in_progress ),
    .X(_0326_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__and2_4 _0922_ (.A(\configy.read_transaction_in_progress ),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__nor3_4 _0923_ (.A(_0324_),
    .B(_0325_),
    .C(_0328_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(wbs_data_i[0]),
    .Y(_0329_));
 sky130_fd_sc_hd__buf_2 _0925_ (.A(wbs_sel_i[0]),
    .X(_0330_));
 sky130_fd_sc_hd__and4_4 _0926_ (.A(_0138_),
    .B(_0330_),
    .C(_0326_),
    .D(_0132_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_2 _0927_ (.A(wb_rst_i),
    .X(_0332_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__o21ai_4 _0929_ (.A1(\configy.free_run ),
    .A2(_0331_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21oi_4 _0930_ (.A1(_0329_),
    .A2(_0331_),
    .B1(_0334_),
    .Y(_0074_));
 sky130_fd_sc_hd__and3_4 _0931_ (.A(wbs_addr_i[3]),
    .B(\configy.write_transaction_in_progress ),
    .C(_0132_),
    .X(_0335_));
 sky130_fd_sc_hd__buf_2 _0932_ (.A(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_4 _0933_ (.A(wbs_sel_i[3]),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__buf_2 _0934_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__buf_2 _0935_ (.A(\configy.output_initiated ),
    .X(_0339_));
 sky130_fd_sc_hd__buf_2 _0936_ (.A(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__buf_2 _0937_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_2 _0938_ (.A(_0336_),
    .X(_0342_));
 sky130_fd_sc_hd__and4_4 _0939_ (.A(\configy.charged[3] ),
    .B(\configy.charged[2] ),
    .C(\configy.charged[1] ),
    .D(\configy.charged[0] ),
    .X(_0343_));
 sky130_fd_sc_hd__or2_4 _0940_ (.A(wb_rst_i),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__a21oi_4 _0941_ (.A1(_0341_),
    .A2(_0342_),
    .B1(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__o21a_4 _0942_ (.A1(\configy.charged[3] ),
    .A2(_0338_),
    .B1(_0345_),
    .X(_0073_));
 sky130_fd_sc_hd__and2_4 _0943_ (.A(wbs_sel_i[2]),
    .B(_0336_),
    .X(_0346_));
 sky130_fd_sc_hd__buf_2 _0944_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__o21a_4 _0945_ (.A1(\configy.charged[2] ),
    .A2(_0347_),
    .B1(_0345_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_4 _0946_ (.A(wbs_sel_i[1]),
    .B(_0335_),
    .X(_0348_));
 sky130_fd_sc_hd__buf_2 _0947_ (.A(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__o21a_4 _0948_ (.A1(\configy.charged[1] ),
    .A2(_0349_),
    .B1(_0345_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_4 _0949_ (.A(_0330_),
    .B(_0335_),
    .X(_0350_));
 sky130_fd_sc_hd__buf_2 _0950_ (.A(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__o21a_4 _0951_ (.A1(\configy.charged[0] ),
    .A2(_0351_),
    .B1(_0345_),
    .X(_0070_));
 sky130_fd_sc_hd__buf_2 _0952_ (.A(\configy.bits_index[2] ),
    .X(_0352_));
 sky130_fd_sc_hd__buf_2 _0953_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_4 _0954_ (.A(\configy.bits_index[1] ),
    .B(\configy.bits_index[0] ),
    .X(_0354_));
 sky130_fd_sc_hd__or2_4 _0955_ (.A(_0353_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_4 _0956_ (.A(_0353_),
    .B(_0354_),
    .X(_0356_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__buf_2 _0958_ (.A(\configy.output_initiated ),
    .X(_0358_));
 sky130_fd_sc_hd__buf_2 _0959_ (.A(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__buf_2 _0960_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nor2_4 _0961_ (.A(_0360_),
    .B(_0336_),
    .Y(_0361_));
 sky130_fd_sc_hd__a32o_4 _0962_ (.A1(_0341_),
    .A2(_0355_),
    .A3(_0357_),
    .B1(_0361_),
    .B2(_0353_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_4 _0963_ (.A(_0333_),
    .B(_0362_),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _0964_ (.A(\configy.output_initiated ),
    .Y(_0363_));
 sky130_fd_sc_hd__buf_2 _0965_ (.A(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__buf_2 _0966_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_2 _0967_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__buf_2 _0968_ (.A(\configy.bits_index[1] ),
    .X(_0367_));
 sky130_fd_sc_hd__a2bb2o_4 _0969_ (.A1_N(_0366_),
    .A2_N(_0354_),
    .B1(_0361_),
    .B2(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(\configy.bits_index[1] ),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(\configy.bits_index[0] ),
    .Y(_0370_));
 sky130_fd_sc_hd__and2_4 _0972_ (.A(_0369_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_4 _0973_ (.A(_0323_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__and2_4 _0974_ (.A(_0368_),
    .B(_0372_),
    .X(_0068_));
 sky130_fd_sc_hd__buf_2 _0975_ (.A(_0370_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_4 _0976_ (.A(_0373_),
    .B(_0361_),
    .X(_0374_));
 sky130_fd_sc_hd__buf_2 _0977_ (.A(\configy.bits_index[0] ),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _0978_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__or2_4 _0979_ (.A(_0376_),
    .B(_0341_),
    .X(_0377_));
 sky130_fd_sc_hd__and3_4 _0980_ (.A(_0333_),
    .B(_0374_),
    .C(_0377_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_2 _0981_ (.A(_0358_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_4 _0982_ (.A(wbs_data_i[7]),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__or4_4 _0983_ (.A(\configy.counter_a[3] ),
    .B(\configy.counter_a[2] ),
    .C(\configy.counter_a[1] ),
    .D(\configy.counter_a[0] ),
    .X(_0380_));
 sky130_fd_sc_hd__or4_4 _0984_ (.A(\configy.counter_a[6] ),
    .B(_0293_),
    .C(\configy.counter_a[4] ),
    .D(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__buf_2 _0985_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__and4_4 _0986_ (.A(\configy.counter_a[5] ),
    .B(\configy.counter_a[4] ),
    .C(\configy.counter_a[3] ),
    .D(\configy.counter_a[2] ),
    .X(_0383_));
 sky130_fd_sc_hd__and4_4 _0987_ (.A(\configy.counter_a[7] ),
    .B(\configy.counter_a[6] ),
    .C(\configy.counter_a[1] ),
    .D(\configy.counter_a[0] ),
    .X(_0384_));
 sky130_fd_sc_hd__buf_2 _0988_ (.A(_0364_),
    .X(_0385_));
 sky130_fd_sc_hd__a21oi_4 _0989_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a41oi_4 _0990_ (.A1(_0330_),
    .A2(_0326_),
    .A3(_0365_),
    .A4(_0241_),
    .B1(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__buf_2 _0991_ (.A(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a21o_4 _0992_ (.A1(_0379_),
    .A2(_0382_),
    .B1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__buf_2 _0993_ (.A(\configy.write_transaction_in_progress ),
    .X(_0390_));
 sky130_fd_sc_hd__buf_2 _0994_ (.A(_0363_),
    .X(_0391_));
 sky130_fd_sc_hd__buf_2 _0995_ (.A(_0139_),
    .X(_0392_));
 sky130_fd_sc_hd__a41o_4 _0996_ (.A1(wbs_sel_i[0]),
    .A2(_0390_),
    .A3(_0391_),
    .A4(_0392_),
    .B1(_0386_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_2 _0997_ (.A(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_4 _0998_ (.A1(\configy.counter_a[7] ),
    .A2(_0382_),
    .B1(_0360_),
    .Y(_0395_));
 sky130_fd_sc_hd__and3_4 _0999_ (.A(_0394_),
    .B(_0379_),
    .C(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__buf_2 _1000_ (.A(_0332_),
    .X(_0397_));
 sky130_fd_sc_hd__a211o_4 _1001_ (.A1(\configy.counter_a[7] ),
    .A2(_0389_),
    .B1(_0396_),
    .C1(_0397_),
    .X(_0066_));
 sky130_fd_sc_hd__buf_2 _1002_ (.A(_0358_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_2 _1003_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_4 _1004_ (.A(_0399_),
    .B(_0382_),
    .Y(_0400_));
 sky130_fd_sc_hd__buf_2 _1005_ (.A(_0358_),
    .X(_0401_));
 sky130_fd_sc_hd__or2_4 _1006_ (.A(wbs_data_i[6]),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and3_4 _1007_ (.A(_0393_),
    .B(_0400_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__or2_4 _1008_ (.A(\configy.counter_a[4] ),
    .B(_0380_),
    .X(_0404_));
 sky130_fd_sc_hd__o21a_4 _1009_ (.A1(_0293_),
    .A2(_0404_),
    .B1(_0378_),
    .X(_0405_));
 sky130_fd_sc_hd__o21a_4 _1010_ (.A1(_0387_),
    .A2(_0405_),
    .B1(\configy.counter_a[6] ),
    .X(_0406_));
 sky130_fd_sc_hd__or3_4 _1011_ (.A(_0323_),
    .B(_0403_),
    .C(_0406_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_2 _1012_ (.A(_0340_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_4 _1013_ (.A(wbs_data_i[5]),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__a2bb2o_4 _1014_ (.A1_N(_0387_),
    .A2_N(_0405_),
    .B1(_0404_),
    .B2(_0293_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_4 _1015_ (.A(_0293_),
    .B(_0388_),
    .X(_0410_));
 sky130_fd_sc_hd__a211o_4 _1016_ (.A1(_0408_),
    .A2(_0409_),
    .B1(_0410_),
    .C1(_0397_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_4 _1017_ (.A(_0407_),
    .B(_0380_),
    .Y(_0411_));
 sky130_fd_sc_hd__nand2_4 _1018_ (.A(_0394_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_4 _1019_ (.A(_0360_),
    .B(_0404_),
    .Y(_0413_));
 sky130_fd_sc_hd__buf_2 _1020_ (.A(_0339_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_4 _1021_ (.A(wbs_data_i[4]),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__and3_4 _1022_ (.A(_0394_),
    .B(_0413_),
    .C(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__a211o_4 _1023_ (.A1(\configy.counter_a[4] ),
    .A2(_0412_),
    .B1(_0416_),
    .C1(_0397_),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_4 _1024_ (.A1(_0394_),
    .A2(_0411_),
    .B1(\configy.counter_a[3] ),
    .X(_0417_));
 sky130_fd_sc_hd__buf_2 _1025_ (.A(_0398_),
    .X(_0418_));
 sky130_fd_sc_hd__or4_4 _1026_ (.A(\configy.counter_a[2] ),
    .B(_0312_),
    .C(\configy.counter_a[0] ),
    .D(_0385_),
    .X(_0419_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(\configy.counter_a[3] ),
    .Y(_0420_));
 sky130_fd_sc_hd__o22a_4 _1028_ (.A1(wbs_data_i[3]),
    .A2(_0418_),
    .B1(_0419_),
    .B2(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__or2_4 _1029_ (.A(_0388_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__a21o_4 _1030_ (.A1(_0417_),
    .A2(_0422_),
    .B1(_0324_),
    .X(_0062_));
 sky130_fd_sc_hd__a21bo_4 _1031_ (.A1(wbs_data_i[2]),
    .A2(_0366_),
    .B1_N(_0419_),
    .X(_0423_));
 sky130_fd_sc_hd__o21a_4 _1032_ (.A1(_0312_),
    .A2(_0319_),
    .B1(_0339_),
    .X(_0424_));
 sky130_fd_sc_hd__o21a_4 _1033_ (.A1(_0387_),
    .A2(_0424_),
    .B1(\configy.counter_a[2] ),
    .X(_0425_));
 sky130_fd_sc_hd__a211o_4 _1034_ (.A1(_0394_),
    .A2(_0423_),
    .B1(_0425_),
    .C1(_0397_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_2 _1035_ (.A(_0398_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_4 _1036_ (.A(wbs_data_i[1]),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__a21bo_4 _1037_ (.A1(_0312_),
    .A2(_0319_),
    .B1_N(_0424_),
    .X(_0428_));
 sky130_fd_sc_hd__and3_4 _1038_ (.A(_0393_),
    .B(_0427_),
    .C(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a211o_4 _1039_ (.A1(_0312_),
    .A2(_0388_),
    .B1(_0429_),
    .C1(_0397_),
    .X(_0060_));
 sky130_fd_sc_hd__or2_4 _1040_ (.A(wbs_data_i[0]),
    .B(_0426_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_2 _1041_ (.A(_0401_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_4 _1042_ (.A(_0319_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__and3_4 _1043_ (.A(_0393_),
    .B(_0430_),
    .C(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_2 _1044_ (.A(_0332_),
    .X(_0434_));
 sky130_fd_sc_hd__a211o_4 _1045_ (.A1(_0319_),
    .A2(_0388_),
    .B1(_0433_),
    .C1(_0434_),
    .X(_0059_));
 sky130_fd_sc_hd__or4_4 _1046_ (.A(\configy.counter_b[3] ),
    .B(\configy.counter_b[2] ),
    .C(\configy.counter_b[1] ),
    .D(\configy.counter_b[0] ),
    .X(_0435_));
 sky130_fd_sc_hd__or4_4 _1047_ (.A(\configy.counter_b[6] ),
    .B(_0246_),
    .C(\configy.counter_b[4] ),
    .D(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__buf_2 _1048_ (.A(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__or2_4 _1049_ (.A(wbs_data_i[15]),
    .B(_0359_),
    .X(_0438_));
 sky130_fd_sc_hd__and4_4 _1050_ (.A(\configy.counter_b[5] ),
    .B(\configy.counter_b[4] ),
    .C(\configy.counter_b[3] ),
    .D(\configy.counter_b[2] ),
    .X(_0439_));
 sky130_fd_sc_hd__and4_4 _1051_ (.A(\configy.counter_b[7] ),
    .B(\configy.counter_b[6] ),
    .C(\configy.counter_b[1] ),
    .D(\configy.counter_b[0] ),
    .X(_0440_));
 sky130_fd_sc_hd__a21oi_4 _1052_ (.A1(_0439_),
    .A2(_0440_),
    .B1(_0364_),
    .Y(_0441_));
 sky130_fd_sc_hd__a41oi_4 _1053_ (.A1(_0390_),
    .A2(_0391_),
    .A3(wbs_sel_i[1]),
    .A4(_0392_),
    .B1(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__buf_2 _1054_ (.A(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__a21o_4 _1055_ (.A1(_0437_),
    .A2(_0438_),
    .B1(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a41o_4 _1056_ (.A1(\configy.write_transaction_in_progress ),
    .A2(_0391_),
    .A3(wbs_sel_i[1]),
    .A4(_0139_),
    .B1(_0441_),
    .X(_0445_));
 sky130_fd_sc_hd__buf_2 _1057_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__o21ai_4 _1058_ (.A1(\configy.counter_b[7] ),
    .A2(_0437_),
    .B1(_0431_),
    .Y(_0447_));
 sky130_fd_sc_hd__and3_4 _1059_ (.A(_0446_),
    .B(_0438_),
    .C(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__a211o_4 _1060_ (.A1(\configy.counter_b[7] ),
    .A2(_0444_),
    .B1(_0448_),
    .C1(_0434_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_2 _1061_ (.A(wb_rst_i),
    .X(_0449_));
 sky130_fd_sc_hd__nand2_4 _1062_ (.A(_0399_),
    .B(_0437_),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_4 _1063_ (.A(wbs_data_i[14]),
    .B(_0401_),
    .X(_0451_));
 sky130_fd_sc_hd__and3_4 _1064_ (.A(_0446_),
    .B(_0450_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or2_4 _1065_ (.A(\configy.counter_b[4] ),
    .B(_0435_),
    .X(_0453_));
 sky130_fd_sc_hd__o21a_4 _1066_ (.A1(_0246_),
    .A2(_0453_),
    .B1(_0378_),
    .X(_0454_));
 sky130_fd_sc_hd__o21a_4 _1067_ (.A1(_0443_),
    .A2(_0454_),
    .B1(\configy.counter_b[6] ),
    .X(_0455_));
 sky130_fd_sc_hd__or3_4 _1068_ (.A(_0449_),
    .B(_0452_),
    .C(_0455_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_4 _1069_ (.A(wbs_data_i[13]),
    .B(_0407_),
    .X(_0456_));
 sky130_fd_sc_hd__a2bb2o_4 _1070_ (.A1_N(_0443_),
    .A2_N(_0454_),
    .B1(_0453_),
    .B2(_0246_),
    .X(_0457_));
 sky130_fd_sc_hd__buf_2 _1071_ (.A(_0442_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_4 _1072_ (.A(_0246_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a211o_4 _1073_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0459_),
    .C1(_0434_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_4 _1074_ (.A(_0418_),
    .B(_0453_),
    .Y(_0460_));
 sky130_fd_sc_hd__or2_4 _1075_ (.A(wbs_data_i[12]),
    .B(_0401_),
    .X(_0461_));
 sky130_fd_sc_hd__and3_4 _1076_ (.A(_0445_),
    .B(_0460_),
    .C(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and2_4 _1077_ (.A(_0340_),
    .B(_0435_),
    .X(_0463_));
 sky130_fd_sc_hd__o21a_4 _1078_ (.A1(_0443_),
    .A2(_0463_),
    .B1(\configy.counter_b[4] ),
    .X(_0464_));
 sky130_fd_sc_hd__or3_4 _1079_ (.A(_0449_),
    .B(_0462_),
    .C(_0464_),
    .X(_0055_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(\configy.counter_b[3] ),
    .Y(_0465_));
 sky130_fd_sc_hd__o21ai_4 _1081_ (.A1(_0458_),
    .A2(_0463_),
    .B1(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__or4_4 _1082_ (.A(\configy.counter_b[2] ),
    .B(_0268_),
    .C(\configy.counter_b[0] ),
    .D(_0385_),
    .X(_0467_));
 sky130_fd_sc_hd__o22a_4 _1083_ (.A1(wbs_data_i[11]),
    .A2(_0418_),
    .B1(_0467_),
    .B2(_0465_),
    .X(_0468_));
 sky130_fd_sc_hd__or2_4 _1084_ (.A(_0458_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a21o_4 _1085_ (.A1(_0466_),
    .A2(_0469_),
    .B1(_0324_),
    .X(_0054_));
 sky130_fd_sc_hd__a21bo_4 _1086_ (.A1(wbs_data_i[10]),
    .A2(_0366_),
    .B1_N(_0467_),
    .X(_0470_));
 sky130_fd_sc_hd__o21a_4 _1087_ (.A1(_0268_),
    .A2(_0275_),
    .B1(_0339_),
    .X(_0471_));
 sky130_fd_sc_hd__o21a_4 _1088_ (.A1(_0443_),
    .A2(_0471_),
    .B1(\configy.counter_b[2] ),
    .X(_0472_));
 sky130_fd_sc_hd__a211o_4 _1089_ (.A1(_0446_),
    .A2(_0470_),
    .B1(_0472_),
    .C1(_0434_),
    .X(_0053_));
 sky130_fd_sc_hd__or2_4 _1090_ (.A(wbs_data_i[9]),
    .B(_0426_),
    .X(_0473_));
 sky130_fd_sc_hd__a21bo_4 _1091_ (.A1(_0268_),
    .A2(_0275_),
    .B1_N(_0471_),
    .X(_0474_));
 sky130_fd_sc_hd__and3_4 _1092_ (.A(_0446_),
    .B(_0473_),
    .C(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__a211o_4 _1093_ (.A1(_0268_),
    .A2(_0458_),
    .B1(_0475_),
    .C1(_0434_),
    .X(_0052_));
 sky130_fd_sc_hd__or2_4 _1094_ (.A(wbs_data_i[8]),
    .B(_0426_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_4 _1095_ (.A(_0275_),
    .B(_0431_),
    .Y(_0477_));
 sky130_fd_sc_hd__and3_4 _1096_ (.A(_0446_),
    .B(_0476_),
    .C(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_2 _1097_ (.A(_0332_),
    .X(_0479_));
 sky130_fd_sc_hd__a211o_4 _1098_ (.A1(_0275_),
    .A2(_0458_),
    .B1(_0478_),
    .C1(_0479_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_4 _1099_ (.A(wbs_data_i[23]),
    .B(_0378_),
    .X(_0480_));
 sky130_fd_sc_hd__or4_4 _1100_ (.A(\configy.counter_c[3] ),
    .B(\configy.counter_c[2] ),
    .C(\configy.counter_c[1] ),
    .D(\configy.counter_c[0] ),
    .X(_0481_));
 sky130_fd_sc_hd__or4_4 _1101_ (.A(\configy.counter_c[6] ),
    .B(_0199_),
    .C(\configy.counter_c[4] ),
    .D(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_2 _1102_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__and4_4 _1103_ (.A(\configy.counter_c[5] ),
    .B(\configy.counter_c[4] ),
    .C(\configy.counter_c[3] ),
    .D(\configy.counter_c[2] ),
    .X(_0484_));
 sky130_fd_sc_hd__and4_4 _1104_ (.A(\configy.counter_c[7] ),
    .B(\configy.counter_c[6] ),
    .C(\configy.counter_c[1] ),
    .D(\configy.counter_c[0] ),
    .X(_0485_));
 sky130_fd_sc_hd__a21oi_4 _1105_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_0385_),
    .Y(_0486_));
 sky130_fd_sc_hd__a41oi_4 _1106_ (.A1(_0326_),
    .A2(_0365_),
    .A3(wbs_sel_i[2]),
    .A4(_0241_),
    .B1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__buf_2 _1107_ (.A(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_4 _1108_ (.A1(_0480_),
    .A2(_0483_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a41o_4 _1109_ (.A1(_0390_),
    .A2(_0365_),
    .A3(wbs_sel_i[2]),
    .A4(_0392_),
    .B1(_0486_),
    .X(_0490_));
 sky130_fd_sc_hd__buf_2 _1110_ (.A(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o21ai_4 _1111_ (.A1(\configy.counter_c[7] ),
    .A2(_0483_),
    .B1(_0431_),
    .Y(_0492_));
 sky130_fd_sc_hd__and3_4 _1112_ (.A(_0491_),
    .B(_0480_),
    .C(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__a211o_4 _1113_ (.A1(\configy.counter_c[7] ),
    .A2(_0489_),
    .B1(_0493_),
    .C1(_0479_),
    .X(_0050_));
 sky130_fd_sc_hd__nand2_4 _1114_ (.A(_0418_),
    .B(_0483_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_4 _1115_ (.A(wbs_data_i[22]),
    .B(_0398_),
    .X(_0495_));
 sky130_fd_sc_hd__and3_4 _1116_ (.A(_0490_),
    .B(_0494_),
    .C(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__or2_4 _1117_ (.A(\configy.counter_c[4] ),
    .B(_0481_),
    .X(_0497_));
 sky130_fd_sc_hd__o21a_4 _1118_ (.A1(_0199_),
    .A2(_0497_),
    .B1(_0359_),
    .X(_0498_));
 sky130_fd_sc_hd__o21a_4 _1119_ (.A1(_0487_),
    .A2(_0498_),
    .B1(\configy.counter_c[6] ),
    .X(_0499_));
 sky130_fd_sc_hd__or3_4 _1120_ (.A(_0449_),
    .B(_0496_),
    .C(_0499_),
    .X(_0049_));
 sky130_fd_sc_hd__or2_4 _1121_ (.A(wbs_data_i[21]),
    .B(_0407_),
    .X(_0500_));
 sky130_fd_sc_hd__a2bb2o_4 _1122_ (.A1_N(_0487_),
    .A2_N(_0498_),
    .B1(_0497_),
    .B2(_0199_),
    .X(_0501_));
 sky130_fd_sc_hd__and2_4 _1123_ (.A(_0199_),
    .B(_0488_),
    .X(_0502_));
 sky130_fd_sc_hd__a211o_4 _1124_ (.A1(_0500_),
    .A2(_0501_),
    .B1(_0502_),
    .C1(_0479_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_4 _1125_ (.A(_0407_),
    .B(_0481_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_4 _1126_ (.A(_0491_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_4 _1127_ (.A(_0360_),
    .B(_0497_),
    .Y(_0505_));
 sky130_fd_sc_hd__or2_4 _1128_ (.A(wbs_data_i[20]),
    .B(_0378_),
    .X(_0506_));
 sky130_fd_sc_hd__and3_4 _1129_ (.A(_0491_),
    .B(_0505_),
    .C(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a211o_4 _1130_ (.A1(\configy.counter_c[4] ),
    .A2(_0504_),
    .B1(_0507_),
    .C1(_0479_),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_4 _1131_ (.A1(_0491_),
    .A2(_0503_),
    .B1(\configy.counter_c[3] ),
    .X(_0508_));
 sky130_fd_sc_hd__or4_4 _1132_ (.A(\configy.counter_c[2] ),
    .B(_0220_),
    .C(\configy.counter_c[0] ),
    .D(_0385_),
    .X(_0509_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(\configy.counter_c[3] ),
    .Y(_0510_));
 sky130_fd_sc_hd__o22a_4 _1134_ (.A1(wbs_data_i[19]),
    .A2(_0340_),
    .B1(_0509_),
    .B2(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_4 _1135_ (.A(_0488_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a21o_4 _1136_ (.A1(_0508_),
    .A2(_0512_),
    .B1(_0324_),
    .X(_0046_));
 sky130_fd_sc_hd__a21bo_4 _1137_ (.A1(wbs_data_i[18]),
    .A2(_0366_),
    .B1_N(_0509_),
    .X(_0513_));
 sky130_fd_sc_hd__o21a_4 _1138_ (.A1(_0220_),
    .A2(_0228_),
    .B1(_0339_),
    .X(_0514_));
 sky130_fd_sc_hd__o21a_4 _1139_ (.A1(_0487_),
    .A2(_0514_),
    .B1(\configy.counter_c[2] ),
    .X(_0515_));
 sky130_fd_sc_hd__a211o_4 _1140_ (.A1(_0491_),
    .A2(_0513_),
    .B1(_0515_),
    .C1(_0479_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_4 _1141_ (.A(wbs_data_i[17]),
    .B(_0414_),
    .X(_0516_));
 sky130_fd_sc_hd__a21bo_4 _1142_ (.A1(_0220_),
    .A2(_0228_),
    .B1_N(_0514_),
    .X(_0517_));
 sky130_fd_sc_hd__and3_4 _1143_ (.A(_0490_),
    .B(_0516_),
    .C(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_2 _1144_ (.A(_0332_),
    .X(_0519_));
 sky130_fd_sc_hd__a211o_4 _1145_ (.A1(_0220_),
    .A2(_0488_),
    .B1(_0518_),
    .C1(_0519_),
    .X(_0044_));
 sky130_fd_sc_hd__or2_4 _1146_ (.A(wbs_data_i[16]),
    .B(_0414_),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_4 _1147_ (.A(_0228_),
    .B(_0399_),
    .Y(_0521_));
 sky130_fd_sc_hd__and3_4 _1148_ (.A(_0490_),
    .B(_0520_),
    .C(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__a211o_4 _1149_ (.A1(_0228_),
    .A2(_0488_),
    .B1(_0522_),
    .C1(_0519_),
    .X(_0043_));
 sky130_fd_sc_hd__or4_4 _1150_ (.A(\configy.counter_d[3] ),
    .B(\configy.counter_d[2] ),
    .C(\configy.counter_d[1] ),
    .D(\configy.counter_d[0] ),
    .X(_0523_));
 sky130_fd_sc_hd__or4_4 _1151_ (.A(\configy.counter_d[6] ),
    .B(_0149_),
    .C(\configy.counter_d[4] ),
    .D(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__buf_2 _1152_ (.A(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_4 _1153_ (.A(wbs_data_i[31]),
    .B(_0401_),
    .X(_0526_));
 sky130_fd_sc_hd__and4_4 _1154_ (.A(\configy.counter_d[5] ),
    .B(\configy.counter_d[4] ),
    .C(\configy.counter_d[3] ),
    .D(\configy.counter_d[2] ),
    .X(_0527_));
 sky130_fd_sc_hd__and4_4 _1155_ (.A(\configy.counter_d[7] ),
    .B(\configy.counter_d[6] ),
    .C(\configy.counter_d[1] ),
    .D(\configy.counter_d[0] ),
    .X(_0528_));
 sky130_fd_sc_hd__a21oi_4 _1156_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0364_),
    .Y(_0529_));
 sky130_fd_sc_hd__a41oi_4 _1157_ (.A1(_0390_),
    .A2(_0391_),
    .A3(wbs_sel_i[3]),
    .A4(_0392_),
    .B1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__buf_2 _1158_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_4 _1159_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__a41o_4 _1160_ (.A1(_0390_),
    .A2(_0391_),
    .A3(wbs_sel_i[3]),
    .A4(_0392_),
    .B1(_0529_),
    .X(_0533_));
 sky130_fd_sc_hd__buf_2 _1161_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__o21ai_4 _1162_ (.A1(\configy.counter_d[7] ),
    .A2(_0525_),
    .B1(_0431_),
    .Y(_0535_));
 sky130_fd_sc_hd__and3_4 _1163_ (.A(_0534_),
    .B(_0526_),
    .C(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a211o_4 _1164_ (.A1(\configy.counter_d[7] ),
    .A2(_0532_),
    .B1(_0536_),
    .C1(_0519_),
    .X(_0042_));
 sky130_fd_sc_hd__or2_4 _1165_ (.A(\configy.counter_d[4] ),
    .B(_0523_),
    .X(_0537_));
 sky130_fd_sc_hd__o21a_4 _1166_ (.A1(_0149_),
    .A2(_0537_),
    .B1(_0359_),
    .X(_0538_));
 sky130_fd_sc_hd__o21a_4 _1167_ (.A1(_0531_),
    .A2(_0538_),
    .B1(\configy.counter_d[6] ),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_4 _1168_ (.A(_0399_),
    .B(_0525_),
    .Y(_0540_));
 sky130_fd_sc_hd__or2_4 _1169_ (.A(wbs_data_i[30]),
    .B(_0359_),
    .X(_0541_));
 sky130_fd_sc_hd__and3_4 _1170_ (.A(_0534_),
    .B(_0540_),
    .C(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__or3_4 _1171_ (.A(_0449_),
    .B(_0539_),
    .C(_0542_),
    .X(_0041_));
 sky130_fd_sc_hd__or2_4 _1172_ (.A(wbs_data_i[29]),
    .B(_0360_),
    .X(_0543_));
 sky130_fd_sc_hd__a2bb2o_4 _1173_ (.A1_N(_0531_),
    .A2_N(_0538_),
    .B1(_0537_),
    .B2(_0149_),
    .X(_0544_));
 sky130_fd_sc_hd__buf_2 _1174_ (.A(_0530_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_4 _1175_ (.A(_0149_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__a211o_4 _1176_ (.A1(_0543_),
    .A2(_0544_),
    .B1(_0546_),
    .C1(_0519_),
    .X(_0040_));
 sky130_fd_sc_hd__nand2_4 _1177_ (.A(_0418_),
    .B(_0537_),
    .Y(_0547_));
 sky130_fd_sc_hd__or2_4 _1178_ (.A(wbs_data_i[28]),
    .B(_0398_),
    .X(_0548_));
 sky130_fd_sc_hd__and3_4 _1179_ (.A(_0533_),
    .B(_0547_),
    .C(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__and2_4 _1180_ (.A(_0426_),
    .B(_0523_),
    .X(_0550_));
 sky130_fd_sc_hd__o21a_4 _1181_ (.A1(_0531_),
    .A2(_0550_),
    .B1(\configy.counter_d[4] ),
    .X(_0551_));
 sky130_fd_sc_hd__or3_4 _1182_ (.A(_0449_),
    .B(_0549_),
    .C(_0551_),
    .X(_0039_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(\configy.counter_d[3] ),
    .Y(_0552_));
 sky130_fd_sc_hd__o21ai_4 _1184_ (.A1(_0545_),
    .A2(_0550_),
    .B1(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__or4_4 _1185_ (.A(\configy.counter_d[2] ),
    .B(_0176_),
    .C(\configy.counter_d[0] ),
    .D(_0364_),
    .X(_0554_));
 sky130_fd_sc_hd__o22a_4 _1186_ (.A1(wbs_data_i[27]),
    .A2(_0340_),
    .B1(_0554_),
    .B2(_0552_),
    .X(_0555_));
 sky130_fd_sc_hd__or2_4 _1187_ (.A(_0545_),
    .B(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_4 _1188_ (.A1(_0553_),
    .A2(_0556_),
    .B1(_0324_),
    .X(_0038_));
 sky130_fd_sc_hd__a21bo_4 _1189_ (.A1(wbs_data_i[26]),
    .A2(_0366_),
    .B1_N(_0554_),
    .X(_0557_));
 sky130_fd_sc_hd__o21a_4 _1190_ (.A1(_0176_),
    .A2(_0181_),
    .B1(_0358_),
    .X(_0558_));
 sky130_fd_sc_hd__o21a_4 _1191_ (.A1(_0531_),
    .A2(_0558_),
    .B1(\configy.counter_d[2] ),
    .X(_0559_));
 sky130_fd_sc_hd__a211o_4 _1192_ (.A1(_0534_),
    .A2(_0557_),
    .B1(_0559_),
    .C1(_0519_),
    .X(_0037_));
 sky130_fd_sc_hd__or2_4 _1193_ (.A(wbs_data_i[25]),
    .B(_0414_),
    .X(_0560_));
 sky130_fd_sc_hd__a21bo_4 _1194_ (.A1(_0176_),
    .A2(_0181_),
    .B1_N(_0558_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_4 _1195_ (.A(_0534_),
    .B(_0560_),
    .C(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a211o_4 _1196_ (.A1(_0176_),
    .A2(_0545_),
    .B1(_0562_),
    .C1(_0323_),
    .X(_0036_));
 sky130_fd_sc_hd__or2_4 _1197_ (.A(wbs_data_i[24]),
    .B(_0414_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_4 _1198_ (.A(_0181_),
    .B(_0399_),
    .Y(_0564_));
 sky130_fd_sc_hd__and3_4 _1199_ (.A(_0534_),
    .B(_0563_),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__a211o_4 _1200_ (.A1(_0181_),
    .A2(_0545_),
    .B1(_0565_),
    .C1(_0323_),
    .X(_0035_));
 sky130_fd_sc_hd__o22a_4 _1201_ (.A1(\configy.charged[0] ),
    .A2(_0330_),
    .B1(wbs_sel_i[2]),
    .B2(\configy.charged[2] ),
    .X(_0566_));
 sky130_fd_sc_hd__o22a_4 _1202_ (.A1(\configy.charged[3] ),
    .A2(wbs_sel_i[3]),
    .B1(wbs_sel_i[1]),
    .B2(\configy.charged[1] ),
    .X(_0567_));
 sky130_fd_sc_hd__and3_4 _1203_ (.A(_0342_),
    .B(_0566_),
    .C(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_4 _1204_ (.A(\configy.read_transaction_in_progress ),
    .B(_0326_),
    .Y(_0569_));
 sky130_fd_sc_hd__and4_4 _1205_ (.A(wbs_we_i),
    .B(_0164_),
    .C(_0166_),
    .D(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__buf_2 _1206_ (.A(_0365_),
    .X(_0571_));
 sky130_fd_sc_hd__o21a_4 _1207_ (.A1(_0571_),
    .A2(_0357_),
    .B1(_0333_),
    .X(_0572_));
 sky130_fd_sc_hd__o21a_4 _1208_ (.A1(_0568_),
    .A2(_0570_),
    .B1(_0572_),
    .X(_0034_));
 sky130_fd_sc_hd__buf_2 _1209_ (.A(_0341_),
    .X(_0573_));
 sky130_fd_sc_hd__o21a_4 _1210_ (.A1(_0573_),
    .A2(_0343_),
    .B1(_0572_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_4 _1211_ (.A(_0110_),
    .B(_0328_),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_4 _1212_ (.A(wbs_sel_i[1]),
    .B(_0342_),
    .Y(_0574_));
 sky130_fd_sc_hd__buf_2 _1213_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__and2_4 _1214_ (.A(wbs_data_i[15]),
    .B(_0349_),
    .X(_0576_));
 sky130_fd_sc_hd__a21o_4 _1215_ (.A1(\configy.bits_b[7] ),
    .A2(_0575_),
    .B1(_0576_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_4 _1216_ (.A(wbs_data_i[14]),
    .B(_0349_),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_4 _1217_ (.A1(\configy.bits_b[6] ),
    .A2(_0575_),
    .B1(_0577_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_4 _1218_ (.A(wbs_data_i[13]),
    .B(_0349_),
    .X(_0578_));
 sky130_fd_sc_hd__a21o_4 _1219_ (.A1(\configy.bits_b[5] ),
    .A2(_0575_),
    .B1(_0578_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_4 _1220_ (.A(wbs_data_i[12]),
    .B(_0349_),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_4 _1221_ (.A1(\configy.bits_b[4] ),
    .A2(_0575_),
    .B1(_0579_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_4 _1222_ (.A(wbs_data_i[11]),
    .B(_0348_),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_4 _1223_ (.A1(\configy.bits_b[3] ),
    .A2(_0575_),
    .B1(_0580_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_4 _1224_ (.A(wbs_data_i[10]),
    .B(_0348_),
    .X(_0581_));
 sky130_fd_sc_hd__a21o_4 _1225_ (.A1(\configy.bits_b[2] ),
    .A2(_0574_),
    .B1(_0581_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_4 _1226_ (.A(wbs_data_i[9]),
    .B(_0348_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_4 _1227_ (.A1(\configy.bits_b[1] ),
    .A2(_0574_),
    .B1(_0582_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_4 _1228_ (.A(wbs_data_i[8]),
    .B(_0348_),
    .X(_0583_));
 sky130_fd_sc_hd__a21o_4 _1229_ (.A1(\configy.bits_b[0] ),
    .A2(_0574_),
    .B1(_0583_),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_4 _1230_ (.A(wbs_sel_i[2]),
    .B(_0342_),
    .Y(_0584_));
 sky130_fd_sc_hd__buf_2 _1231_ (.A(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__and2_4 _1232_ (.A(wbs_data_i[23]),
    .B(_0347_),
    .X(_0586_));
 sky130_fd_sc_hd__a21o_4 _1233_ (.A1(\configy.bits_c[7] ),
    .A2(_0585_),
    .B1(_0586_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_4 _1234_ (.A(wbs_data_i[22]),
    .B(_0347_),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_4 _1235_ (.A1(\configy.bits_c[6] ),
    .A2(_0585_),
    .B1(_0587_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_4 _1236_ (.A(wbs_data_i[21]),
    .B(_0347_),
    .X(_0588_));
 sky130_fd_sc_hd__a21o_4 _1237_ (.A1(\configy.bits_c[5] ),
    .A2(_0585_),
    .B1(_0588_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_4 _1238_ (.A(wbs_data_i[20]),
    .B(_0347_),
    .X(_0589_));
 sky130_fd_sc_hd__a21o_4 _1239_ (.A1(\configy.bits_c[4] ),
    .A2(_0585_),
    .B1(_0589_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_4 _1240_ (.A(wbs_data_i[19]),
    .B(_0346_),
    .X(_0590_));
 sky130_fd_sc_hd__a21o_4 _1241_ (.A1(\configy.bits_c[3] ),
    .A2(_0585_),
    .B1(_0590_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_4 _1242_ (.A(wbs_data_i[18]),
    .B(_0346_),
    .X(_0591_));
 sky130_fd_sc_hd__a21o_4 _1243_ (.A1(\configy.bits_c[2] ),
    .A2(_0584_),
    .B1(_0591_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_4 _1244_ (.A(wbs_data_i[17]),
    .B(_0346_),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_4 _1245_ (.A1(\configy.bits_c[1] ),
    .A2(_0584_),
    .B1(_0592_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_4 _1246_ (.A(wbs_data_i[16]),
    .B(_0346_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_4 _1247_ (.A1(\configy.bits_c[0] ),
    .A2(_0584_),
    .B1(_0593_),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_4 _1248_ (.A(wbs_sel_i[3]),
    .B(_0342_),
    .Y(_0594_));
 sky130_fd_sc_hd__buf_2 _1249_ (.A(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__and2_4 _1250_ (.A(wbs_data_i[31]),
    .B(_0338_),
    .X(_0596_));
 sky130_fd_sc_hd__a21o_4 _1251_ (.A1(\configy.bits_d[7] ),
    .A2(_0595_),
    .B1(_0596_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_4 _1252_ (.A(wbs_data_i[30]),
    .B(_0338_),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_4 _1253_ (.A1(\configy.bits_d[6] ),
    .A2(_0595_),
    .B1(_0597_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_4 _1254_ (.A(wbs_data_i[29]),
    .B(_0338_),
    .X(_0598_));
 sky130_fd_sc_hd__a21o_4 _1255_ (.A1(\configy.bits_d[5] ),
    .A2(_0595_),
    .B1(_0598_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_4 _1256_ (.A(wbs_data_i[28]),
    .B(_0338_),
    .X(_0599_));
 sky130_fd_sc_hd__a21o_4 _1257_ (.A1(\configy.bits_d[4] ),
    .A2(_0595_),
    .B1(_0599_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_4 _1258_ (.A(wbs_data_i[27]),
    .B(_0337_),
    .X(_0600_));
 sky130_fd_sc_hd__a21o_4 _1259_ (.A1(\configy.bits_d[3] ),
    .A2(_0595_),
    .B1(_0600_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_4 _1260_ (.A(wbs_data_i[26]),
    .B(_0337_),
    .X(_0601_));
 sky130_fd_sc_hd__a21o_4 _1261_ (.A1(\configy.bits_d[2] ),
    .A2(_0594_),
    .B1(_0601_),
    .X(_0010_));
 sky130_fd_sc_hd__and2_4 _1262_ (.A(wbs_data_i[25]),
    .B(_0337_),
    .X(_0602_));
 sky130_fd_sc_hd__a21o_4 _1263_ (.A1(\configy.bits_d[1] ),
    .A2(_0594_),
    .B1(_0602_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_4 _1264_ (.A(wbs_data_i[24]),
    .B(_0337_),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_4 _1265_ (.A1(\configy.bits_d[0] ),
    .A2(_0594_),
    .B1(_0603_),
    .X(_0008_));
 sky130_fd_sc_hd__nand2_4 _1266_ (.A(_0330_),
    .B(_0336_),
    .Y(_0604_));
 sky130_fd_sc_hd__buf_2 _1267_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__and2_4 _1268_ (.A(wbs_data_i[7]),
    .B(_0351_),
    .X(_0606_));
 sky130_fd_sc_hd__a21o_4 _1269_ (.A1(\configy.bits_a[7] ),
    .A2(_0605_),
    .B1(_0606_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_4 _1270_ (.A(wbs_data_i[6]),
    .B(_0351_),
    .X(_0607_));
 sky130_fd_sc_hd__a21o_4 _1271_ (.A1(\configy.bits_a[6] ),
    .A2(_0605_),
    .B1(_0607_),
    .X(_0006_));
 sky130_fd_sc_hd__and2_4 _1272_ (.A(wbs_data_i[5]),
    .B(_0351_),
    .X(_0608_));
 sky130_fd_sc_hd__a21o_4 _1273_ (.A1(\configy.bits_a[5] ),
    .A2(_0605_),
    .B1(_0608_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_4 _1274_ (.A(wbs_data_i[4]),
    .B(_0351_),
    .X(_0609_));
 sky130_fd_sc_hd__a21o_4 _1275_ (.A1(\configy.bits_a[4] ),
    .A2(_0605_),
    .B1(_0609_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_4 _1276_ (.A(wbs_data_i[3]),
    .B(_0350_),
    .X(_0610_));
 sky130_fd_sc_hd__a21o_4 _1277_ (.A1(\configy.bits_a[3] ),
    .A2(_0605_),
    .B1(_0610_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_4 _1278_ (.A(wbs_data_i[2]),
    .B(_0350_),
    .X(_0611_));
 sky130_fd_sc_hd__a21o_4 _1279_ (.A1(\configy.bits_a[2] ),
    .A2(_0604_),
    .B1(_0611_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_4 _1280_ (.A(wbs_data_i[1]),
    .B(_0350_),
    .X(_0612_));
 sky130_fd_sc_hd__a21o_4 _1281_ (.A1(\configy.bits_a[1] ),
    .A2(_0604_),
    .B1(_0612_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_4 _1282_ (.A(wbs_data_i[0]),
    .B(_0350_),
    .X(_0613_));
 sky130_fd_sc_hd__a21o_4 _1283_ (.A1(\configy.bits_a[0] ),
    .A2(_0604_),
    .B1(_0613_),
    .X(_0000_));
 sky130_fd_sc_hd__nor3_4 _1284_ (.A(\configy.counter_d[7] ),
    .B(_0571_),
    .C(_0525_),
    .Y(set_out[3]));
 sky130_fd_sc_hd__nor3_4 _1285_ (.A(\configy.counter_c[7] ),
    .B(_0571_),
    .C(_0483_),
    .Y(set_out[2]));
 sky130_fd_sc_hd__nor3_4 _1286_ (.A(\configy.counter_b[7] ),
    .B(_0571_),
    .C(_0437_),
    .Y(set_out[1]));
 sky130_fd_sc_hd__nor3_4 _1287_ (.A(\configy.counter_a[7] ),
    .B(_0571_),
    .C(_0382_),
    .Y(set_out[0]));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(\configy.bits_index[2] ),
    .Y(_0614_));
 sky130_fd_sc_hd__buf_2 _1289_ (.A(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__buf_2 _1290_ (.A(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _1291_ (.A(\configy.bits_index[2] ),
    .X(_0617_));
 sky130_fd_sc_hd__or2_4 _1292_ (.A(_0617_),
    .B(\configy.bits_d[2] ),
    .X(_0618_));
 sky130_fd_sc_hd__o21a_4 _1293_ (.A1(_0616_),
    .A2(\configy.bits_d[6] ),
    .B1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__buf_2 _1294_ (.A(_0614_),
    .X(_0620_));
 sky130_fd_sc_hd__or2_4 _1295_ (.A(_0620_),
    .B(\configy.bits_d[7] ),
    .X(_0621_));
 sky130_fd_sc_hd__or2_4 _1296_ (.A(_0352_),
    .B(\configy.bits_d[3] ),
    .X(_0622_));
 sky130_fd_sc_hd__and3_4 _1297_ (.A(_0376_),
    .B(_0621_),
    .C(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__a211o_4 _1298_ (.A1(_0373_),
    .A2(_0619_),
    .B1(_0623_),
    .C1(_0369_),
    .X(_0624_));
 sky130_fd_sc_hd__or2_4 _1299_ (.A(_0617_),
    .B(\configy.bits_d[0] ),
    .X(_0625_));
 sky130_fd_sc_hd__o21a_4 _1300_ (.A1(_0616_),
    .A2(\configy.bits_d[4] ),
    .B1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or2_4 _1301_ (.A(_0620_),
    .B(\configy.bits_d[5] ),
    .X(_0627_));
 sky130_fd_sc_hd__buf_2 _1302_ (.A(\configy.bits_index[2] ),
    .X(_0628_));
 sky130_fd_sc_hd__or2_4 _1303_ (.A(_0628_),
    .B(\configy.bits_d[1] ),
    .X(_0629_));
 sky130_fd_sc_hd__and3_4 _1304_ (.A(_0375_),
    .B(_0627_),
    .C(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__a211o_4 _1305_ (.A1(_0373_),
    .A2(_0626_),
    .B1(_0630_),
    .C1(_0367_),
    .X(_0631_));
 sky130_fd_sc_hd__and3_4 _1306_ (.A(_0573_),
    .B(_0624_),
    .C(_0631_),
    .X(shift_out[3]));
 sky130_fd_sc_hd__or2_4 _1307_ (.A(_0616_),
    .B(\configy.bits_c[5] ),
    .X(_0632_));
 sky130_fd_sc_hd__or2_4 _1308_ (.A(_0353_),
    .B(\configy.bits_c[1] ),
    .X(_0633_));
 sky130_fd_sc_hd__and4_4 _1309_ (.A(_0369_),
    .B(_0376_),
    .C(_0632_),
    .D(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__or2_4 _1310_ (.A(_0353_),
    .B(\configy.bits_c[0] ),
    .X(_0635_));
 sky130_fd_sc_hd__or2_4 _1311_ (.A(_0615_),
    .B(\configy.bits_c[4] ),
    .X(_0636_));
 sky130_fd_sc_hd__or2_4 _1312_ (.A(_0628_),
    .B(\configy.bits_c[2] ),
    .X(_0637_));
 sky130_fd_sc_hd__or2_4 _1313_ (.A(_0614_),
    .B(\configy.bits_c[6] ),
    .X(_0638_));
 sky130_fd_sc_hd__or2_4 _1314_ (.A(_0352_),
    .B(\configy.bits_c[3] ),
    .X(_0639_));
 sky130_fd_sc_hd__o21a_4 _1315_ (.A1(_0615_),
    .A2(\configy.bits_c[7] ),
    .B1(_0375_),
    .X(_0640_));
 sky130_fd_sc_hd__a32o_4 _1316_ (.A1(_0370_),
    .A2(_0637_),
    .A3(_0638_),
    .B1(_0639_),
    .B2(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__a32o_4 _1317_ (.A1(_0371_),
    .A2(_0635_),
    .A3(_0636_),
    .B1(_0641_),
    .B2(_0367_),
    .X(_0642_));
 sky130_fd_sc_hd__o21a_4 _1318_ (.A1(_0634_),
    .A2(_0642_),
    .B1(_0573_),
    .X(shift_out[2]));
 sky130_fd_sc_hd__or2_4 _1319_ (.A(_0617_),
    .B(\configy.bits_b[2] ),
    .X(_0643_));
 sky130_fd_sc_hd__o21a_4 _1320_ (.A1(_0616_),
    .A2(\configy.bits_b[6] ),
    .B1(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__or2_4 _1321_ (.A(_0620_),
    .B(\configy.bits_b[7] ),
    .X(_0645_));
 sky130_fd_sc_hd__or2_4 _1322_ (.A(_0352_),
    .B(\configy.bits_b[3] ),
    .X(_0646_));
 sky130_fd_sc_hd__and3_4 _1323_ (.A(_0376_),
    .B(_0645_),
    .C(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__a211o_4 _1324_ (.A1(_0373_),
    .A2(_0644_),
    .B1(_0647_),
    .C1(_0369_),
    .X(_0648_));
 sky130_fd_sc_hd__or2_4 _1325_ (.A(_0352_),
    .B(\configy.bits_b[0] ),
    .X(_0649_));
 sky130_fd_sc_hd__o21a_4 _1326_ (.A1(_0616_),
    .A2(\configy.bits_b[4] ),
    .B1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__or2_4 _1327_ (.A(_0620_),
    .B(\configy.bits_b[5] ),
    .X(_0651_));
 sky130_fd_sc_hd__or2_4 _1328_ (.A(_0628_),
    .B(\configy.bits_b[1] ),
    .X(_0652_));
 sky130_fd_sc_hd__and3_4 _1329_ (.A(_0375_),
    .B(_0651_),
    .C(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__a211o_4 _1330_ (.A1(_0373_),
    .A2(_0650_),
    .B1(_0653_),
    .C1(_0367_),
    .X(_0654_));
 sky130_fd_sc_hd__and3_4 _1331_ (.A(_0573_),
    .B(_0648_),
    .C(_0654_),
    .X(shift_out[1]));
 sky130_fd_sc_hd__or2_4 _1332_ (.A(_0628_),
    .B(\configy.bits_a[2] ),
    .X(_0655_));
 sky130_fd_sc_hd__or2_4 _1333_ (.A(_0614_),
    .B(\configy.bits_a[6] ),
    .X(_0656_));
 sky130_fd_sc_hd__or2_4 _1334_ (.A(_0628_),
    .B(\configy.bits_a[3] ),
    .X(_0657_));
 sky130_fd_sc_hd__o21a_4 _1335_ (.A1(_0620_),
    .A2(\configy.bits_a[7] ),
    .B1(_0375_),
    .X(_0658_));
 sky130_fd_sc_hd__a32o_4 _1336_ (.A1(_0370_),
    .A2(_0655_),
    .A3(_0656_),
    .B1(_0657_),
    .B2(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__or2_4 _1337_ (.A(_0617_),
    .B(\configy.bits_a[0] ),
    .X(_0660_));
 sky130_fd_sc_hd__or2_4 _1338_ (.A(_0615_),
    .B(\configy.bits_a[4] ),
    .X(_0661_));
 sky130_fd_sc_hd__and3_4 _1339_ (.A(_0371_),
    .B(_0660_),
    .C(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_4 _1340_ (.A(_0615_),
    .B(\configy.bits_a[5] ),
    .X(_0663_));
 sky130_fd_sc_hd__or2_4 _1341_ (.A(_0617_),
    .B(\configy.bits_a[1] ),
    .X(_0664_));
 sky130_fd_sc_hd__and4_4 _1342_ (.A(_0369_),
    .B(_0376_),
    .C(_0663_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__a211o_4 _1343_ (.A1(_0367_),
    .A2(_0659_),
    .B1(_0662_),
    .C1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__and2_4 _1344_ (.A(_0573_),
    .B(_0666_),
    .X(shift_out[0]));
 sky130_fd_sc_hd__or2_4 _1345_ (.A(\configy.free_run ),
    .B(_0341_),
    .X(cen));
 sky130_fd_sc_hd__a21o_4 _1346_ (.A1(_0164_),
    .A2(_0166_),
    .B1(wbs_data_o[31]),
    .X(_0667_));
 sky130_fd_sc_hd__and2_4 _1347_ (.A(\configy.counter_d[7] ),
    .B(_0298_),
    .X(_0668_));
 sky130_fd_sc_hd__and2_4 _1348_ (.A(\configy.bits_d[7] ),
    .B(_0300_),
    .X(_0669_));
 sky130_fd_sc_hd__or4_4 _1349_ (.A(_0173_),
    .B(_0145_),
    .C(_0668_),
    .D(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_4 _1350_ (.A(_0109_),
    .B(_0667_),
    .C(_0670_),
    .X(_0107_));
 sky130_fd_sc_hd__dfxtp_4 _1351_ (.D(_0000_),
    .Q(\configy.bits_a[0] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1352_ (.D(_0001_),
    .Q(\configy.bits_a[1] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1353_ (.D(_0002_),
    .Q(\configy.bits_a[2] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1354_ (.D(_0003_),
    .Q(\configy.bits_a[3] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1355_ (.D(_0004_),
    .Q(\configy.bits_a[4] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1356_ (.D(_0005_),
    .Q(\configy.bits_a[5] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1357_ (.D(_0006_),
    .Q(\configy.bits_a[6] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1358_ (.D(_0007_),
    .Q(\configy.bits_a[7] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1359_ (.D(_0008_),
    .Q(\configy.bits_d[0] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1360_ (.D(_0009_),
    .Q(\configy.bits_d[1] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1361_ (.D(_0010_),
    .Q(\configy.bits_d[2] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1362_ (.D(_0011_),
    .Q(\configy.bits_d[3] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1363_ (.D(_0012_),
    .Q(\configy.bits_d[4] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1364_ (.D(_0013_),
    .Q(\configy.bits_d[5] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1365_ (.D(_0014_),
    .Q(\configy.bits_d[6] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1366_ (.D(_0015_),
    .Q(\configy.bits_d[7] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1367_ (.D(_0016_),
    .Q(\configy.bits_c[0] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1368_ (.D(_0017_),
    .Q(\configy.bits_c[1] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1369_ (.D(_0018_),
    .Q(\configy.bits_c[2] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1370_ (.D(_0019_),
    .Q(\configy.bits_c[3] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1371_ (.D(_0020_),
    .Q(\configy.bits_c[4] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1372_ (.D(_0021_),
    .Q(\configy.bits_c[5] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1373_ (.D(_0022_),
    .Q(\configy.bits_c[6] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1374_ (.D(_0023_),
    .Q(\configy.bits_c[7] ),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1375_ (.D(_0024_),
    .Q(\configy.bits_b[0] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1376_ (.D(_0025_),
    .Q(\configy.bits_b[1] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1377_ (.D(_0026_),
    .Q(\configy.bits_b[2] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1378_ (.D(_0027_),
    .Q(\configy.bits_b[3] ),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1379_ (.D(_0028_),
    .Q(\configy.bits_b[4] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1380_ (.D(_0029_),
    .Q(\configy.bits_b[5] ),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1381_ (.D(_0030_),
    .Q(\configy.bits_b[6] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1382_ (.D(_0031_),
    .Q(\configy.bits_b[7] ),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1383_ (.D(_0032_),
    .Q(wbs_ack_o),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1384_ (.D(_0033_),
    .Q(\configy.output_initiated ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1385_ (.D(_0034_),
    .Q(\configy.write_transaction_in_progress ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1386_ (.D(_0035_),
    .Q(\configy.counter_d[0] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1387_ (.D(_0036_),
    .Q(\configy.counter_d[1] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1388_ (.D(_0037_),
    .Q(\configy.counter_d[2] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1389_ (.D(_0038_),
    .Q(\configy.counter_d[3] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1390_ (.D(_0039_),
    .Q(\configy.counter_d[4] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1391_ (.D(_0040_),
    .Q(\configy.counter_d[5] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1392_ (.D(_0041_),
    .Q(\configy.counter_d[6] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1393_ (.D(_0042_),
    .Q(\configy.counter_d[7] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1394_ (.D(_0043_),
    .Q(\configy.counter_c[0] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1395_ (.D(_0044_),
    .Q(\configy.counter_c[1] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1396_ (.D(_0045_),
    .Q(\configy.counter_c[2] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1397_ (.D(_0046_),
    .Q(\configy.counter_c[3] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1398_ (.D(_0047_),
    .Q(\configy.counter_c[4] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1399_ (.D(_0048_),
    .Q(\configy.counter_c[5] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1400_ (.D(_0049_),
    .Q(\configy.counter_c[6] ),
    .CLK(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1401_ (.D(_0050_),
    .Q(\configy.counter_c[7] ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1402_ (.D(_0051_),
    .Q(\configy.counter_b[0] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1403_ (.D(_0052_),
    .Q(\configy.counter_b[1] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1404_ (.D(_0053_),
    .Q(\configy.counter_b[2] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1405_ (.D(_0054_),
    .Q(\configy.counter_b[3] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1406_ (.D(_0055_),
    .Q(\configy.counter_b[4] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1407_ (.D(_0056_),
    .Q(\configy.counter_b[5] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1408_ (.D(_0057_),
    .Q(\configy.counter_b[6] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1409_ (.D(_0058_),
    .Q(\configy.counter_b[7] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1410_ (.D(_0059_),
    .Q(\configy.counter_a[0] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1411_ (.D(_0060_),
    .Q(\configy.counter_a[1] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1412_ (.D(_0061_),
    .Q(\configy.counter_a[2] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1413_ (.D(_0062_),
    .Q(\configy.counter_a[3] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1414_ (.D(_0063_),
    .Q(\configy.counter_a[4] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1415_ (.D(_0064_),
    .Q(\configy.counter_a[5] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1416_ (.D(_0065_),
    .Q(\configy.counter_a[6] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1417_ (.D(_0066_),
    .Q(\configy.counter_a[7] ),
    .CLK(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1418_ (.D(_0067_),
    .Q(\configy.bits_index[0] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1419_ (.D(_0068_),
    .Q(\configy.bits_index[1] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1420_ (.D(_0069_),
    .Q(\configy.bits_index[2] ),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1421_ (.D(_0070_),
    .Q(\configy.charged[0] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1422_ (.D(_0071_),
    .Q(\configy.charged[1] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1423_ (.D(_0072_),
    .Q(\configy.charged[2] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1424_ (.D(_0073_),
    .Q(\configy.charged[3] ),
    .CLK(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1425_ (.D(_0074_),
    .Q(\configy.free_run ),
    .CLK(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1426_ (.D(_0075_),
    .Q(\configy.read_transaction_in_progress ),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1427_ (.D(_0076_),
    .Q(wbs_data_o[0]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1428_ (.D(_0077_),
    .Q(wbs_data_o[1]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1429_ (.D(_0078_),
    .Q(wbs_data_o[2]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1430_ (.D(_0079_),
    .Q(wbs_data_o[3]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1431_ (.D(_0080_),
    .Q(wbs_data_o[4]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1432_ (.D(_0081_),
    .Q(wbs_data_o[5]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1433_ (.D(_0082_),
    .Q(wbs_data_o[6]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1434_ (.D(_0083_),
    .Q(wbs_data_o[7]),
    .CLK(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1435_ (.D(_0084_),
    .Q(wbs_data_o[8]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1436_ (.D(_0085_),
    .Q(wbs_data_o[9]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1437_ (.D(_0086_),
    .Q(wbs_data_o[10]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1438_ (.D(_0087_),
    .Q(wbs_data_o[11]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1439_ (.D(_0088_),
    .Q(wbs_data_o[12]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1440_ (.D(_0089_),
    .Q(wbs_data_o[13]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1441_ (.D(_0090_),
    .Q(wbs_data_o[14]),
    .CLK(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1442_ (.D(_0091_),
    .Q(wbs_data_o[15]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1443_ (.D(_0092_),
    .Q(wbs_data_o[16]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1444_ (.D(_0093_),
    .Q(wbs_data_o[17]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1445_ (.D(_0094_),
    .Q(wbs_data_o[18]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1446_ (.D(_0095_),
    .Q(wbs_data_o[19]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1447_ (.D(_0096_),
    .Q(wbs_data_o[20]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1448_ (.D(_0097_),
    .Q(wbs_data_o[21]),
    .CLK(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1449_ (.D(_0098_),
    .Q(wbs_data_o[22]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1450_ (.D(_0099_),
    .Q(wbs_data_o[23]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1451_ (.D(_0100_),
    .Q(wbs_data_o[24]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1452_ (.D(_0101_),
    .Q(wbs_data_o[25]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1453_ (.D(_0102_),
    .Q(wbs_data_o[26]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1454_ (.D(_0103_),
    .Q(wbs_data_o[27]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1455_ (.D(_0104_),
    .Q(wbs_data_o[28]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1456_ (.D(_0105_),
    .Q(wbs_data_o[29]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1457_ (.D(_0106_),
    .Q(wbs_data_o[30]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__dfxtp_4 _1458_ (.D(_0107_),
    .Q(wbs_data_o[31]),
    .CLK(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_0 (.DIODE(wbs_data_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(wbs_data_i[29]));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_590 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_276 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_313 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_480 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_602 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_367 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_594 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_437 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_522 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_574 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_646 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_267 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_298 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_92 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_396 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_514 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_580 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_628 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_646 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_484 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_532 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_213 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_325 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_519 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_556 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_467 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_548 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_606 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_566 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_628 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_406 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_467 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_579 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_605 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_639 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_651 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_663 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_358 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_388 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_463 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_476 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_646 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_222 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_311 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_366 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_398 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_640 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_22 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_396 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_619 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_641 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_100 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_459 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_157 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_522 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_562 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_602 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_630 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_280 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_471 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_673 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_76 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_400 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_436 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_550 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_624 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_644 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_227 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_368 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_423 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_487 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_518 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_527 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_596 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_633 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_649 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_574 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_644 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_48 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_549 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_638 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_312 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_554 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_578 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_608 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_647 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_170 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_552 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_600 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_639 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_241 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_266 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_382 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_463 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_518 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_554 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_602 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_630 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_243 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_406 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_450 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_459 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_572 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_593 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_637 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_254 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_297 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_364 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_367 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_440 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_462 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_521 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_586 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_598 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_611 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_623 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_635 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_647 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_672 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_304 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_356 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_456 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_459 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_471 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_511 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_578 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_581 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_593 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_605 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_629 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_674 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_240 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_302 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_462 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_466 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_524 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_588 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_590 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_621 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_645 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_672 ();
endmodule
