VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_tile
  CLASS BLOCK ;
  FOREIGN mac_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 2198.860 BY 2286.000 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.330 44.120 2122.610 48.120 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2132.910 44.120 2133.190 48.120 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2237.840 2149.480 2238.440 ;
    END
  END cset
  PIN cset_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2143.490 44.120 2143.770 48.120 ;
    END
  END cset_out
  PIN east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 49.600 2149.480 50.200 ;
    END
  END east[0]
  PIN east[100]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1177.040 2149.480 1177.640 ;
    END
  END east[100]
  PIN east[101]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1188.600 2149.480 1189.200 ;
    END
  END east[101]
  PIN east[102]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1200.160 2149.480 1200.760 ;
    END
  END east[102]
  PIN east[103]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1211.040 2149.480 1211.640 ;
    END
  END east[103]
  PIN east[104]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1222.600 2149.480 1223.200 ;
    END
  END east[104]
  PIN east[105]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1233.480 2149.480 1234.080 ;
    END
  END east[105]
  PIN east[106]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1245.040 2149.480 1245.640 ;
    END
  END east[106]
  PIN east[107]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1256.600 2149.480 1257.200 ;
    END
  END east[107]
  PIN east[108]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1267.480 2149.480 1268.080 ;
    END
  END east[108]
  PIN east[109]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1279.040 2149.480 1279.640 ;
    END
  END east[109]
  PIN east[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 161.800 2149.480 162.400 ;
    END
  END east[10]
  PIN east[110]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1289.920 2149.480 1290.520 ;
    END
  END east[110]
  PIN east[111]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1301.480 2149.480 1302.080 ;
    END
  END east[111]
  PIN east[112]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1313.040 2149.480 1313.640 ;
    END
  END east[112]
  PIN east[113]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1323.920 2149.480 1324.520 ;
    END
  END east[113]
  PIN east[114]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1335.480 2149.480 1336.080 ;
    END
  END east[114]
  PIN east[115]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1346.360 2149.480 1346.960 ;
    END
  END east[115]
  PIN east[116]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1357.920 2149.480 1358.520 ;
    END
  END east[116]
  PIN east[117]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1369.480 2149.480 1370.080 ;
    END
  END east[117]
  PIN east[118]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1380.360 2149.480 1380.960 ;
    END
  END east[118]
  PIN east[119]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1391.920 2149.480 1392.520 ;
    END
  END east[119]
  PIN east[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 173.360 2149.480 173.960 ;
    END
  END east[11]
  PIN east[120]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1402.800 2149.480 1403.400 ;
    END
  END east[120]
  PIN east[121]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1414.360 2149.480 1414.960 ;
    END
  END east[121]
  PIN east[122]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1425.240 2149.480 1425.840 ;
    END
  END east[122]
  PIN east[123]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1436.800 2149.480 1437.400 ;
    END
  END east[123]
  PIN east[124]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1448.360 2149.480 1448.960 ;
    END
  END east[124]
  PIN east[125]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1459.240 2149.480 1459.840 ;
    END
  END east[125]
  PIN east[126]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1470.800 2149.480 1471.400 ;
    END
  END east[126]
  PIN east[127]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1481.680 2149.480 1482.280 ;
    END
  END east[127]
  PIN east[128]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1493.240 2149.480 1493.840 ;
    END
  END east[128]
  PIN east[129]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1504.800 2149.480 1505.400 ;
    END
  END east[129]
  PIN east[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 184.920 2149.480 185.520 ;
    END
  END east[12]
  PIN east[130]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1515.680 2149.480 1516.280 ;
    END
  END east[130]
  PIN east[131]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1527.240 2149.480 1527.840 ;
    END
  END east[131]
  PIN east[132]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1538.120 2149.480 1538.720 ;
    END
  END east[132]
  PIN east[133]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1549.680 2149.480 1550.280 ;
    END
  END east[133]
  PIN east[134]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1561.240 2149.480 1561.840 ;
    END
  END east[134]
  PIN east[135]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1572.120 2149.480 1572.720 ;
    END
  END east[135]
  PIN east[136]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1583.680 2149.480 1584.280 ;
    END
  END east[136]
  PIN east[137]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1594.560 2149.480 1595.160 ;
    END
  END east[137]
  PIN east[138]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1606.120 2149.480 1606.720 ;
    END
  END east[138]
  PIN east[139]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1617.000 2149.480 1617.600 ;
    END
  END east[139]
  PIN east[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 195.800 2149.480 196.400 ;
    END
  END east[13]
  PIN east[140]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1628.560 2149.480 1629.160 ;
    END
  END east[140]
  PIN east[141]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1640.120 2149.480 1640.720 ;
    END
  END east[141]
  PIN east[142]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1651.000 2149.480 1651.600 ;
    END
  END east[142]
  PIN east[143]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1662.560 2149.480 1663.160 ;
    END
  END east[143]
  PIN east[144]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1673.440 2149.480 1674.040 ;
    END
  END east[144]
  PIN east[145]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1685.000 2149.480 1685.600 ;
    END
  END east[145]
  PIN east[146]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1696.560 2149.480 1697.160 ;
    END
  END east[146]
  PIN east[147]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1707.440 2149.480 1708.040 ;
    END
  END east[147]
  PIN east[148]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1719.000 2149.480 1719.600 ;
    END
  END east[148]
  PIN east[149]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1729.880 2149.480 1730.480 ;
    END
  END east[149]
  PIN east[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 207.360 2149.480 207.960 ;
    END
  END east[14]
  PIN east[150]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1741.440 2149.480 1742.040 ;
    END
  END east[150]
  PIN east[151]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1753.000 2149.480 1753.600 ;
    END
  END east[151]
  PIN east[152]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1763.880 2149.480 1764.480 ;
    END
  END east[152]
  PIN east[153]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1775.440 2149.480 1776.040 ;
    END
  END east[153]
  PIN east[154]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1786.320 2149.480 1786.920 ;
    END
  END east[154]
  PIN east[155]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1797.880 2149.480 1798.480 ;
    END
  END east[155]
  PIN east[156]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1809.440 2149.480 1810.040 ;
    END
  END east[156]
  PIN east[157]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1820.320 2149.480 1820.920 ;
    END
  END east[157]
  PIN east[158]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1831.880 2149.480 1832.480 ;
    END
  END east[158]
  PIN east[159]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1842.760 2149.480 1843.360 ;
    END
  END east[159]
  PIN east[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 218.240 2149.480 218.840 ;
    END
  END east[15]
  PIN east[160]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1854.320 2149.480 1854.920 ;
    END
  END east[160]
  PIN east[161]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1865.200 2149.480 1865.800 ;
    END
  END east[161]
  PIN east[162]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1876.760 2149.480 1877.360 ;
    END
  END east[162]
  PIN east[163]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1888.320 2149.480 1888.920 ;
    END
  END east[163]
  PIN east[164]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1899.200 2149.480 1899.800 ;
    END
  END east[164]
  PIN east[165]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1910.760 2149.480 1911.360 ;
    END
  END east[165]
  PIN east[166]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1921.640 2149.480 1922.240 ;
    END
  END east[166]
  PIN east[167]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1933.200 2149.480 1933.800 ;
    END
  END east[167]
  PIN east[168]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1944.760 2149.480 1945.360 ;
    END
  END east[168]
  PIN east[169]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1955.640 2149.480 1956.240 ;
    END
  END east[169]
  PIN east[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 229.800 2149.480 230.400 ;
    END
  END east[16]
  PIN east[170]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1967.200 2149.480 1967.800 ;
    END
  END east[170]
  PIN east[171]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1978.080 2149.480 1978.680 ;
    END
  END east[171]
  PIN east[172]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1989.640 2149.480 1990.240 ;
    END
  END east[172]
  PIN east[173]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2001.200 2149.480 2001.800 ;
    END
  END east[173]
  PIN east[174]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2012.080 2149.480 2012.680 ;
    END
  END east[174]
  PIN east[175]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2023.640 2149.480 2024.240 ;
    END
  END east[175]
  PIN east[176]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2034.520 2149.480 2035.120 ;
    END
  END east[176]
  PIN east[177]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2046.080 2149.480 2046.680 ;
    END
  END east[177]
  PIN east[178]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2056.960 2149.480 2057.560 ;
    END
  END east[178]
  PIN east[179]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2068.520 2149.480 2069.120 ;
    END
  END east[179]
  PIN east[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 241.360 2149.480 241.960 ;
    END
  END east[17]
  PIN east[180]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2080.080 2149.480 2080.680 ;
    END
  END east[180]
  PIN east[181]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2090.960 2149.480 2091.560 ;
    END
  END east[181]
  PIN east[182]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2102.520 2149.480 2103.120 ;
    END
  END east[182]
  PIN east[183]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2113.400 2149.480 2114.000 ;
    END
  END east[183]
  PIN east[184]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2124.960 2149.480 2125.560 ;
    END
  END east[184]
  PIN east[185]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2136.520 2149.480 2137.120 ;
    END
  END east[185]
  PIN east[186]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2147.400 2149.480 2148.000 ;
    END
  END east[186]
  PIN east[187]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2158.960 2149.480 2159.560 ;
    END
  END east[187]
  PIN east[188]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2169.840 2149.480 2170.440 ;
    END
  END east[188]
  PIN east[189]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2181.400 2149.480 2182.000 ;
    END
  END east[189]
  PIN east[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 252.240 2149.480 252.840 ;
    END
  END east[18]
  PIN east[190]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2192.960 2149.480 2193.560 ;
    END
  END east[190]
  PIN east[191]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2203.840 2149.480 2204.440 ;
    END
  END east[191]
  PIN east[192]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2215.400 2149.480 2216.000 ;
    END
  END east[192]
  PIN east[193]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 2226.280 2149.480 2226.880 ;
    END
  END east[193]
  PIN east[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 263.800 2149.480 264.400 ;
    END
  END east[19]
  PIN east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 60.480 2149.480 61.080 ;
    END
  END east[1]
  PIN east[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 274.680 2149.480 275.280 ;
    END
  END east[20]
  PIN east[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 286.240 2149.480 286.840 ;
    END
  END east[21]
  PIN east[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 297.120 2149.480 297.720 ;
    END
  END east[22]
  PIN east[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 308.680 2149.480 309.280 ;
    END
  END east[23]
  PIN east[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 320.240 2149.480 320.840 ;
    END
  END east[24]
  PIN east[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 331.120 2149.480 331.720 ;
    END
  END east[25]
  PIN east[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 342.680 2149.480 343.280 ;
    END
  END east[26]
  PIN east[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 353.560 2149.480 354.160 ;
    END
  END east[27]
  PIN east[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 365.120 2149.480 365.720 ;
    END
  END east[28]
  PIN east[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 376.680 2149.480 377.280 ;
    END
  END east[29]
  PIN east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 72.040 2149.480 72.640 ;
    END
  END east[2]
  PIN east[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 387.560 2149.480 388.160 ;
    END
  END east[30]
  PIN east[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 399.120 2149.480 399.720 ;
    END
  END east[31]
  PIN east[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 410.000 2149.480 410.600 ;
    END
  END east[32]
  PIN east[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 421.560 2149.480 422.160 ;
    END
  END east[33]
  PIN east[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 433.120 2149.480 433.720 ;
    END
  END east[34]
  PIN east[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 444.000 2149.480 444.600 ;
    END
  END east[35]
  PIN east[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 455.560 2149.480 456.160 ;
    END
  END east[36]
  PIN east[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 466.440 2149.480 467.040 ;
    END
  END east[37]
  PIN east[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 478.000 2149.480 478.600 ;
    END
  END east[38]
  PIN east[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 489.560 2149.480 490.160 ;
    END
  END east[39]
  PIN east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 82.920 2149.480 83.520 ;
    END
  END east[3]
  PIN east[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 500.440 2149.480 501.040 ;
    END
  END east[40]
  PIN east[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 512.000 2149.480 512.600 ;
    END
  END east[41]
  PIN east[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 522.880 2149.480 523.480 ;
    END
  END east[42]
  PIN east[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 534.440 2149.480 535.040 ;
    END
  END east[43]
  PIN east[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 545.320 2149.480 545.920 ;
    END
  END east[44]
  PIN east[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 556.880 2149.480 557.480 ;
    END
  END east[45]
  PIN east[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 568.440 2149.480 569.040 ;
    END
  END east[46]
  PIN east[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 579.320 2149.480 579.920 ;
    END
  END east[47]
  PIN east[48]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 590.880 2149.480 591.480 ;
    END
  END east[48]
  PIN east[49]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 601.760 2149.480 602.360 ;
    END
  END east[49]
  PIN east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 94.480 2149.480 95.080 ;
    END
  END east[4]
  PIN east[50]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 613.320 2149.480 613.920 ;
    END
  END east[50]
  PIN east[51]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 624.880 2149.480 625.480 ;
    END
  END east[51]
  PIN east[52]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 635.760 2149.480 636.360 ;
    END
  END east[52]
  PIN east[53]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 647.320 2149.480 647.920 ;
    END
  END east[53]
  PIN east[54]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 658.200 2149.480 658.800 ;
    END
  END east[54]
  PIN east[55]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 669.760 2149.480 670.360 ;
    END
  END east[55]
  PIN east[56]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 681.320 2149.480 681.920 ;
    END
  END east[56]
  PIN east[57]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 692.200 2149.480 692.800 ;
    END
  END east[57]
  PIN east[58]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 703.760 2149.480 704.360 ;
    END
  END east[58]
  PIN east[59]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 714.640 2149.480 715.240 ;
    END
  END east[59]
  PIN east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 105.360 2149.480 105.960 ;
    END
  END east[5]
  PIN east[60]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 726.200 2149.480 726.800 ;
    END
  END east[60]
  PIN east[61]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 737.080 2149.480 737.680 ;
    END
  END east[61]
  PIN east[62]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 748.640 2149.480 749.240 ;
    END
  END east[62]
  PIN east[63]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 760.200 2149.480 760.800 ;
    END
  END east[63]
  PIN east[64]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 771.080 2149.480 771.680 ;
    END
  END east[64]
  PIN east[65]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 782.640 2149.480 783.240 ;
    END
  END east[65]
  PIN east[66]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 793.520 2149.480 794.120 ;
    END
  END east[66]
  PIN east[67]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 805.080 2149.480 805.680 ;
    END
  END east[67]
  PIN east[68]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 816.640 2149.480 817.240 ;
    END
  END east[68]
  PIN east[69]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 827.520 2149.480 828.120 ;
    END
  END east[69]
  PIN east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 116.920 2149.480 117.520 ;
    END
  END east[6]
  PIN east[70]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 839.080 2149.480 839.680 ;
    END
  END east[70]
  PIN east[71]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 849.960 2149.480 850.560 ;
    END
  END east[71]
  PIN east[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 861.520 2149.480 862.120 ;
    END
  END east[72]
  PIN east[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 873.080 2149.480 873.680 ;
    END
  END east[73]
  PIN east[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 883.960 2149.480 884.560 ;
    END
  END east[74]
  PIN east[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 895.520 2149.480 896.120 ;
    END
  END east[75]
  PIN east[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 906.400 2149.480 907.000 ;
    END
  END east[76]
  PIN east[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 917.960 2149.480 918.560 ;
    END
  END east[77]
  PIN east[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 929.520 2149.480 930.120 ;
    END
  END east[78]
  PIN east[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 940.400 2149.480 941.000 ;
    END
  END east[79]
  PIN east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 128.480 2149.480 129.080 ;
    END
  END east[7]
  PIN east[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 951.960 2149.480 952.560 ;
    END
  END east[80]
  PIN east[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 962.840 2149.480 963.440 ;
    END
  END east[81]
  PIN east[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 974.400 2149.480 975.000 ;
    END
  END east[82]
  PIN east[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 985.280 2149.480 985.880 ;
    END
  END east[83]
  PIN east[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 996.840 2149.480 997.440 ;
    END
  END east[84]
  PIN east[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1008.400 2149.480 1009.000 ;
    END
  END east[85]
  PIN east[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1019.280 2149.480 1019.880 ;
    END
  END east[86]
  PIN east[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1030.840 2149.480 1031.440 ;
    END
  END east[87]
  PIN east[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1041.720 2149.480 1042.320 ;
    END
  END east[88]
  PIN east[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1053.280 2149.480 1053.880 ;
    END
  END east[89]
  PIN east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 139.360 2149.480 139.960 ;
    END
  END east[8]
  PIN east[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1064.840 2149.480 1065.440 ;
    END
  END east[90]
  PIN east[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1075.720 2149.480 1076.320 ;
    END
  END east[91]
  PIN east[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1087.280 2149.480 1087.880 ;
    END
  END east[92]
  PIN east[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1098.160 2149.480 1098.760 ;
    END
  END east[93]
  PIN east[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1109.720 2149.480 1110.320 ;
    END
  END east[94]
  PIN east[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1121.280 2149.480 1121.880 ;
    END
  END east[95]
  PIN east[96]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1132.160 2149.480 1132.760 ;
    END
  END east[96]
  PIN east[97]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1143.720 2149.480 1144.320 ;
    END
  END east[97]
  PIN east[98]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1154.600 2149.480 1155.200 ;
    END
  END east[98]
  PIN east[99]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 1166.160 2149.480 1166.760 ;
    END
  END east[99]
  PIN east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2145.480 150.920 2149.480 151.520 ;
    END
  END east[9]
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2226.280 53.480 2226.880 ;
    END
  END en
  PIN north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.630 2240.120 54.910 2244.120 ;
    END
  END north[0]
  PIN north[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1131.490 2240.120 1131.770 2244.120 ;
    END
  END north[100]
  PIN north[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1142.070 2240.120 1142.350 2244.120 ;
    END
  END north[101]
  PIN north[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1152.650 2240.120 1152.930 2244.120 ;
    END
  END north[102]
  PIN north[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1163.690 2240.120 1163.970 2244.120 ;
    END
  END north[103]
  PIN north[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1174.270 2240.120 1174.550 2244.120 ;
    END
  END north[104]
  PIN north[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1185.310 2240.120 1185.590 2244.120 ;
    END
  END north[105]
  PIN north[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1195.890 2240.120 1196.170 2244.120 ;
    END
  END north[106]
  PIN north[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1206.470 2240.120 1206.750 2244.120 ;
    END
  END north[107]
  PIN north[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1217.510 2240.120 1217.790 2244.120 ;
    END
  END north[108]
  PIN north[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1228.090 2240.120 1228.370 2244.120 ;
    END
  END north[109]
  PIN north[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 162.270 2240.120 162.550 2244.120 ;
    END
  END north[10]
  PIN north[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1239.130 2240.120 1239.410 2244.120 ;
    END
  END north[110]
  PIN north[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1249.710 2240.120 1249.990 2244.120 ;
    END
  END north[111]
  PIN north[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1260.290 2240.120 1260.570 2244.120 ;
    END
  END north[112]
  PIN north[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1271.330 2240.120 1271.610 2244.120 ;
    END
  END north[113]
  PIN north[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1281.910 2240.120 1282.190 2244.120 ;
    END
  END north[114]
  PIN north[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1292.950 2240.120 1293.230 2244.120 ;
    END
  END north[115]
  PIN north[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1303.530 2240.120 1303.810 2244.120 ;
    END
  END north[116]
  PIN north[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1314.570 2240.120 1314.850 2244.120 ;
    END
  END north[117]
  PIN north[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1325.150 2240.120 1325.430 2244.120 ;
    END
  END north[118]
  PIN north[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1335.730 2240.120 1336.010 2244.120 ;
    END
  END north[119]
  PIN north[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 172.850 2240.120 173.130 2244.120 ;
    END
  END north[11]
  PIN north[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1346.770 2240.120 1347.050 2244.120 ;
    END
  END north[120]
  PIN north[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1357.350 2240.120 1357.630 2244.120 ;
    END
  END north[121]
  PIN north[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1368.390 2240.120 1368.670 2244.120 ;
    END
  END north[122]
  PIN north[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1378.970 2240.120 1379.250 2244.120 ;
    END
  END north[123]
  PIN north[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1389.550 2240.120 1389.830 2244.120 ;
    END
  END north[124]
  PIN north[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1400.590 2240.120 1400.870 2244.120 ;
    END
  END north[125]
  PIN north[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1411.170 2240.120 1411.450 2244.120 ;
    END
  END north[126]
  PIN north[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1422.210 2240.120 1422.490 2244.120 ;
    END
  END north[127]
  PIN north[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1432.790 2240.120 1433.070 2244.120 ;
    END
  END north[128]
  PIN north[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1443.370 2240.120 1443.650 2244.120 ;
    END
  END north[129]
  PIN north[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 183.430 2240.120 183.710 2244.120 ;
    END
  END north[12]
  PIN north[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1454.410 2240.120 1454.690 2244.120 ;
    END
  END north[130]
  PIN north[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1464.990 2240.120 1465.270 2244.120 ;
    END
  END north[131]
  PIN north[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1476.030 2240.120 1476.310 2244.120 ;
    END
  END north[132]
  PIN north[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1486.610 2240.120 1486.890 2244.120 ;
    END
  END north[133]
  PIN north[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1497.190 2240.120 1497.470 2244.120 ;
    END
  END north[134]
  PIN north[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1508.230 2240.120 1508.510 2244.120 ;
    END
  END north[135]
  PIN north[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1518.810 2240.120 1519.090 2244.120 ;
    END
  END north[136]
  PIN north[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1529.850 2240.120 1530.130 2244.120 ;
    END
  END north[137]
  PIN north[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1540.430 2240.120 1540.710 2244.120 ;
    END
  END north[138]
  PIN north[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1551.470 2240.120 1551.750 2244.120 ;
    END
  END north[139]
  PIN north[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 194.470 2240.120 194.750 2244.120 ;
    END
  END north[13]
  PIN north[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1562.050 2240.120 1562.330 2244.120 ;
    END
  END north[140]
  PIN north[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1572.630 2240.120 1572.910 2244.120 ;
    END
  END north[141]
  PIN north[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1583.670 2240.120 1583.950 2244.120 ;
    END
  END north[142]
  PIN north[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1594.250 2240.120 1594.530 2244.120 ;
    END
  END north[143]
  PIN north[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1605.290 2240.120 1605.570 2244.120 ;
    END
  END north[144]
  PIN north[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1615.870 2240.120 1616.150 2244.120 ;
    END
  END north[145]
  PIN north[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1626.450 2240.120 1626.730 2244.120 ;
    END
  END north[146]
  PIN north[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1637.490 2240.120 1637.770 2244.120 ;
    END
  END north[147]
  PIN north[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1648.070 2240.120 1648.350 2244.120 ;
    END
  END north[148]
  PIN north[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1659.110 2240.120 1659.390 2244.120 ;
    END
  END north[149]
  PIN north[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 205.050 2240.120 205.330 2244.120 ;
    END
  END north[14]
  PIN north[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1669.690 2240.120 1669.970 2244.120 ;
    END
  END north[150]
  PIN north[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1680.270 2240.120 1680.550 2244.120 ;
    END
  END north[151]
  PIN north[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1691.310 2240.120 1691.590 2244.120 ;
    END
  END north[152]
  PIN north[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1701.890 2240.120 1702.170 2244.120 ;
    END
  END north[153]
  PIN north[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1712.930 2240.120 1713.210 2244.120 ;
    END
  END north[154]
  PIN north[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1723.510 2240.120 1723.790 2244.120 ;
    END
  END north[155]
  PIN north[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1734.550 2240.120 1734.830 2244.120 ;
    END
  END north[156]
  PIN north[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1745.130 2240.120 1745.410 2244.120 ;
    END
  END north[157]
  PIN north[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1755.710 2240.120 1755.990 2244.120 ;
    END
  END north[158]
  PIN north[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1766.750 2240.120 1767.030 2244.120 ;
    END
  END north[159]
  PIN north[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 216.090 2240.120 216.370 2244.120 ;
    END
  END north[15]
  PIN north[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1777.330 2240.120 1777.610 2244.120 ;
    END
  END north[160]
  PIN north[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1788.370 2240.120 1788.650 2244.120 ;
    END
  END north[161]
  PIN north[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1798.950 2240.120 1799.230 2244.120 ;
    END
  END north[162]
  PIN north[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1809.530 2240.120 1809.810 2244.120 ;
    END
  END north[163]
  PIN north[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1820.570 2240.120 1820.850 2244.120 ;
    END
  END north[164]
  PIN north[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1831.150 2240.120 1831.430 2244.120 ;
    END
  END north[165]
  PIN north[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1842.190 2240.120 1842.470 2244.120 ;
    END
  END north[166]
  PIN north[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1852.770 2240.120 1853.050 2244.120 ;
    END
  END north[167]
  PIN north[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1863.350 2240.120 1863.630 2244.120 ;
    END
  END north[168]
  PIN north[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1874.390 2240.120 1874.670 2244.120 ;
    END
  END north[169]
  PIN north[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 226.670 2240.120 226.950 2244.120 ;
    END
  END north[16]
  PIN north[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1884.970 2240.120 1885.250 2244.120 ;
    END
  END north[170]
  PIN north[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1896.010 2240.120 1896.290 2244.120 ;
    END
  END north[171]
  PIN north[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1906.590 2240.120 1906.870 2244.120 ;
    END
  END north[172]
  PIN north[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1917.170 2240.120 1917.450 2244.120 ;
    END
  END north[173]
  PIN north[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1928.210 2240.120 1928.490 2244.120 ;
    END
  END north[174]
  PIN north[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1938.790 2240.120 1939.070 2244.120 ;
    END
  END north[175]
  PIN north[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1949.830 2240.120 1950.110 2244.120 ;
    END
  END north[176]
  PIN north[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1960.410 2240.120 1960.690 2244.120 ;
    END
  END north[177]
  PIN north[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1971.450 2240.120 1971.730 2244.120 ;
    END
  END north[178]
  PIN north[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1982.030 2240.120 1982.310 2244.120 ;
    END
  END north[179]
  PIN north[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 237.250 2240.120 237.530 2244.120 ;
    END
  END north[17]
  PIN north[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1992.610 2240.120 1992.890 2244.120 ;
    END
  END north[180]
  PIN north[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2003.650 2240.120 2003.930 2244.120 ;
    END
  END north[181]
  PIN north[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2014.230 2240.120 2014.510 2244.120 ;
    END
  END north[182]
  PIN north[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2025.270 2240.120 2025.550 2244.120 ;
    END
  END north[183]
  PIN north[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2035.850 2240.120 2036.130 2244.120 ;
    END
  END north[184]
  PIN north[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2046.430 2240.120 2046.710 2244.120 ;
    END
  END north[185]
  PIN north[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2057.470 2240.120 2057.750 2244.120 ;
    END
  END north[186]
  PIN north[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2068.050 2240.120 2068.330 2244.120 ;
    END
  END north[187]
  PIN north[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2079.090 2240.120 2079.370 2244.120 ;
    END
  END north[188]
  PIN north[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2089.670 2240.120 2089.950 2244.120 ;
    END
  END north[189]
  PIN north[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 248.290 2240.120 248.570 2244.120 ;
    END
  END north[18]
  PIN north[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2100.250 2240.120 2100.530 2244.120 ;
    END
  END north[190]
  PIN north[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2111.290 2240.120 2111.570 2244.120 ;
    END
  END north[191]
  PIN north[192]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2121.870 2240.120 2122.150 2244.120 ;
    END
  END north[192]
  PIN north[193]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2132.910 2240.120 2133.190 2244.120 ;
    END
  END north[193]
  PIN north[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 258.870 2240.120 259.150 2244.120 ;
    END
  END north[19]
  PIN north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 65.210 2240.120 65.490 2244.120 ;
    END
  END north[1]
  PIN north[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 269.910 2240.120 270.190 2244.120 ;
    END
  END north[20]
  PIN north[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 280.490 2240.120 280.770 2244.120 ;
    END
  END north[21]
  PIN north[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 291.530 2240.120 291.810 2244.120 ;
    END
  END north[22]
  PIN north[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 302.110 2240.120 302.390 2244.120 ;
    END
  END north[23]
  PIN north[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 312.690 2240.120 312.970 2244.120 ;
    END
  END north[24]
  PIN north[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 323.730 2240.120 324.010 2244.120 ;
    END
  END north[25]
  PIN north[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 334.310 2240.120 334.590 2244.120 ;
    END
  END north[26]
  PIN north[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 345.350 2240.120 345.630 2244.120 ;
    END
  END north[27]
  PIN north[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 355.930 2240.120 356.210 2244.120 ;
    END
  END north[28]
  PIN north[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 366.510 2240.120 366.790 2244.120 ;
    END
  END north[29]
  PIN north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.790 2240.120 76.070 2244.120 ;
    END
  END north[2]
  PIN north[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 377.550 2240.120 377.830 2244.120 ;
    END
  END north[30]
  PIN north[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 388.130 2240.120 388.410 2244.120 ;
    END
  END north[31]
  PIN north[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 399.170 2240.120 399.450 2244.120 ;
    END
  END north[32]
  PIN north[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 409.750 2240.120 410.030 2244.120 ;
    END
  END north[33]
  PIN north[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 420.330 2240.120 420.610 2244.120 ;
    END
  END north[34]
  PIN north[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 431.370 2240.120 431.650 2244.120 ;
    END
  END north[35]
  PIN north[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 441.950 2240.120 442.230 2244.120 ;
    END
  END north[36]
  PIN north[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 452.990 2240.120 453.270 2244.120 ;
    END
  END north[37]
  PIN north[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 463.570 2240.120 463.850 2244.120 ;
    END
  END north[38]
  PIN north[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 474.610 2240.120 474.890 2244.120 ;
    END
  END north[39]
  PIN north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 86.830 2240.120 87.110 2244.120 ;
    END
  END north[3]
  PIN north[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 485.190 2240.120 485.470 2244.120 ;
    END
  END north[40]
  PIN north[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 495.770 2240.120 496.050 2244.120 ;
    END
  END north[41]
  PIN north[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 506.810 2240.120 507.090 2244.120 ;
    END
  END north[42]
  PIN north[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 517.390 2240.120 517.670 2244.120 ;
    END
  END north[43]
  PIN north[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 528.430 2240.120 528.710 2244.120 ;
    END
  END north[44]
  PIN north[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 539.010 2240.120 539.290 2244.120 ;
    END
  END north[45]
  PIN north[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 549.590 2240.120 549.870 2244.120 ;
    END
  END north[46]
  PIN north[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 560.630 2240.120 560.910 2244.120 ;
    END
  END north[47]
  PIN north[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 571.210 2240.120 571.490 2244.120 ;
    END
  END north[48]
  PIN north[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 582.250 2240.120 582.530 2244.120 ;
    END
  END north[49]
  PIN north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 97.410 2240.120 97.690 2244.120 ;
    END
  END north[4]
  PIN north[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 592.830 2240.120 593.110 2244.120 ;
    END
  END north[50]
  PIN north[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 603.410 2240.120 603.690 2244.120 ;
    END
  END north[51]
  PIN north[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 614.450 2240.120 614.730 2244.120 ;
    END
  END north[52]
  PIN north[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 625.030 2240.120 625.310 2244.120 ;
    END
  END north[53]
  PIN north[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 636.070 2240.120 636.350 2244.120 ;
    END
  END north[54]
  PIN north[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 646.650 2240.120 646.930 2244.120 ;
    END
  END north[55]
  PIN north[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 657.230 2240.120 657.510 2244.120 ;
    END
  END north[56]
  PIN north[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 668.270 2240.120 668.550 2244.120 ;
    END
  END north[57]
  PIN north[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 678.850 2240.120 679.130 2244.120 ;
    END
  END north[58]
  PIN north[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 689.890 2240.120 690.170 2244.120 ;
    END
  END north[59]
  PIN north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 108.450 2240.120 108.730 2244.120 ;
    END
  END north[5]
  PIN north[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 700.470 2240.120 700.750 2244.120 ;
    END
  END north[60]
  PIN north[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 711.510 2240.120 711.790 2244.120 ;
    END
  END north[61]
  PIN north[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 722.090 2240.120 722.370 2244.120 ;
    END
  END north[62]
  PIN north[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 732.670 2240.120 732.950 2244.120 ;
    END
  END north[63]
  PIN north[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 743.710 2240.120 743.990 2244.120 ;
    END
  END north[64]
  PIN north[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 754.290 2240.120 754.570 2244.120 ;
    END
  END north[65]
  PIN north[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 765.330 2240.120 765.610 2244.120 ;
    END
  END north[66]
  PIN north[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 775.910 2240.120 776.190 2244.120 ;
    END
  END north[67]
  PIN north[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 786.490 2240.120 786.770 2244.120 ;
    END
  END north[68]
  PIN north[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 797.530 2240.120 797.810 2244.120 ;
    END
  END north[69]
  PIN north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 119.030 2240.120 119.310 2244.120 ;
    END
  END north[6]
  PIN north[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 808.110 2240.120 808.390 2244.120 ;
    END
  END north[70]
  PIN north[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 819.150 2240.120 819.430 2244.120 ;
    END
  END north[71]
  PIN north[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 829.730 2240.120 830.010 2244.120 ;
    END
  END north[72]
  PIN north[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 840.310 2240.120 840.590 2244.120 ;
    END
  END north[73]
  PIN north[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 851.350 2240.120 851.630 2244.120 ;
    END
  END north[74]
  PIN north[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 861.930 2240.120 862.210 2244.120 ;
    END
  END north[75]
  PIN north[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 872.970 2240.120 873.250 2244.120 ;
    END
  END north[76]
  PIN north[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 883.550 2240.120 883.830 2244.120 ;
    END
  END north[77]
  PIN north[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 894.590 2240.120 894.870 2244.120 ;
    END
  END north[78]
  PIN north[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 905.170 2240.120 905.450 2244.120 ;
    END
  END north[79]
  PIN north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 129.610 2240.120 129.890 2244.120 ;
    END
  END north[7]
  PIN north[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 915.750 2240.120 916.030 2244.120 ;
    END
  END north[80]
  PIN north[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 926.790 2240.120 927.070 2244.120 ;
    END
  END north[81]
  PIN north[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 937.370 2240.120 937.650 2244.120 ;
    END
  END north[82]
  PIN north[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 948.410 2240.120 948.690 2244.120 ;
    END
  END north[83]
  PIN north[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 958.990 2240.120 959.270 2244.120 ;
    END
  END north[84]
  PIN north[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 969.570 2240.120 969.850 2244.120 ;
    END
  END north[85]
  PIN north[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 980.610 2240.120 980.890 2244.120 ;
    END
  END north[86]
  PIN north[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 991.190 2240.120 991.470 2244.120 ;
    END
  END north[87]
  PIN north[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1002.230 2240.120 1002.510 2244.120 ;
    END
  END north[88]
  PIN north[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1012.810 2240.120 1013.090 2244.120 ;
    END
  END north[89]
  PIN north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 140.650 2240.120 140.930 2244.120 ;
    END
  END north[8]
  PIN north[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1023.390 2240.120 1023.670 2244.120 ;
    END
  END north[90]
  PIN north[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1034.430 2240.120 1034.710 2244.120 ;
    END
  END north[91]
  PIN north[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1045.010 2240.120 1045.290 2244.120 ;
    END
  END north[92]
  PIN north[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1056.050 2240.120 1056.330 2244.120 ;
    END
  END north[93]
  PIN north[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1066.630 2240.120 1066.910 2244.120 ;
    END
  END north[94]
  PIN north[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1077.210 2240.120 1077.490 2244.120 ;
    END
  END north[95]
  PIN north[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1088.250 2240.120 1088.530 2244.120 ;
    END
  END north[96]
  PIN north[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1098.830 2240.120 1099.110 2244.120 ;
    END
  END north[97]
  PIN north[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1109.870 2240.120 1110.150 2244.120 ;
    END
  END north[98]
  PIN north[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1120.450 2240.120 1120.730 2244.120 ;
    END
  END north[99]
  PIN north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 151.230 2240.120 151.510 2244.120 ;
    END
  END north[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2237.840 53.480 2238.440 ;
    END
  END rst
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2111.750 44.120 2112.030 48.120 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2143.490 2240.120 2143.770 2244.120 ;
    END
  END shift_out
  PIN south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.630 44.120 54.910 48.120 ;
    END
  END south[0]
  PIN south[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1114.930 44.120 1115.210 48.120 ;
    END
  END south[100]
  PIN south[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1125.510 44.120 1125.790 48.120 ;
    END
  END south[101]
  PIN south[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1136.090 44.120 1136.370 48.120 ;
    END
  END south[102]
  PIN south[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1146.670 44.120 1146.950 48.120 ;
    END
  END south[103]
  PIN south[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1157.250 44.120 1157.530 48.120 ;
    END
  END south[104]
  PIN south[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1167.830 44.120 1168.110 48.120 ;
    END
  END south[105]
  PIN south[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1178.410 44.120 1178.690 48.120 ;
    END
  END south[106]
  PIN south[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1188.990 44.120 1189.270 48.120 ;
    END
  END south[107]
  PIN south[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1200.030 44.120 1200.310 48.120 ;
    END
  END south[108]
  PIN south[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1210.610 44.120 1210.890 48.120 ;
    END
  END south[109]
  PIN south[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 160.430 44.120 160.710 48.120 ;
    END
  END south[10]
  PIN south[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1221.190 44.120 1221.470 48.120 ;
    END
  END south[110]
  PIN south[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1231.770 44.120 1232.050 48.120 ;
    END
  END south[111]
  PIN south[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1242.350 44.120 1242.630 48.120 ;
    END
  END south[112]
  PIN south[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1252.930 44.120 1253.210 48.120 ;
    END
  END south[113]
  PIN south[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1263.510 44.120 1263.790 48.120 ;
    END
  END south[114]
  PIN south[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1274.090 44.120 1274.370 48.120 ;
    END
  END south[115]
  PIN south[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1284.670 44.120 1284.950 48.120 ;
    END
  END south[116]
  PIN south[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1295.250 44.120 1295.530 48.120 ;
    END
  END south[117]
  PIN south[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1305.830 44.120 1306.110 48.120 ;
    END
  END south[118]
  PIN south[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1316.410 44.120 1316.690 48.120 ;
    END
  END south[119]
  PIN south[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 171.010 44.120 171.290 48.120 ;
    END
  END south[11]
  PIN south[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1326.990 44.120 1327.270 48.120 ;
    END
  END south[120]
  PIN south[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1337.570 44.120 1337.850 48.120 ;
    END
  END south[121]
  PIN south[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1348.150 44.120 1348.430 48.120 ;
    END
  END south[122]
  PIN south[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1358.730 44.120 1359.010 48.120 ;
    END
  END south[123]
  PIN south[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1369.310 44.120 1369.590 48.120 ;
    END
  END south[124]
  PIN south[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1379.890 44.120 1380.170 48.120 ;
    END
  END south[125]
  PIN south[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1390.930 44.120 1391.210 48.120 ;
    END
  END south[126]
  PIN south[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1401.510 44.120 1401.790 48.120 ;
    END
  END south[127]
  PIN south[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1412.090 44.120 1412.370 48.120 ;
    END
  END south[128]
  PIN south[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1422.670 44.120 1422.950 48.120 ;
    END
  END south[129]
  PIN south[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 181.590 44.120 181.870 48.120 ;
    END
  END south[12]
  PIN south[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1433.250 44.120 1433.530 48.120 ;
    END
  END south[130]
  PIN south[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1443.830 44.120 1444.110 48.120 ;
    END
  END south[131]
  PIN south[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1454.410 44.120 1454.690 48.120 ;
    END
  END south[132]
  PIN south[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1464.990 44.120 1465.270 48.120 ;
    END
  END south[133]
  PIN south[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1475.570 44.120 1475.850 48.120 ;
    END
  END south[134]
  PIN south[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1486.150 44.120 1486.430 48.120 ;
    END
  END south[135]
  PIN south[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1496.730 44.120 1497.010 48.120 ;
    END
  END south[136]
  PIN south[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1507.310 44.120 1507.590 48.120 ;
    END
  END south[137]
  PIN south[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1517.890 44.120 1518.170 48.120 ;
    END
  END south[138]
  PIN south[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1528.470 44.120 1528.750 48.120 ;
    END
  END south[139]
  PIN south[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 192.170 44.120 192.450 48.120 ;
    END
  END south[13]
  PIN south[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1539.050 44.120 1539.330 48.120 ;
    END
  END south[140]
  PIN south[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1549.630 44.120 1549.910 48.120 ;
    END
  END south[141]
  PIN south[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1560.210 44.120 1560.490 48.120 ;
    END
  END south[142]
  PIN south[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1570.790 44.120 1571.070 48.120 ;
    END
  END south[143]
  PIN south[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.830 44.120 1582.110 48.120 ;
    END
  END south[144]
  PIN south[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1592.410 44.120 1592.690 48.120 ;
    END
  END south[145]
  PIN south[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1602.990 44.120 1603.270 48.120 ;
    END
  END south[146]
  PIN south[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1613.570 44.120 1613.850 48.120 ;
    END
  END south[147]
  PIN south[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1624.150 44.120 1624.430 48.120 ;
    END
  END south[148]
  PIN south[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1634.730 44.120 1635.010 48.120 ;
    END
  END south[149]
  PIN south[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 202.750 44.120 203.030 48.120 ;
    END
  END south[14]
  PIN south[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1645.310 44.120 1645.590 48.120 ;
    END
  END south[150]
  PIN south[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1655.890 44.120 1656.170 48.120 ;
    END
  END south[151]
  PIN south[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1666.470 44.120 1666.750 48.120 ;
    END
  END south[152]
  PIN south[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1677.050 44.120 1677.330 48.120 ;
    END
  END south[153]
  PIN south[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1687.630 44.120 1687.910 48.120 ;
    END
  END south[154]
  PIN south[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1698.210 44.120 1698.490 48.120 ;
    END
  END south[155]
  PIN south[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1708.790 44.120 1709.070 48.120 ;
    END
  END south[156]
  PIN south[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1719.370 44.120 1719.650 48.120 ;
    END
  END south[157]
  PIN south[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1729.950 44.120 1730.230 48.120 ;
    END
  END south[158]
  PIN south[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1740.530 44.120 1740.810 48.120 ;
    END
  END south[159]
  PIN south[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 213.330 44.120 213.610 48.120 ;
    END
  END south[15]
  PIN south[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1751.110 44.120 1751.390 48.120 ;
    END
  END south[160]
  PIN south[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1761.690 44.120 1761.970 48.120 ;
    END
  END south[161]
  PIN south[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1772.730 44.120 1773.010 48.120 ;
    END
  END south[162]
  PIN south[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1783.310 44.120 1783.590 48.120 ;
    END
  END south[163]
  PIN south[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1793.890 44.120 1794.170 48.120 ;
    END
  END south[164]
  PIN south[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1804.470 44.120 1804.750 48.120 ;
    END
  END south[165]
  PIN south[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1815.050 44.120 1815.330 48.120 ;
    END
  END south[166]
  PIN south[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1825.630 44.120 1825.910 48.120 ;
    END
  END south[167]
  PIN south[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1836.210 44.120 1836.490 48.120 ;
    END
  END south[168]
  PIN south[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1846.790 44.120 1847.070 48.120 ;
    END
  END south[169]
  PIN south[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 223.910 44.120 224.190 48.120 ;
    END
  END south[16]
  PIN south[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1857.370 44.120 1857.650 48.120 ;
    END
  END south[170]
  PIN south[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1867.950 44.120 1868.230 48.120 ;
    END
  END south[171]
  PIN south[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1878.530 44.120 1878.810 48.120 ;
    END
  END south[172]
  PIN south[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1889.110 44.120 1889.390 48.120 ;
    END
  END south[173]
  PIN south[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1899.690 44.120 1899.970 48.120 ;
    END
  END south[174]
  PIN south[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1910.270 44.120 1910.550 48.120 ;
    END
  END south[175]
  PIN south[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1920.850 44.120 1921.130 48.120 ;
    END
  END south[176]
  PIN south[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1931.430 44.120 1931.710 48.120 ;
    END
  END south[177]
  PIN south[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1942.010 44.120 1942.290 48.120 ;
    END
  END south[178]
  PIN south[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1952.590 44.120 1952.870 48.120 ;
    END
  END south[179]
  PIN south[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 234.490 44.120 234.770 48.120 ;
    END
  END south[17]
  PIN south[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1963.630 44.120 1963.910 48.120 ;
    END
  END south[180]
  PIN south[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1974.210 44.120 1974.490 48.120 ;
    END
  END south[181]
  PIN south[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1984.790 44.120 1985.070 48.120 ;
    END
  END south[182]
  PIN south[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1995.370 44.120 1995.650 48.120 ;
    END
  END south[183]
  PIN south[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2005.950 44.120 2006.230 48.120 ;
    END
  END south[184]
  PIN south[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2016.530 44.120 2016.810 48.120 ;
    END
  END south[185]
  PIN south[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2027.110 44.120 2027.390 48.120 ;
    END
  END south[186]
  PIN south[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2037.690 44.120 2037.970 48.120 ;
    END
  END south[187]
  PIN south[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2048.270 44.120 2048.550 48.120 ;
    END
  END south[188]
  PIN south[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2058.850 44.120 2059.130 48.120 ;
    END
  END south[189]
  PIN south[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 245.530 44.120 245.810 48.120 ;
    END
  END south[18]
  PIN south[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2069.430 44.120 2069.710 48.120 ;
    END
  END south[190]
  PIN south[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2080.010 44.120 2080.290 48.120 ;
    END
  END south[191]
  PIN south[192]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2090.590 44.120 2090.870 48.120 ;
    END
  END south[192]
  PIN south[193]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2101.170 44.120 2101.450 48.120 ;
    END
  END south[193]
  PIN south[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 256.110 44.120 256.390 48.120 ;
    END
  END south[19]
  PIN south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 65.210 44.120 65.490 48.120 ;
    END
  END south[1]
  PIN south[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 266.690 44.120 266.970 48.120 ;
    END
  END south[20]
  PIN south[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 277.270 44.120 277.550 48.120 ;
    END
  END south[21]
  PIN south[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 287.850 44.120 288.130 48.120 ;
    END
  END south[22]
  PIN south[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 298.430 44.120 298.710 48.120 ;
    END
  END south[23]
  PIN south[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 309.010 44.120 309.290 48.120 ;
    END
  END south[24]
  PIN south[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 319.590 44.120 319.870 48.120 ;
    END
  END south[25]
  PIN south[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 330.170 44.120 330.450 48.120 ;
    END
  END south[26]
  PIN south[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 340.750 44.120 341.030 48.120 ;
    END
  END south[27]
  PIN south[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 351.330 44.120 351.610 48.120 ;
    END
  END south[28]
  PIN south[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 361.910 44.120 362.190 48.120 ;
    END
  END south[29]
  PIN south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.790 44.120 76.070 48.120 ;
    END
  END south[2]
  PIN south[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 372.490 44.120 372.770 48.120 ;
    END
  END south[30]
  PIN south[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 383.070 44.120 383.350 48.120 ;
    END
  END south[31]
  PIN south[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 393.650 44.120 393.930 48.120 ;
    END
  END south[32]
  PIN south[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 404.230 44.120 404.510 48.120 ;
    END
  END south[33]
  PIN south[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 414.810 44.120 415.090 48.120 ;
    END
  END south[34]
  PIN south[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 425.390 44.120 425.670 48.120 ;
    END
  END south[35]
  PIN south[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 436.430 44.120 436.710 48.120 ;
    END
  END south[36]
  PIN south[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 447.010 44.120 447.290 48.120 ;
    END
  END south[37]
  PIN south[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 457.590 44.120 457.870 48.120 ;
    END
  END south[38]
  PIN south[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 468.170 44.120 468.450 48.120 ;
    END
  END south[39]
  PIN south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 86.370 44.120 86.650 48.120 ;
    END
  END south[3]
  PIN south[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 478.750 44.120 479.030 48.120 ;
    END
  END south[40]
  PIN south[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 489.330 44.120 489.610 48.120 ;
    END
  END south[41]
  PIN south[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 499.910 44.120 500.190 48.120 ;
    END
  END south[42]
  PIN south[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 510.490 44.120 510.770 48.120 ;
    END
  END south[43]
  PIN south[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 521.070 44.120 521.350 48.120 ;
    END
  END south[44]
  PIN south[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 531.650 44.120 531.930 48.120 ;
    END
  END south[45]
  PIN south[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 542.230 44.120 542.510 48.120 ;
    END
  END south[46]
  PIN south[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 552.810 44.120 553.090 48.120 ;
    END
  END south[47]
  PIN south[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 563.390 44.120 563.670 48.120 ;
    END
  END south[48]
  PIN south[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 573.970 44.120 574.250 48.120 ;
    END
  END south[49]
  PIN south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 96.950 44.120 97.230 48.120 ;
    END
  END south[4]
  PIN south[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 584.550 44.120 584.830 48.120 ;
    END
  END south[50]
  PIN south[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 595.130 44.120 595.410 48.120 ;
    END
  END south[51]
  PIN south[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.710 44.120 605.990 48.120 ;
    END
  END south[52]
  PIN south[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 616.290 44.120 616.570 48.120 ;
    END
  END south[53]
  PIN south[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 627.330 44.120 627.610 48.120 ;
    END
  END south[54]
  PIN south[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 637.910 44.120 638.190 48.120 ;
    END
  END south[55]
  PIN south[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 648.490 44.120 648.770 48.120 ;
    END
  END south[56]
  PIN south[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 659.070 44.120 659.350 48.120 ;
    END
  END south[57]
  PIN south[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 669.650 44.120 669.930 48.120 ;
    END
  END south[58]
  PIN south[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 680.230 44.120 680.510 48.120 ;
    END
  END south[59]
  PIN south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 107.530 44.120 107.810 48.120 ;
    END
  END south[5]
  PIN south[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 690.810 44.120 691.090 48.120 ;
    END
  END south[60]
  PIN south[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 701.390 44.120 701.670 48.120 ;
    END
  END south[61]
  PIN south[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 711.970 44.120 712.250 48.120 ;
    END
  END south[62]
  PIN south[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 722.550 44.120 722.830 48.120 ;
    END
  END south[63]
  PIN south[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 733.130 44.120 733.410 48.120 ;
    END
  END south[64]
  PIN south[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 743.710 44.120 743.990 48.120 ;
    END
  END south[65]
  PIN south[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 754.290 44.120 754.570 48.120 ;
    END
  END south[66]
  PIN south[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 764.870 44.120 765.150 48.120 ;
    END
  END south[67]
  PIN south[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 775.450 44.120 775.730 48.120 ;
    END
  END south[68]
  PIN south[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 786.030 44.120 786.310 48.120 ;
    END
  END south[69]
  PIN south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 118.110 44.120 118.390 48.120 ;
    END
  END south[6]
  PIN south[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 796.610 44.120 796.890 48.120 ;
    END
  END south[70]
  PIN south[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 807.190 44.120 807.470 48.120 ;
    END
  END south[71]
  PIN south[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 818.230 44.120 818.510 48.120 ;
    END
  END south[72]
  PIN south[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 828.810 44.120 829.090 48.120 ;
    END
  END south[73]
  PIN south[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 839.390 44.120 839.670 48.120 ;
    END
  END south[74]
  PIN south[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 849.970 44.120 850.250 48.120 ;
    END
  END south[75]
  PIN south[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 860.550 44.120 860.830 48.120 ;
    END
  END south[76]
  PIN south[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 871.130 44.120 871.410 48.120 ;
    END
  END south[77]
  PIN south[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 881.710 44.120 881.990 48.120 ;
    END
  END south[78]
  PIN south[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 892.290 44.120 892.570 48.120 ;
    END
  END south[79]
  PIN south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 128.690 44.120 128.970 48.120 ;
    END
  END south[7]
  PIN south[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 902.870 44.120 903.150 48.120 ;
    END
  END south[80]
  PIN south[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 913.450 44.120 913.730 48.120 ;
    END
  END south[81]
  PIN south[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 924.030 44.120 924.310 48.120 ;
    END
  END south[82]
  PIN south[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 934.610 44.120 934.890 48.120 ;
    END
  END south[83]
  PIN south[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 945.190 44.120 945.470 48.120 ;
    END
  END south[84]
  PIN south[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 955.770 44.120 956.050 48.120 ;
    END
  END south[85]
  PIN south[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 966.350 44.120 966.630 48.120 ;
    END
  END south[86]
  PIN south[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 976.930 44.120 977.210 48.120 ;
    END
  END south[87]
  PIN south[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 987.510 44.120 987.790 48.120 ;
    END
  END south[88]
  PIN south[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 998.090 44.120 998.370 48.120 ;
    END
  END south[89]
  PIN south[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 139.270 44.120 139.550 48.120 ;
    END
  END south[8]
  PIN south[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1009.130 44.120 1009.410 48.120 ;
    END
  END south[90]
  PIN south[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1019.710 44.120 1019.990 48.120 ;
    END
  END south[91]
  PIN south[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1030.290 44.120 1030.570 48.120 ;
    END
  END south[92]
  PIN south[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1040.870 44.120 1041.150 48.120 ;
    END
  END south[93]
  PIN south[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1051.450 44.120 1051.730 48.120 ;
    END
  END south[94]
  PIN south[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1062.030 44.120 1062.310 48.120 ;
    END
  END south[95]
  PIN south[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1072.610 44.120 1072.890 48.120 ;
    END
  END south[96]
  PIN south[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1083.190 44.120 1083.470 48.120 ;
    END
  END south[97]
  PIN south[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1093.770 44.120 1094.050 48.120 ;
    END
  END south[98]
  PIN south[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1104.350 44.120 1104.630 48.120 ;
    END
  END south[99]
  PIN south[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 149.850 44.120 150.130 48.120 ;
    END
  END south[9]
  PIN west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 49.600 53.480 50.200 ;
    END
  END west[0]
  PIN west[100]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1171.600 53.480 1172.200 ;
    END
  END west[100]
  PIN west[101]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1183.160 53.480 1183.760 ;
    END
  END west[101]
  PIN west[102]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1194.040 53.480 1194.640 ;
    END
  END west[102]
  PIN west[103]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1205.600 53.480 1206.200 ;
    END
  END west[103]
  PIN west[104]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1216.480 53.480 1217.080 ;
    END
  END west[104]
  PIN west[105]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1228.040 53.480 1228.640 ;
    END
  END west[105]
  PIN west[106]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1238.920 53.480 1239.520 ;
    END
  END west[106]
  PIN west[107]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1250.480 53.480 1251.080 ;
    END
  END west[107]
  PIN west[108]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1261.360 53.480 1261.960 ;
    END
  END west[108]
  PIN west[109]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1272.920 53.480 1273.520 ;
    END
  END west[109]
  PIN west[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 161.800 53.480 162.400 ;
    END
  END west[10]
  PIN west[110]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1283.800 53.480 1284.400 ;
    END
  END west[110]
  PIN west[111]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1295.360 53.480 1295.960 ;
    END
  END west[111]
  PIN west[112]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1306.240 53.480 1306.840 ;
    END
  END west[112]
  PIN west[113]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1317.800 53.480 1318.400 ;
    END
  END west[113]
  PIN west[114]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1328.680 53.480 1329.280 ;
    END
  END west[114]
  PIN west[115]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1340.240 53.480 1340.840 ;
    END
  END west[115]
  PIN west[116]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1351.120 53.480 1351.720 ;
    END
  END west[116]
  PIN west[117]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1362.680 53.480 1363.280 ;
    END
  END west[117]
  PIN west[118]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1373.560 53.480 1374.160 ;
    END
  END west[118]
  PIN west[119]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1385.120 53.480 1385.720 ;
    END
  END west[119]
  PIN west[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 172.680 53.480 173.280 ;
    END
  END west[11]
  PIN west[120]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1396.000 53.480 1396.600 ;
    END
  END west[120]
  PIN west[121]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1407.560 53.480 1408.160 ;
    END
  END west[121]
  PIN west[122]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1418.440 53.480 1419.040 ;
    END
  END west[122]
  PIN west[123]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1430.000 53.480 1430.600 ;
    END
  END west[123]
  PIN west[124]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1440.880 53.480 1441.480 ;
    END
  END west[124]
  PIN west[125]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1452.440 53.480 1453.040 ;
    END
  END west[125]
  PIN west[126]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1463.320 53.480 1463.920 ;
    END
  END west[126]
  PIN west[127]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1474.880 53.480 1475.480 ;
    END
  END west[127]
  PIN west[128]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1485.760 53.480 1486.360 ;
    END
  END west[128]
  PIN west[129]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1497.320 53.480 1497.920 ;
    END
  END west[129]
  PIN west[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 184.240 53.480 184.840 ;
    END
  END west[12]
  PIN west[130]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1508.200 53.480 1508.800 ;
    END
  END west[130]
  PIN west[131]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1519.760 53.480 1520.360 ;
    END
  END west[131]
  PIN west[132]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1530.640 53.480 1531.240 ;
    END
  END west[132]
  PIN west[133]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1542.200 53.480 1542.800 ;
    END
  END west[133]
  PIN west[134]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1553.080 53.480 1553.680 ;
    END
  END west[134]
  PIN west[135]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1564.640 53.480 1565.240 ;
    END
  END west[135]
  PIN west[136]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1575.520 53.480 1576.120 ;
    END
  END west[136]
  PIN west[137]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1587.080 53.480 1587.680 ;
    END
  END west[137]
  PIN west[138]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1597.960 53.480 1598.560 ;
    END
  END west[138]
  PIN west[139]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1609.520 53.480 1610.120 ;
    END
  END west[139]
  PIN west[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 195.120 53.480 195.720 ;
    END
  END west[13]
  PIN west[140]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1620.400 53.480 1621.000 ;
    END
  END west[140]
  PIN west[141]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1631.960 53.480 1632.560 ;
    END
  END west[141]
  PIN west[142]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1642.840 53.480 1643.440 ;
    END
  END west[142]
  PIN west[143]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1654.400 53.480 1655.000 ;
    END
  END west[143]
  PIN west[144]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1665.280 53.480 1665.880 ;
    END
  END west[144]
  PIN west[145]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1676.840 53.480 1677.440 ;
    END
  END west[145]
  PIN west[146]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1687.720 53.480 1688.320 ;
    END
  END west[146]
  PIN west[147]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1699.280 53.480 1699.880 ;
    END
  END west[147]
  PIN west[148]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1710.160 53.480 1710.760 ;
    END
  END west[148]
  PIN west[149]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1721.720 53.480 1722.320 ;
    END
  END west[149]
  PIN west[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 206.680 53.480 207.280 ;
    END
  END west[14]
  PIN west[150]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1732.600 53.480 1733.200 ;
    END
  END west[150]
  PIN west[151]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1744.160 53.480 1744.760 ;
    END
  END west[151]
  PIN west[152]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1755.040 53.480 1755.640 ;
    END
  END west[152]
  PIN west[153]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1766.600 53.480 1767.200 ;
    END
  END west[153]
  PIN west[154]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1777.480 53.480 1778.080 ;
    END
  END west[154]
  PIN west[155]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1789.040 53.480 1789.640 ;
    END
  END west[155]
  PIN west[156]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1799.920 53.480 1800.520 ;
    END
  END west[156]
  PIN west[157]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1811.480 53.480 1812.080 ;
    END
  END west[157]
  PIN west[158]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1822.360 53.480 1822.960 ;
    END
  END west[158]
  PIN west[159]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1833.920 53.480 1834.520 ;
    END
  END west[159]
  PIN west[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 217.560 53.480 218.160 ;
    END
  END west[15]
  PIN west[160]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1844.800 53.480 1845.400 ;
    END
  END west[160]
  PIN west[161]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1856.360 53.480 1856.960 ;
    END
  END west[161]
  PIN west[162]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1867.240 53.480 1867.840 ;
    END
  END west[162]
  PIN west[163]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1878.800 53.480 1879.400 ;
    END
  END west[163]
  PIN west[164]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1889.680 53.480 1890.280 ;
    END
  END west[164]
  PIN west[165]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1901.240 53.480 1901.840 ;
    END
  END west[165]
  PIN west[166]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1912.120 53.480 1912.720 ;
    END
  END west[166]
  PIN west[167]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1923.680 53.480 1924.280 ;
    END
  END west[167]
  PIN west[168]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1934.560 53.480 1935.160 ;
    END
  END west[168]
  PIN west[169]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1946.120 53.480 1946.720 ;
    END
  END west[169]
  PIN west[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 229.120 53.480 229.720 ;
    END
  END west[16]
  PIN west[170]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1957.000 53.480 1957.600 ;
    END
  END west[170]
  PIN west[171]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1968.560 53.480 1969.160 ;
    END
  END west[171]
  PIN west[172]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1979.440 53.480 1980.040 ;
    END
  END west[172]
  PIN west[173]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1991.000 53.480 1991.600 ;
    END
  END west[173]
  PIN west[174]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2001.880 53.480 2002.480 ;
    END
  END west[174]
  PIN west[175]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2013.440 53.480 2014.040 ;
    END
  END west[175]
  PIN west[176]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2024.320 53.480 2024.920 ;
    END
  END west[176]
  PIN west[177]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2035.880 53.480 2036.480 ;
    END
  END west[177]
  PIN west[178]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2046.760 53.480 2047.360 ;
    END
  END west[178]
  PIN west[179]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2058.320 53.480 2058.920 ;
    END
  END west[179]
  PIN west[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 240.000 53.480 240.600 ;
    END
  END west[17]
  PIN west[180]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2069.200 53.480 2069.800 ;
    END
  END west[180]
  PIN west[181]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2080.760 53.480 2081.360 ;
    END
  END west[181]
  PIN west[182]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2091.640 53.480 2092.240 ;
    END
  END west[182]
  PIN west[183]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2103.200 53.480 2103.800 ;
    END
  END west[183]
  PIN west[184]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2114.080 53.480 2114.680 ;
    END
  END west[184]
  PIN west[185]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2125.640 53.480 2126.240 ;
    END
  END west[185]
  PIN west[186]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2136.520 53.480 2137.120 ;
    END
  END west[186]
  PIN west[187]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2148.080 53.480 2148.680 ;
    END
  END west[187]
  PIN west[188]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2158.960 53.480 2159.560 ;
    END
  END west[188]
  PIN west[189]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2170.520 53.480 2171.120 ;
    END
  END west[189]
  PIN west[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 251.560 53.480 252.160 ;
    END
  END west[18]
  PIN west[190]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2181.400 53.480 2182.000 ;
    END
  END west[190]
  PIN west[191]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2192.960 53.480 2193.560 ;
    END
  END west[191]
  PIN west[192]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2203.840 53.480 2204.440 ;
    END
  END west[192]
  PIN west[193]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2215.400 53.480 2216.000 ;
    END
  END west[193]
  PIN west[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 262.440 53.480 263.040 ;
    END
  END west[19]
  PIN west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 60.480 53.480 61.080 ;
    END
  END west[1]
  PIN west[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 274.000 53.480 274.600 ;
    END
  END west[20]
  PIN west[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 284.880 53.480 285.480 ;
    END
  END west[21]
  PIN west[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 296.440 53.480 297.040 ;
    END
  END west[22]
  PIN west[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 307.320 53.480 307.920 ;
    END
  END west[23]
  PIN west[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 318.880 53.480 319.480 ;
    END
  END west[24]
  PIN west[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 329.760 53.480 330.360 ;
    END
  END west[25]
  PIN west[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 341.320 53.480 341.920 ;
    END
  END west[26]
  PIN west[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 352.200 53.480 352.800 ;
    END
  END west[27]
  PIN west[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 363.760 53.480 364.360 ;
    END
  END west[28]
  PIN west[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 374.640 53.480 375.240 ;
    END
  END west[29]
  PIN west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 72.040 53.480 72.640 ;
    END
  END west[2]
  PIN west[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 386.200 53.480 386.800 ;
    END
  END west[30]
  PIN west[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 397.080 53.480 397.680 ;
    END
  END west[31]
  PIN west[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 408.640 53.480 409.240 ;
    END
  END west[32]
  PIN west[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 419.520 53.480 420.120 ;
    END
  END west[33]
  PIN west[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 431.080 53.480 431.680 ;
    END
  END west[34]
  PIN west[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 441.960 53.480 442.560 ;
    END
  END west[35]
  PIN west[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 453.520 53.480 454.120 ;
    END
  END west[36]
  PIN west[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 464.400 53.480 465.000 ;
    END
  END west[37]
  PIN west[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 475.960 53.480 476.560 ;
    END
  END west[38]
  PIN west[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 486.840 53.480 487.440 ;
    END
  END west[39]
  PIN west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 82.920 53.480 83.520 ;
    END
  END west[3]
  PIN west[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 498.400 53.480 499.000 ;
    END
  END west[40]
  PIN west[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 509.280 53.480 509.880 ;
    END
  END west[41]
  PIN west[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 520.840 53.480 521.440 ;
    END
  END west[42]
  PIN west[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 531.720 53.480 532.320 ;
    END
  END west[43]
  PIN west[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 543.280 53.480 543.880 ;
    END
  END west[44]
  PIN west[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 554.160 53.480 554.760 ;
    END
  END west[45]
  PIN west[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 565.720 53.480 566.320 ;
    END
  END west[46]
  PIN west[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 576.600 53.480 577.200 ;
    END
  END west[47]
  PIN west[48]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 588.160 53.480 588.760 ;
    END
  END west[48]
  PIN west[49]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 599.040 53.480 599.640 ;
    END
  END west[49]
  PIN west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 94.480 53.480 95.080 ;
    END
  END west[4]
  PIN west[50]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 610.600 53.480 611.200 ;
    END
  END west[50]
  PIN west[51]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 621.480 53.480 622.080 ;
    END
  END west[51]
  PIN west[52]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 633.040 53.480 633.640 ;
    END
  END west[52]
  PIN west[53]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 643.920 53.480 644.520 ;
    END
  END west[53]
  PIN west[54]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 655.480 53.480 656.080 ;
    END
  END west[54]
  PIN west[55]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 666.360 53.480 666.960 ;
    END
  END west[55]
  PIN west[56]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 677.920 53.480 678.520 ;
    END
  END west[56]
  PIN west[57]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 688.800 53.480 689.400 ;
    END
  END west[57]
  PIN west[58]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 700.360 53.480 700.960 ;
    END
  END west[58]
  PIN west[59]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 711.240 53.480 711.840 ;
    END
  END west[59]
  PIN west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 105.360 53.480 105.960 ;
    END
  END west[5]
  PIN west[60]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 722.800 53.480 723.400 ;
    END
  END west[60]
  PIN west[61]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 733.680 53.480 734.280 ;
    END
  END west[61]
  PIN west[62]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 745.240 53.480 745.840 ;
    END
  END west[62]
  PIN west[63]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 756.120 53.480 756.720 ;
    END
  END west[63]
  PIN west[64]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 767.680 53.480 768.280 ;
    END
  END west[64]
  PIN west[65]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 778.560 53.480 779.160 ;
    END
  END west[65]
  PIN west[66]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 790.120 53.480 790.720 ;
    END
  END west[66]
  PIN west[67]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 801.000 53.480 801.600 ;
    END
  END west[67]
  PIN west[68]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 812.560 53.480 813.160 ;
    END
  END west[68]
  PIN west[69]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 823.440 53.480 824.040 ;
    END
  END west[69]
  PIN west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 116.920 53.480 117.520 ;
    END
  END west[6]
  PIN west[70]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 835.000 53.480 835.600 ;
    END
  END west[70]
  PIN west[71]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 845.880 53.480 846.480 ;
    END
  END west[71]
  PIN west[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 857.440 53.480 858.040 ;
    END
  END west[72]
  PIN west[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 868.320 53.480 868.920 ;
    END
  END west[73]
  PIN west[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 879.880 53.480 880.480 ;
    END
  END west[74]
  PIN west[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 890.760 53.480 891.360 ;
    END
  END west[75]
  PIN west[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 902.320 53.480 902.920 ;
    END
  END west[76]
  PIN west[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 913.200 53.480 913.800 ;
    END
  END west[77]
  PIN west[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 924.760 53.480 925.360 ;
    END
  END west[78]
  PIN west[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 935.640 53.480 936.240 ;
    END
  END west[79]
  PIN west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 127.800 53.480 128.400 ;
    END
  END west[7]
  PIN west[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 947.200 53.480 947.800 ;
    END
  END west[80]
  PIN west[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 958.080 53.480 958.680 ;
    END
  END west[81]
  PIN west[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 969.640 53.480 970.240 ;
    END
  END west[82]
  PIN west[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 980.520 53.480 981.120 ;
    END
  END west[83]
  PIN west[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 992.080 53.480 992.680 ;
    END
  END west[84]
  PIN west[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1002.960 53.480 1003.560 ;
    END
  END west[85]
  PIN west[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1014.520 53.480 1015.120 ;
    END
  END west[86]
  PIN west[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1025.400 53.480 1026.000 ;
    END
  END west[87]
  PIN west[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1036.960 53.480 1037.560 ;
    END
  END west[88]
  PIN west[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1047.840 53.480 1048.440 ;
    END
  END west[89]
  PIN west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 139.360 53.480 139.960 ;
    END
  END west[8]
  PIN west[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1059.400 53.480 1060.000 ;
    END
  END west[90]
  PIN west[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1070.280 53.480 1070.880 ;
    END
  END west[91]
  PIN west[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1081.840 53.480 1082.440 ;
    END
  END west[92]
  PIN west[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1092.720 53.480 1093.320 ;
    END
  END west[93]
  PIN west[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1104.280 53.480 1104.880 ;
    END
  END west[94]
  PIN west[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1115.160 53.480 1115.760 ;
    END
  END west[95]
  PIN west[96]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1126.720 53.480 1127.320 ;
    END
  END west[96]
  PIN west[97]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1137.600 53.480 1138.200 ;
    END
  END west[97]
  PIN west[98]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1149.160 53.480 1149.760 ;
    END
  END west[98]
  PIN west[99]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1160.720 53.480 1161.320 ;
    END
  END west[99]
  PIN west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 150.240 53.480 150.840 ;
    END
  END west[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2173.860 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2198.860 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 2143.860 2231.085 ;
      LAYER met1 ;
        RECT 55.000 45.860 2143.860 2239.800 ;
      LAYER met2 ;
        RECT 55.190 2239.840 64.930 2240.120 ;
        RECT 65.770 2239.840 75.510 2240.120 ;
        RECT 76.350 2239.840 86.550 2240.120 ;
        RECT 87.390 2239.840 97.130 2240.120 ;
        RECT 97.970 2239.840 108.170 2240.120 ;
        RECT 109.010 2239.840 118.750 2240.120 ;
        RECT 119.590 2239.840 129.330 2240.120 ;
        RECT 130.170 2239.840 140.370 2240.120 ;
        RECT 141.210 2239.840 150.950 2240.120 ;
        RECT 151.790 2239.840 161.990 2240.120 ;
        RECT 162.830 2239.840 172.570 2240.120 ;
        RECT 173.410 2239.840 183.150 2240.120 ;
        RECT 183.990 2239.840 194.190 2240.120 ;
        RECT 195.030 2239.840 204.770 2240.120 ;
        RECT 205.610 2239.840 215.810 2240.120 ;
        RECT 216.650 2239.840 226.390 2240.120 ;
        RECT 227.230 2239.840 236.970 2240.120 ;
        RECT 237.810 2239.840 248.010 2240.120 ;
        RECT 248.850 2239.840 258.590 2240.120 ;
        RECT 259.430 2239.840 269.630 2240.120 ;
        RECT 270.470 2239.840 280.210 2240.120 ;
        RECT 281.050 2239.840 291.250 2240.120 ;
        RECT 292.090 2239.840 301.830 2240.120 ;
        RECT 302.670 2239.840 312.410 2240.120 ;
        RECT 313.250 2239.840 323.450 2240.120 ;
        RECT 324.290 2239.840 334.030 2240.120 ;
        RECT 334.870 2239.840 345.070 2240.120 ;
        RECT 345.910 2239.840 355.650 2240.120 ;
        RECT 356.490 2239.840 366.230 2240.120 ;
        RECT 367.070 2239.840 377.270 2240.120 ;
        RECT 378.110 2239.840 387.850 2240.120 ;
        RECT 388.690 2239.840 398.890 2240.120 ;
        RECT 399.730 2239.840 409.470 2240.120 ;
        RECT 410.310 2239.840 420.050 2240.120 ;
        RECT 420.890 2239.840 431.090 2240.120 ;
        RECT 431.930 2239.840 441.670 2240.120 ;
        RECT 442.510 2239.840 452.710 2240.120 ;
        RECT 453.550 2239.840 463.290 2240.120 ;
        RECT 464.130 2239.840 474.330 2240.120 ;
        RECT 475.170 2239.840 484.910 2240.120 ;
        RECT 485.750 2239.840 495.490 2240.120 ;
        RECT 496.330 2239.840 506.530 2240.120 ;
        RECT 507.370 2239.840 517.110 2240.120 ;
        RECT 517.950 2239.840 528.150 2240.120 ;
        RECT 528.990 2239.840 538.730 2240.120 ;
        RECT 539.570 2239.840 549.310 2240.120 ;
        RECT 550.150 2239.840 560.350 2240.120 ;
        RECT 561.190 2239.840 570.930 2240.120 ;
        RECT 571.770 2239.840 581.970 2240.120 ;
        RECT 582.810 2239.840 592.550 2240.120 ;
        RECT 593.390 2239.840 603.130 2240.120 ;
        RECT 603.970 2239.840 614.170 2240.120 ;
        RECT 615.010 2239.840 624.750 2240.120 ;
        RECT 625.590 2239.840 635.790 2240.120 ;
        RECT 636.630 2239.840 646.370 2240.120 ;
        RECT 647.210 2239.840 656.950 2240.120 ;
        RECT 657.790 2239.840 667.990 2240.120 ;
        RECT 668.830 2239.840 678.570 2240.120 ;
        RECT 679.410 2239.840 689.610 2240.120 ;
        RECT 690.450 2239.840 700.190 2240.120 ;
        RECT 701.030 2239.840 711.230 2240.120 ;
        RECT 712.070 2239.840 721.810 2240.120 ;
        RECT 722.650 2239.840 732.390 2240.120 ;
        RECT 733.230 2239.840 743.430 2240.120 ;
        RECT 744.270 2239.840 754.010 2240.120 ;
        RECT 754.850 2239.840 765.050 2240.120 ;
        RECT 765.890 2239.840 775.630 2240.120 ;
        RECT 776.470 2239.840 786.210 2240.120 ;
        RECT 787.050 2239.840 797.250 2240.120 ;
        RECT 798.090 2239.840 807.830 2240.120 ;
        RECT 808.670 2239.840 818.870 2240.120 ;
        RECT 819.710 2239.840 829.450 2240.120 ;
        RECT 830.290 2239.840 840.030 2240.120 ;
        RECT 840.870 2239.840 851.070 2240.120 ;
        RECT 851.910 2239.840 861.650 2240.120 ;
        RECT 862.490 2239.840 872.690 2240.120 ;
        RECT 873.530 2239.840 883.270 2240.120 ;
        RECT 884.110 2239.840 894.310 2240.120 ;
        RECT 895.150 2239.840 904.890 2240.120 ;
        RECT 905.730 2239.840 915.470 2240.120 ;
        RECT 916.310 2239.840 926.510 2240.120 ;
        RECT 927.350 2239.840 937.090 2240.120 ;
        RECT 937.930 2239.840 948.130 2240.120 ;
        RECT 948.970 2239.840 958.710 2240.120 ;
        RECT 959.550 2239.840 969.290 2240.120 ;
        RECT 970.130 2239.840 980.330 2240.120 ;
        RECT 981.170 2239.840 990.910 2240.120 ;
        RECT 991.750 2239.840 1001.950 2240.120 ;
        RECT 1002.790 2239.840 1012.530 2240.120 ;
        RECT 1013.370 2239.840 1023.110 2240.120 ;
        RECT 1023.950 2239.840 1034.150 2240.120 ;
        RECT 1034.990 2239.840 1044.730 2240.120 ;
        RECT 1045.570 2239.840 1055.770 2240.120 ;
        RECT 1056.610 2239.840 1066.350 2240.120 ;
        RECT 1067.190 2239.840 1076.930 2240.120 ;
        RECT 1077.770 2239.840 1087.970 2240.120 ;
        RECT 1088.810 2239.840 1098.550 2240.120 ;
        RECT 1099.390 2239.840 1109.590 2240.120 ;
        RECT 1110.430 2239.840 1120.170 2240.120 ;
        RECT 1121.010 2239.840 1131.210 2240.120 ;
        RECT 1132.050 2239.840 1141.790 2240.120 ;
        RECT 1142.630 2239.840 1152.370 2240.120 ;
        RECT 1153.210 2239.840 1163.410 2240.120 ;
        RECT 1164.250 2239.840 1173.990 2240.120 ;
        RECT 1174.830 2239.840 1185.030 2240.120 ;
        RECT 1185.870 2239.840 1195.610 2240.120 ;
        RECT 1196.450 2239.840 1206.190 2240.120 ;
        RECT 1207.030 2239.840 1217.230 2240.120 ;
        RECT 1218.070 2239.840 1227.810 2240.120 ;
        RECT 1228.650 2239.840 1238.850 2240.120 ;
        RECT 1239.690 2239.840 1249.430 2240.120 ;
        RECT 1250.270 2239.840 1260.010 2240.120 ;
        RECT 1260.850 2239.840 1271.050 2240.120 ;
        RECT 1271.890 2239.840 1281.630 2240.120 ;
        RECT 1282.470 2239.840 1292.670 2240.120 ;
        RECT 1293.510 2239.840 1303.250 2240.120 ;
        RECT 1304.090 2239.840 1314.290 2240.120 ;
        RECT 1315.130 2239.840 1324.870 2240.120 ;
        RECT 1325.710 2239.840 1335.450 2240.120 ;
        RECT 1336.290 2239.840 1346.490 2240.120 ;
        RECT 1347.330 2239.840 1357.070 2240.120 ;
        RECT 1357.910 2239.840 1368.110 2240.120 ;
        RECT 1368.950 2239.840 1378.690 2240.120 ;
        RECT 1379.530 2239.840 1389.270 2240.120 ;
        RECT 1390.110 2239.840 1400.310 2240.120 ;
        RECT 1401.150 2239.840 1410.890 2240.120 ;
        RECT 1411.730 2239.840 1421.930 2240.120 ;
        RECT 1422.770 2239.840 1432.510 2240.120 ;
        RECT 1433.350 2239.840 1443.090 2240.120 ;
        RECT 1443.930 2239.840 1454.130 2240.120 ;
        RECT 1454.970 2239.840 1464.710 2240.120 ;
        RECT 1465.550 2239.840 1475.750 2240.120 ;
        RECT 1476.590 2239.840 1486.330 2240.120 ;
        RECT 1487.170 2239.840 1496.910 2240.120 ;
        RECT 1497.750 2239.840 1507.950 2240.120 ;
        RECT 1508.790 2239.840 1518.530 2240.120 ;
        RECT 1519.370 2239.840 1529.570 2240.120 ;
        RECT 1530.410 2239.840 1540.150 2240.120 ;
        RECT 1540.990 2239.840 1551.190 2240.120 ;
        RECT 1552.030 2239.840 1561.770 2240.120 ;
        RECT 1562.610 2239.840 1572.350 2240.120 ;
        RECT 1573.190 2239.840 1583.390 2240.120 ;
        RECT 1584.230 2239.840 1593.970 2240.120 ;
        RECT 1594.810 2239.840 1605.010 2240.120 ;
        RECT 1605.850 2239.840 1615.590 2240.120 ;
        RECT 1616.430 2239.840 1626.170 2240.120 ;
        RECT 1627.010 2239.840 1637.210 2240.120 ;
        RECT 1638.050 2239.840 1647.790 2240.120 ;
        RECT 1648.630 2239.840 1658.830 2240.120 ;
        RECT 1659.670 2239.840 1669.410 2240.120 ;
        RECT 1670.250 2239.840 1679.990 2240.120 ;
        RECT 1680.830 2239.840 1691.030 2240.120 ;
        RECT 1691.870 2239.840 1701.610 2240.120 ;
        RECT 1702.450 2239.840 1712.650 2240.120 ;
        RECT 1713.490 2239.840 1723.230 2240.120 ;
        RECT 1724.070 2239.840 1734.270 2240.120 ;
        RECT 1735.110 2239.840 1744.850 2240.120 ;
        RECT 1745.690 2239.840 1755.430 2240.120 ;
        RECT 1756.270 2239.840 1766.470 2240.120 ;
        RECT 1767.310 2239.840 1777.050 2240.120 ;
        RECT 1777.890 2239.840 1788.090 2240.120 ;
        RECT 1788.930 2239.840 1798.670 2240.120 ;
        RECT 1799.510 2239.840 1809.250 2240.120 ;
        RECT 1810.090 2239.840 1820.290 2240.120 ;
        RECT 1821.130 2239.840 1830.870 2240.120 ;
        RECT 1831.710 2239.840 1841.910 2240.120 ;
        RECT 1842.750 2239.840 1852.490 2240.120 ;
        RECT 1853.330 2239.840 1863.070 2240.120 ;
        RECT 1863.910 2239.840 1874.110 2240.120 ;
        RECT 1874.950 2239.840 1884.690 2240.120 ;
        RECT 1885.530 2239.840 1895.730 2240.120 ;
        RECT 1896.570 2239.840 1906.310 2240.120 ;
        RECT 1907.150 2239.840 1916.890 2240.120 ;
        RECT 1917.730 2239.840 1927.930 2240.120 ;
        RECT 1928.770 2239.840 1938.510 2240.120 ;
        RECT 1939.350 2239.840 1949.550 2240.120 ;
        RECT 1950.390 2239.840 1960.130 2240.120 ;
        RECT 1960.970 2239.840 1971.170 2240.120 ;
        RECT 1972.010 2239.840 1981.750 2240.120 ;
        RECT 1982.590 2239.840 1992.330 2240.120 ;
        RECT 1993.170 2239.840 2003.370 2240.120 ;
        RECT 2004.210 2239.840 2013.950 2240.120 ;
        RECT 2014.790 2239.840 2024.990 2240.120 ;
        RECT 2025.830 2239.840 2035.570 2240.120 ;
        RECT 2036.410 2239.840 2046.150 2240.120 ;
        RECT 2046.990 2239.840 2057.190 2240.120 ;
        RECT 2058.030 2239.840 2067.770 2240.120 ;
        RECT 2068.610 2239.840 2078.810 2240.120 ;
        RECT 2079.650 2239.840 2089.390 2240.120 ;
        RECT 2090.230 2239.840 2099.970 2240.120 ;
        RECT 2100.810 2239.840 2111.010 2240.120 ;
        RECT 2111.850 2239.840 2121.590 2240.120 ;
        RECT 2122.430 2239.840 2132.630 2240.120 ;
        RECT 2133.470 2239.840 2143.210 2240.120 ;
        RECT 54.700 48.400 2143.770 2239.840 ;
        RECT 55.190 44.955 64.930 48.400 ;
        RECT 65.770 44.955 75.510 48.400 ;
        RECT 76.350 44.955 86.090 48.400 ;
        RECT 86.930 44.955 96.670 48.400 ;
        RECT 97.510 44.955 107.250 48.400 ;
        RECT 108.090 44.955 117.830 48.400 ;
        RECT 118.670 44.955 128.410 48.400 ;
        RECT 129.250 44.955 138.990 48.400 ;
        RECT 139.830 44.955 149.570 48.400 ;
        RECT 150.410 44.955 160.150 48.400 ;
        RECT 160.990 44.955 170.730 48.400 ;
        RECT 171.570 44.955 181.310 48.400 ;
        RECT 182.150 44.955 191.890 48.400 ;
        RECT 192.730 44.955 202.470 48.400 ;
        RECT 203.310 44.955 213.050 48.400 ;
        RECT 213.890 44.955 223.630 48.400 ;
        RECT 224.470 44.955 234.210 48.400 ;
        RECT 235.050 44.955 245.250 48.400 ;
        RECT 246.090 44.955 255.830 48.400 ;
        RECT 256.670 44.955 266.410 48.400 ;
        RECT 267.250 44.955 276.990 48.400 ;
        RECT 277.830 44.955 287.570 48.400 ;
        RECT 288.410 44.955 298.150 48.400 ;
        RECT 298.990 44.955 308.730 48.400 ;
        RECT 309.570 44.955 319.310 48.400 ;
        RECT 320.150 44.955 329.890 48.400 ;
        RECT 330.730 44.955 340.470 48.400 ;
        RECT 341.310 44.955 351.050 48.400 ;
        RECT 351.890 44.955 361.630 48.400 ;
        RECT 362.470 44.955 372.210 48.400 ;
        RECT 373.050 44.955 382.790 48.400 ;
        RECT 383.630 44.955 393.370 48.400 ;
        RECT 394.210 44.955 403.950 48.400 ;
        RECT 404.790 44.955 414.530 48.400 ;
        RECT 415.370 44.955 425.110 48.400 ;
        RECT 425.950 44.955 436.150 48.400 ;
        RECT 436.990 44.955 446.730 48.400 ;
        RECT 447.570 44.955 457.310 48.400 ;
        RECT 458.150 44.955 467.890 48.400 ;
        RECT 468.730 44.955 478.470 48.400 ;
        RECT 479.310 44.955 489.050 48.400 ;
        RECT 489.890 44.955 499.630 48.400 ;
        RECT 500.470 44.955 510.210 48.400 ;
        RECT 511.050 44.955 520.790 48.400 ;
        RECT 521.630 44.955 531.370 48.400 ;
        RECT 532.210 44.955 541.950 48.400 ;
        RECT 542.790 44.955 552.530 48.400 ;
        RECT 553.370 44.955 563.110 48.400 ;
        RECT 563.950 44.955 573.690 48.400 ;
        RECT 574.530 44.955 584.270 48.400 ;
        RECT 585.110 44.955 594.850 48.400 ;
        RECT 595.690 44.955 605.430 48.400 ;
        RECT 606.270 44.955 616.010 48.400 ;
        RECT 616.850 44.955 627.050 48.400 ;
        RECT 627.890 44.955 637.630 48.400 ;
        RECT 638.470 44.955 648.210 48.400 ;
        RECT 649.050 44.955 658.790 48.400 ;
        RECT 659.630 44.955 669.370 48.400 ;
        RECT 670.210 44.955 679.950 48.400 ;
        RECT 680.790 44.955 690.530 48.400 ;
        RECT 691.370 44.955 701.110 48.400 ;
        RECT 701.950 44.955 711.690 48.400 ;
        RECT 712.530 44.955 722.270 48.400 ;
        RECT 723.110 44.955 732.850 48.400 ;
        RECT 733.690 44.955 743.430 48.400 ;
        RECT 744.270 44.955 754.010 48.400 ;
        RECT 754.850 44.955 764.590 48.400 ;
        RECT 765.430 44.955 775.170 48.400 ;
        RECT 776.010 44.955 785.750 48.400 ;
        RECT 786.590 44.955 796.330 48.400 ;
        RECT 797.170 44.955 806.910 48.400 ;
        RECT 807.750 44.955 817.950 48.400 ;
        RECT 818.790 44.955 828.530 48.400 ;
        RECT 829.370 44.955 839.110 48.400 ;
        RECT 839.950 44.955 849.690 48.400 ;
        RECT 850.530 44.955 860.270 48.400 ;
        RECT 861.110 44.955 870.850 48.400 ;
        RECT 871.690 44.955 881.430 48.400 ;
        RECT 882.270 44.955 892.010 48.400 ;
        RECT 892.850 44.955 902.590 48.400 ;
        RECT 903.430 44.955 913.170 48.400 ;
        RECT 914.010 44.955 923.750 48.400 ;
        RECT 924.590 44.955 934.330 48.400 ;
        RECT 935.170 44.955 944.910 48.400 ;
        RECT 945.750 44.955 955.490 48.400 ;
        RECT 956.330 44.955 966.070 48.400 ;
        RECT 966.910 44.955 976.650 48.400 ;
        RECT 977.490 44.955 987.230 48.400 ;
        RECT 988.070 44.955 997.810 48.400 ;
        RECT 998.650 44.955 1008.850 48.400 ;
        RECT 1009.690 44.955 1019.430 48.400 ;
        RECT 1020.270 44.955 1030.010 48.400 ;
        RECT 1030.850 44.955 1040.590 48.400 ;
        RECT 1041.430 44.955 1051.170 48.400 ;
        RECT 1052.010 44.955 1061.750 48.400 ;
        RECT 1062.590 44.955 1072.330 48.400 ;
        RECT 1073.170 44.955 1082.910 48.400 ;
        RECT 1083.750 44.955 1093.490 48.400 ;
        RECT 1094.330 44.955 1104.070 48.400 ;
        RECT 1104.910 44.955 1114.650 48.400 ;
        RECT 1115.490 44.955 1125.230 48.400 ;
        RECT 1126.070 44.955 1135.810 48.400 ;
        RECT 1136.650 44.955 1146.390 48.400 ;
        RECT 1147.230 44.955 1156.970 48.400 ;
        RECT 1157.810 44.955 1167.550 48.400 ;
        RECT 1168.390 44.955 1178.130 48.400 ;
        RECT 1178.970 44.955 1188.710 48.400 ;
        RECT 1189.550 44.955 1199.750 48.400 ;
        RECT 1200.590 44.955 1210.330 48.400 ;
        RECT 1211.170 44.955 1220.910 48.400 ;
        RECT 1221.750 44.955 1231.490 48.400 ;
        RECT 1232.330 44.955 1242.070 48.400 ;
        RECT 1242.910 44.955 1252.650 48.400 ;
        RECT 1253.490 44.955 1263.230 48.400 ;
        RECT 1264.070 44.955 1273.810 48.400 ;
        RECT 1274.650 44.955 1284.390 48.400 ;
        RECT 1285.230 44.955 1294.970 48.400 ;
        RECT 1295.810 44.955 1305.550 48.400 ;
        RECT 1306.390 44.955 1316.130 48.400 ;
        RECT 1316.970 44.955 1326.710 48.400 ;
        RECT 1327.550 44.955 1337.290 48.400 ;
        RECT 1338.130 44.955 1347.870 48.400 ;
        RECT 1348.710 44.955 1358.450 48.400 ;
        RECT 1359.290 44.955 1369.030 48.400 ;
        RECT 1369.870 44.955 1379.610 48.400 ;
        RECT 1380.450 44.955 1390.650 48.400 ;
        RECT 1391.490 44.955 1401.230 48.400 ;
        RECT 1402.070 44.955 1411.810 48.400 ;
        RECT 1412.650 44.955 1422.390 48.400 ;
        RECT 1423.230 44.955 1432.970 48.400 ;
        RECT 1433.810 44.955 1443.550 48.400 ;
        RECT 1444.390 44.955 1454.130 48.400 ;
        RECT 1454.970 44.955 1464.710 48.400 ;
        RECT 1465.550 44.955 1475.290 48.400 ;
        RECT 1476.130 44.955 1485.870 48.400 ;
        RECT 1486.710 44.955 1496.450 48.400 ;
        RECT 1497.290 44.955 1507.030 48.400 ;
        RECT 1507.870 44.955 1517.610 48.400 ;
        RECT 1518.450 44.955 1528.190 48.400 ;
        RECT 1529.030 44.955 1538.770 48.400 ;
        RECT 1539.610 44.955 1549.350 48.400 ;
        RECT 1550.190 44.955 1559.930 48.400 ;
        RECT 1560.770 44.955 1570.510 48.400 ;
        RECT 1571.350 44.955 1581.550 48.400 ;
        RECT 1582.390 44.955 1592.130 48.400 ;
        RECT 1592.970 44.955 1602.710 48.400 ;
        RECT 1603.550 44.955 1613.290 48.400 ;
        RECT 1614.130 44.955 1623.870 48.400 ;
        RECT 1624.710 44.955 1634.450 48.400 ;
        RECT 1635.290 44.955 1645.030 48.400 ;
        RECT 1645.870 44.955 1655.610 48.400 ;
        RECT 1656.450 44.955 1666.190 48.400 ;
        RECT 1667.030 44.955 1676.770 48.400 ;
        RECT 1677.610 44.955 1687.350 48.400 ;
        RECT 1688.190 44.955 1697.930 48.400 ;
        RECT 1698.770 44.955 1708.510 48.400 ;
        RECT 1709.350 44.955 1719.090 48.400 ;
        RECT 1719.930 44.955 1729.670 48.400 ;
        RECT 1730.510 44.955 1740.250 48.400 ;
        RECT 1741.090 44.955 1750.830 48.400 ;
        RECT 1751.670 44.955 1761.410 48.400 ;
        RECT 1762.250 44.955 1772.450 48.400 ;
        RECT 1773.290 44.955 1783.030 48.400 ;
        RECT 1783.870 44.955 1793.610 48.400 ;
        RECT 1794.450 44.955 1804.190 48.400 ;
        RECT 1805.030 44.955 1814.770 48.400 ;
        RECT 1815.610 44.955 1825.350 48.400 ;
        RECT 1826.190 44.955 1835.930 48.400 ;
        RECT 1836.770 44.955 1846.510 48.400 ;
        RECT 1847.350 44.955 1857.090 48.400 ;
        RECT 1857.930 44.955 1867.670 48.400 ;
        RECT 1868.510 44.955 1878.250 48.400 ;
        RECT 1879.090 44.955 1888.830 48.400 ;
        RECT 1889.670 44.955 1899.410 48.400 ;
        RECT 1900.250 44.955 1909.990 48.400 ;
        RECT 1910.830 44.955 1920.570 48.400 ;
        RECT 1921.410 44.955 1931.150 48.400 ;
        RECT 1931.990 44.955 1941.730 48.400 ;
        RECT 1942.570 44.955 1952.310 48.400 ;
        RECT 1953.150 44.955 1963.350 48.400 ;
        RECT 1964.190 44.955 1973.930 48.400 ;
        RECT 1974.770 44.955 1984.510 48.400 ;
        RECT 1985.350 44.955 1995.090 48.400 ;
        RECT 1995.930 44.955 2005.670 48.400 ;
        RECT 2006.510 44.955 2016.250 48.400 ;
        RECT 2017.090 44.955 2026.830 48.400 ;
        RECT 2027.670 44.955 2037.410 48.400 ;
        RECT 2038.250 44.955 2047.990 48.400 ;
        RECT 2048.830 44.955 2058.570 48.400 ;
        RECT 2059.410 44.955 2069.150 48.400 ;
        RECT 2069.990 44.955 2079.730 48.400 ;
        RECT 2080.570 44.955 2090.310 48.400 ;
        RECT 2091.150 44.955 2100.890 48.400 ;
        RECT 2101.730 44.955 2111.470 48.400 ;
        RECT 2112.310 44.955 2122.050 48.400 ;
        RECT 2122.890 44.955 2132.630 48.400 ;
        RECT 2133.470 44.955 2143.210 48.400 ;
      LAYER met3 ;
        RECT 53.880 2237.440 2145.080 2238.305 ;
        RECT 53.470 2227.280 2145.480 2237.440 ;
        RECT 53.880 2225.880 2145.080 2227.280 ;
        RECT 53.470 2216.400 2145.480 2225.880 ;
        RECT 53.880 2215.000 2145.080 2216.400 ;
        RECT 53.470 2204.840 2145.480 2215.000 ;
        RECT 53.880 2203.440 2145.080 2204.840 ;
        RECT 53.470 2193.960 2145.480 2203.440 ;
        RECT 53.880 2192.560 2145.080 2193.960 ;
        RECT 53.470 2182.400 2145.480 2192.560 ;
        RECT 53.880 2181.000 2145.080 2182.400 ;
        RECT 53.470 2171.520 2145.480 2181.000 ;
        RECT 53.880 2170.840 2145.480 2171.520 ;
        RECT 53.880 2170.120 2145.080 2170.840 ;
        RECT 53.470 2169.440 2145.080 2170.120 ;
        RECT 53.470 2159.960 2145.480 2169.440 ;
        RECT 53.880 2158.560 2145.080 2159.960 ;
        RECT 53.470 2149.080 2145.480 2158.560 ;
        RECT 53.880 2148.400 2145.480 2149.080 ;
        RECT 53.880 2147.680 2145.080 2148.400 ;
        RECT 53.470 2147.000 2145.080 2147.680 ;
        RECT 53.470 2137.520 2145.480 2147.000 ;
        RECT 53.880 2136.120 2145.080 2137.520 ;
        RECT 53.470 2126.640 2145.480 2136.120 ;
        RECT 53.880 2125.960 2145.480 2126.640 ;
        RECT 53.880 2125.240 2145.080 2125.960 ;
        RECT 53.470 2124.560 2145.080 2125.240 ;
        RECT 53.470 2115.080 2145.480 2124.560 ;
        RECT 53.880 2114.400 2145.480 2115.080 ;
        RECT 53.880 2113.680 2145.080 2114.400 ;
        RECT 53.470 2113.000 2145.080 2113.680 ;
        RECT 53.470 2104.200 2145.480 2113.000 ;
        RECT 53.880 2103.520 2145.480 2104.200 ;
        RECT 53.880 2102.800 2145.080 2103.520 ;
        RECT 53.470 2102.120 2145.080 2102.800 ;
        RECT 53.470 2092.640 2145.480 2102.120 ;
        RECT 53.880 2091.960 2145.480 2092.640 ;
        RECT 53.880 2091.240 2145.080 2091.960 ;
        RECT 53.470 2090.560 2145.080 2091.240 ;
        RECT 53.470 2081.760 2145.480 2090.560 ;
        RECT 53.880 2081.080 2145.480 2081.760 ;
        RECT 53.880 2080.360 2145.080 2081.080 ;
        RECT 53.470 2079.680 2145.080 2080.360 ;
        RECT 53.470 2070.200 2145.480 2079.680 ;
        RECT 53.880 2069.520 2145.480 2070.200 ;
        RECT 53.880 2068.800 2145.080 2069.520 ;
        RECT 53.470 2068.120 2145.080 2068.800 ;
        RECT 53.470 2059.320 2145.480 2068.120 ;
        RECT 53.880 2057.960 2145.480 2059.320 ;
        RECT 53.880 2057.920 2145.080 2057.960 ;
        RECT 53.470 2056.560 2145.080 2057.920 ;
        RECT 53.470 2047.760 2145.480 2056.560 ;
        RECT 53.880 2047.080 2145.480 2047.760 ;
        RECT 53.880 2046.360 2145.080 2047.080 ;
        RECT 53.470 2045.680 2145.080 2046.360 ;
        RECT 53.470 2036.880 2145.480 2045.680 ;
        RECT 53.880 2035.520 2145.480 2036.880 ;
        RECT 53.880 2035.480 2145.080 2035.520 ;
        RECT 53.470 2034.120 2145.080 2035.480 ;
        RECT 53.470 2025.320 2145.480 2034.120 ;
        RECT 53.880 2024.640 2145.480 2025.320 ;
        RECT 53.880 2023.920 2145.080 2024.640 ;
        RECT 53.470 2023.240 2145.080 2023.920 ;
        RECT 53.470 2014.440 2145.480 2023.240 ;
        RECT 53.880 2013.080 2145.480 2014.440 ;
        RECT 53.880 2013.040 2145.080 2013.080 ;
        RECT 53.470 2011.680 2145.080 2013.040 ;
        RECT 53.470 2002.880 2145.480 2011.680 ;
        RECT 53.880 2002.200 2145.480 2002.880 ;
        RECT 53.880 2001.480 2145.080 2002.200 ;
        RECT 53.470 2000.800 2145.080 2001.480 ;
        RECT 53.470 1992.000 2145.480 2000.800 ;
        RECT 53.880 1990.640 2145.480 1992.000 ;
        RECT 53.880 1990.600 2145.080 1990.640 ;
        RECT 53.470 1989.240 2145.080 1990.600 ;
        RECT 53.470 1980.440 2145.480 1989.240 ;
        RECT 53.880 1979.080 2145.480 1980.440 ;
        RECT 53.880 1979.040 2145.080 1979.080 ;
        RECT 53.470 1977.680 2145.080 1979.040 ;
        RECT 53.470 1969.560 2145.480 1977.680 ;
        RECT 53.880 1968.200 2145.480 1969.560 ;
        RECT 53.880 1968.160 2145.080 1968.200 ;
        RECT 53.470 1966.800 2145.080 1968.160 ;
        RECT 53.470 1958.000 2145.480 1966.800 ;
        RECT 53.880 1956.640 2145.480 1958.000 ;
        RECT 53.880 1956.600 2145.080 1956.640 ;
        RECT 53.470 1955.240 2145.080 1956.600 ;
        RECT 53.470 1947.120 2145.480 1955.240 ;
        RECT 53.880 1945.760 2145.480 1947.120 ;
        RECT 53.880 1945.720 2145.080 1945.760 ;
        RECT 53.470 1944.360 2145.080 1945.720 ;
        RECT 53.470 1935.560 2145.480 1944.360 ;
        RECT 53.880 1934.200 2145.480 1935.560 ;
        RECT 53.880 1934.160 2145.080 1934.200 ;
        RECT 53.470 1932.800 2145.080 1934.160 ;
        RECT 53.470 1924.680 2145.480 1932.800 ;
        RECT 53.880 1923.280 2145.480 1924.680 ;
        RECT 53.470 1922.640 2145.480 1923.280 ;
        RECT 53.470 1921.240 2145.080 1922.640 ;
        RECT 53.470 1913.120 2145.480 1921.240 ;
        RECT 53.880 1911.760 2145.480 1913.120 ;
        RECT 53.880 1911.720 2145.080 1911.760 ;
        RECT 53.470 1910.360 2145.080 1911.720 ;
        RECT 53.470 1902.240 2145.480 1910.360 ;
        RECT 53.880 1900.840 2145.480 1902.240 ;
        RECT 53.470 1900.200 2145.480 1900.840 ;
        RECT 53.470 1898.800 2145.080 1900.200 ;
        RECT 53.470 1890.680 2145.480 1898.800 ;
        RECT 53.880 1889.320 2145.480 1890.680 ;
        RECT 53.880 1889.280 2145.080 1889.320 ;
        RECT 53.470 1887.920 2145.080 1889.280 ;
        RECT 53.470 1879.800 2145.480 1887.920 ;
        RECT 53.880 1878.400 2145.480 1879.800 ;
        RECT 53.470 1877.760 2145.480 1878.400 ;
        RECT 53.470 1876.360 2145.080 1877.760 ;
        RECT 53.470 1868.240 2145.480 1876.360 ;
        RECT 53.880 1866.840 2145.480 1868.240 ;
        RECT 53.470 1866.200 2145.480 1866.840 ;
        RECT 53.470 1864.800 2145.080 1866.200 ;
        RECT 53.470 1857.360 2145.480 1864.800 ;
        RECT 53.880 1855.960 2145.480 1857.360 ;
        RECT 53.470 1855.320 2145.480 1855.960 ;
        RECT 53.470 1853.920 2145.080 1855.320 ;
        RECT 53.470 1845.800 2145.480 1853.920 ;
        RECT 53.880 1844.400 2145.480 1845.800 ;
        RECT 53.470 1843.760 2145.480 1844.400 ;
        RECT 53.470 1842.360 2145.080 1843.760 ;
        RECT 53.470 1834.920 2145.480 1842.360 ;
        RECT 53.880 1833.520 2145.480 1834.920 ;
        RECT 53.470 1832.880 2145.480 1833.520 ;
        RECT 53.470 1831.480 2145.080 1832.880 ;
        RECT 53.470 1823.360 2145.480 1831.480 ;
        RECT 53.880 1821.960 2145.480 1823.360 ;
        RECT 53.470 1821.320 2145.480 1821.960 ;
        RECT 53.470 1819.920 2145.080 1821.320 ;
        RECT 53.470 1812.480 2145.480 1819.920 ;
        RECT 53.880 1811.080 2145.480 1812.480 ;
        RECT 53.470 1810.440 2145.480 1811.080 ;
        RECT 53.470 1809.040 2145.080 1810.440 ;
        RECT 53.470 1800.920 2145.480 1809.040 ;
        RECT 53.880 1799.520 2145.480 1800.920 ;
        RECT 53.470 1798.880 2145.480 1799.520 ;
        RECT 53.470 1797.480 2145.080 1798.880 ;
        RECT 53.470 1790.040 2145.480 1797.480 ;
        RECT 53.880 1788.640 2145.480 1790.040 ;
        RECT 53.470 1787.320 2145.480 1788.640 ;
        RECT 53.470 1785.920 2145.080 1787.320 ;
        RECT 53.470 1778.480 2145.480 1785.920 ;
        RECT 53.880 1777.080 2145.480 1778.480 ;
        RECT 53.470 1776.440 2145.480 1777.080 ;
        RECT 53.470 1775.040 2145.080 1776.440 ;
        RECT 53.470 1767.600 2145.480 1775.040 ;
        RECT 53.880 1766.200 2145.480 1767.600 ;
        RECT 53.470 1764.880 2145.480 1766.200 ;
        RECT 53.470 1763.480 2145.080 1764.880 ;
        RECT 53.470 1756.040 2145.480 1763.480 ;
        RECT 53.880 1754.640 2145.480 1756.040 ;
        RECT 53.470 1754.000 2145.480 1754.640 ;
        RECT 53.470 1752.600 2145.080 1754.000 ;
        RECT 53.470 1745.160 2145.480 1752.600 ;
        RECT 53.880 1743.760 2145.480 1745.160 ;
        RECT 53.470 1742.440 2145.480 1743.760 ;
        RECT 53.470 1741.040 2145.080 1742.440 ;
        RECT 53.470 1733.600 2145.480 1741.040 ;
        RECT 53.880 1732.200 2145.480 1733.600 ;
        RECT 53.470 1730.880 2145.480 1732.200 ;
        RECT 53.470 1729.480 2145.080 1730.880 ;
        RECT 53.470 1722.720 2145.480 1729.480 ;
        RECT 53.880 1721.320 2145.480 1722.720 ;
        RECT 53.470 1720.000 2145.480 1721.320 ;
        RECT 53.470 1718.600 2145.080 1720.000 ;
        RECT 53.470 1711.160 2145.480 1718.600 ;
        RECT 53.880 1709.760 2145.480 1711.160 ;
        RECT 53.470 1708.440 2145.480 1709.760 ;
        RECT 53.470 1707.040 2145.080 1708.440 ;
        RECT 53.470 1700.280 2145.480 1707.040 ;
        RECT 53.880 1698.880 2145.480 1700.280 ;
        RECT 53.470 1697.560 2145.480 1698.880 ;
        RECT 53.470 1696.160 2145.080 1697.560 ;
        RECT 53.470 1688.720 2145.480 1696.160 ;
        RECT 53.880 1687.320 2145.480 1688.720 ;
        RECT 53.470 1686.000 2145.480 1687.320 ;
        RECT 53.470 1684.600 2145.080 1686.000 ;
        RECT 53.470 1677.840 2145.480 1684.600 ;
        RECT 53.880 1676.440 2145.480 1677.840 ;
        RECT 53.470 1674.440 2145.480 1676.440 ;
        RECT 53.470 1673.040 2145.080 1674.440 ;
        RECT 53.470 1666.280 2145.480 1673.040 ;
        RECT 53.880 1664.880 2145.480 1666.280 ;
        RECT 53.470 1663.560 2145.480 1664.880 ;
        RECT 53.470 1662.160 2145.080 1663.560 ;
        RECT 53.470 1655.400 2145.480 1662.160 ;
        RECT 53.880 1654.000 2145.480 1655.400 ;
        RECT 53.470 1652.000 2145.480 1654.000 ;
        RECT 53.470 1650.600 2145.080 1652.000 ;
        RECT 53.470 1643.840 2145.480 1650.600 ;
        RECT 53.880 1642.440 2145.480 1643.840 ;
        RECT 53.470 1641.120 2145.480 1642.440 ;
        RECT 53.470 1639.720 2145.080 1641.120 ;
        RECT 53.470 1632.960 2145.480 1639.720 ;
        RECT 53.880 1631.560 2145.480 1632.960 ;
        RECT 53.470 1629.560 2145.480 1631.560 ;
        RECT 53.470 1628.160 2145.080 1629.560 ;
        RECT 53.470 1621.400 2145.480 1628.160 ;
        RECT 53.880 1620.000 2145.480 1621.400 ;
        RECT 53.470 1618.000 2145.480 1620.000 ;
        RECT 53.470 1616.600 2145.080 1618.000 ;
        RECT 53.470 1610.520 2145.480 1616.600 ;
        RECT 53.880 1609.120 2145.480 1610.520 ;
        RECT 53.470 1607.120 2145.480 1609.120 ;
        RECT 53.470 1605.720 2145.080 1607.120 ;
        RECT 53.470 1598.960 2145.480 1605.720 ;
        RECT 53.880 1597.560 2145.480 1598.960 ;
        RECT 53.470 1595.560 2145.480 1597.560 ;
        RECT 53.470 1594.160 2145.080 1595.560 ;
        RECT 53.470 1588.080 2145.480 1594.160 ;
        RECT 53.880 1586.680 2145.480 1588.080 ;
        RECT 53.470 1584.680 2145.480 1586.680 ;
        RECT 53.470 1583.280 2145.080 1584.680 ;
        RECT 53.470 1576.520 2145.480 1583.280 ;
        RECT 53.880 1575.120 2145.480 1576.520 ;
        RECT 53.470 1573.120 2145.480 1575.120 ;
        RECT 53.470 1571.720 2145.080 1573.120 ;
        RECT 53.470 1565.640 2145.480 1571.720 ;
        RECT 53.880 1564.240 2145.480 1565.640 ;
        RECT 53.470 1562.240 2145.480 1564.240 ;
        RECT 53.470 1560.840 2145.080 1562.240 ;
        RECT 53.470 1554.080 2145.480 1560.840 ;
        RECT 53.880 1552.680 2145.480 1554.080 ;
        RECT 53.470 1550.680 2145.480 1552.680 ;
        RECT 53.470 1549.280 2145.080 1550.680 ;
        RECT 53.470 1543.200 2145.480 1549.280 ;
        RECT 53.880 1541.800 2145.480 1543.200 ;
        RECT 53.470 1539.120 2145.480 1541.800 ;
        RECT 53.470 1537.720 2145.080 1539.120 ;
        RECT 53.470 1531.640 2145.480 1537.720 ;
        RECT 53.880 1530.240 2145.480 1531.640 ;
        RECT 53.470 1528.240 2145.480 1530.240 ;
        RECT 53.470 1526.840 2145.080 1528.240 ;
        RECT 53.470 1520.760 2145.480 1526.840 ;
        RECT 53.880 1519.360 2145.480 1520.760 ;
        RECT 53.470 1516.680 2145.480 1519.360 ;
        RECT 53.470 1515.280 2145.080 1516.680 ;
        RECT 53.470 1509.200 2145.480 1515.280 ;
        RECT 53.880 1507.800 2145.480 1509.200 ;
        RECT 53.470 1505.800 2145.480 1507.800 ;
        RECT 53.470 1504.400 2145.080 1505.800 ;
        RECT 53.470 1498.320 2145.480 1504.400 ;
        RECT 53.880 1496.920 2145.480 1498.320 ;
        RECT 53.470 1494.240 2145.480 1496.920 ;
        RECT 53.470 1492.840 2145.080 1494.240 ;
        RECT 53.470 1486.760 2145.480 1492.840 ;
        RECT 53.880 1485.360 2145.480 1486.760 ;
        RECT 53.470 1482.680 2145.480 1485.360 ;
        RECT 53.470 1481.280 2145.080 1482.680 ;
        RECT 53.470 1475.880 2145.480 1481.280 ;
        RECT 53.880 1474.480 2145.480 1475.880 ;
        RECT 53.470 1471.800 2145.480 1474.480 ;
        RECT 53.470 1470.400 2145.080 1471.800 ;
        RECT 53.470 1464.320 2145.480 1470.400 ;
        RECT 53.880 1462.920 2145.480 1464.320 ;
        RECT 53.470 1460.240 2145.480 1462.920 ;
        RECT 53.470 1458.840 2145.080 1460.240 ;
        RECT 53.470 1453.440 2145.480 1458.840 ;
        RECT 53.880 1452.040 2145.480 1453.440 ;
        RECT 53.470 1449.360 2145.480 1452.040 ;
        RECT 53.470 1447.960 2145.080 1449.360 ;
        RECT 53.470 1441.880 2145.480 1447.960 ;
        RECT 53.880 1440.480 2145.480 1441.880 ;
        RECT 53.470 1437.800 2145.480 1440.480 ;
        RECT 53.470 1436.400 2145.080 1437.800 ;
        RECT 53.470 1431.000 2145.480 1436.400 ;
        RECT 53.880 1429.600 2145.480 1431.000 ;
        RECT 53.470 1426.240 2145.480 1429.600 ;
        RECT 53.470 1424.840 2145.080 1426.240 ;
        RECT 53.470 1419.440 2145.480 1424.840 ;
        RECT 53.880 1418.040 2145.480 1419.440 ;
        RECT 53.470 1415.360 2145.480 1418.040 ;
        RECT 53.470 1413.960 2145.080 1415.360 ;
        RECT 53.470 1408.560 2145.480 1413.960 ;
        RECT 53.880 1407.160 2145.480 1408.560 ;
        RECT 53.470 1403.800 2145.480 1407.160 ;
        RECT 53.470 1402.400 2145.080 1403.800 ;
        RECT 53.470 1397.000 2145.480 1402.400 ;
        RECT 53.880 1395.600 2145.480 1397.000 ;
        RECT 53.470 1392.920 2145.480 1395.600 ;
        RECT 53.470 1391.520 2145.080 1392.920 ;
        RECT 53.470 1386.120 2145.480 1391.520 ;
        RECT 53.880 1384.720 2145.480 1386.120 ;
        RECT 53.470 1381.360 2145.480 1384.720 ;
        RECT 53.470 1379.960 2145.080 1381.360 ;
        RECT 53.470 1374.560 2145.480 1379.960 ;
        RECT 53.880 1373.160 2145.480 1374.560 ;
        RECT 53.470 1370.480 2145.480 1373.160 ;
        RECT 53.470 1369.080 2145.080 1370.480 ;
        RECT 53.470 1363.680 2145.480 1369.080 ;
        RECT 53.880 1362.280 2145.480 1363.680 ;
        RECT 53.470 1358.920 2145.480 1362.280 ;
        RECT 53.470 1357.520 2145.080 1358.920 ;
        RECT 53.470 1352.120 2145.480 1357.520 ;
        RECT 53.880 1350.720 2145.480 1352.120 ;
        RECT 53.470 1347.360 2145.480 1350.720 ;
        RECT 53.470 1345.960 2145.080 1347.360 ;
        RECT 53.470 1341.240 2145.480 1345.960 ;
        RECT 53.880 1339.840 2145.480 1341.240 ;
        RECT 53.470 1336.480 2145.480 1339.840 ;
        RECT 53.470 1335.080 2145.080 1336.480 ;
        RECT 53.470 1329.680 2145.480 1335.080 ;
        RECT 53.880 1328.280 2145.480 1329.680 ;
        RECT 53.470 1324.920 2145.480 1328.280 ;
        RECT 53.470 1323.520 2145.080 1324.920 ;
        RECT 53.470 1318.800 2145.480 1323.520 ;
        RECT 53.880 1317.400 2145.480 1318.800 ;
        RECT 53.470 1314.040 2145.480 1317.400 ;
        RECT 53.470 1312.640 2145.080 1314.040 ;
        RECT 53.470 1307.240 2145.480 1312.640 ;
        RECT 53.880 1305.840 2145.480 1307.240 ;
        RECT 53.470 1302.480 2145.480 1305.840 ;
        RECT 53.470 1301.080 2145.080 1302.480 ;
        RECT 53.470 1296.360 2145.480 1301.080 ;
        RECT 53.880 1294.960 2145.480 1296.360 ;
        RECT 53.470 1290.920 2145.480 1294.960 ;
        RECT 53.470 1289.520 2145.080 1290.920 ;
        RECT 53.470 1284.800 2145.480 1289.520 ;
        RECT 53.880 1283.400 2145.480 1284.800 ;
        RECT 53.470 1280.040 2145.480 1283.400 ;
        RECT 53.470 1278.640 2145.080 1280.040 ;
        RECT 53.470 1273.920 2145.480 1278.640 ;
        RECT 53.880 1272.520 2145.480 1273.920 ;
        RECT 53.470 1268.480 2145.480 1272.520 ;
        RECT 53.470 1267.080 2145.080 1268.480 ;
        RECT 53.470 1262.360 2145.480 1267.080 ;
        RECT 53.880 1260.960 2145.480 1262.360 ;
        RECT 53.470 1257.600 2145.480 1260.960 ;
        RECT 53.470 1256.200 2145.080 1257.600 ;
        RECT 53.470 1251.480 2145.480 1256.200 ;
        RECT 53.880 1250.080 2145.480 1251.480 ;
        RECT 53.470 1246.040 2145.480 1250.080 ;
        RECT 53.470 1244.640 2145.080 1246.040 ;
        RECT 53.470 1239.920 2145.480 1244.640 ;
        RECT 53.880 1238.520 2145.480 1239.920 ;
        RECT 53.470 1234.480 2145.480 1238.520 ;
        RECT 53.470 1233.080 2145.080 1234.480 ;
        RECT 53.470 1229.040 2145.480 1233.080 ;
        RECT 53.880 1227.640 2145.480 1229.040 ;
        RECT 53.470 1223.600 2145.480 1227.640 ;
        RECT 53.470 1222.200 2145.080 1223.600 ;
        RECT 53.470 1217.480 2145.480 1222.200 ;
        RECT 53.880 1216.080 2145.480 1217.480 ;
        RECT 53.470 1212.040 2145.480 1216.080 ;
        RECT 53.470 1210.640 2145.080 1212.040 ;
        RECT 53.470 1206.600 2145.480 1210.640 ;
        RECT 53.880 1205.200 2145.480 1206.600 ;
        RECT 53.470 1201.160 2145.480 1205.200 ;
        RECT 53.470 1199.760 2145.080 1201.160 ;
        RECT 53.470 1195.040 2145.480 1199.760 ;
        RECT 53.880 1193.640 2145.480 1195.040 ;
        RECT 53.470 1189.600 2145.480 1193.640 ;
        RECT 53.470 1188.200 2145.080 1189.600 ;
        RECT 53.470 1184.160 2145.480 1188.200 ;
        RECT 53.880 1182.760 2145.480 1184.160 ;
        RECT 53.470 1178.040 2145.480 1182.760 ;
        RECT 53.470 1176.640 2145.080 1178.040 ;
        RECT 53.470 1172.600 2145.480 1176.640 ;
        RECT 53.880 1171.200 2145.480 1172.600 ;
        RECT 53.470 1167.160 2145.480 1171.200 ;
        RECT 53.470 1165.760 2145.080 1167.160 ;
        RECT 53.470 1161.720 2145.480 1165.760 ;
        RECT 53.880 1160.320 2145.480 1161.720 ;
        RECT 53.470 1155.600 2145.480 1160.320 ;
        RECT 53.470 1154.200 2145.080 1155.600 ;
        RECT 53.470 1150.160 2145.480 1154.200 ;
        RECT 53.880 1148.760 2145.480 1150.160 ;
        RECT 53.470 1144.720 2145.480 1148.760 ;
        RECT 53.470 1143.320 2145.080 1144.720 ;
        RECT 53.470 1138.600 2145.480 1143.320 ;
        RECT 53.880 1137.200 2145.480 1138.600 ;
        RECT 53.470 1133.160 2145.480 1137.200 ;
        RECT 53.470 1131.760 2145.080 1133.160 ;
        RECT 53.470 1127.720 2145.480 1131.760 ;
        RECT 53.880 1126.320 2145.480 1127.720 ;
        RECT 53.470 1122.280 2145.480 1126.320 ;
        RECT 53.470 1120.880 2145.080 1122.280 ;
        RECT 53.470 1116.160 2145.480 1120.880 ;
        RECT 53.880 1114.760 2145.480 1116.160 ;
        RECT 53.470 1110.720 2145.480 1114.760 ;
        RECT 53.470 1109.320 2145.080 1110.720 ;
        RECT 53.470 1105.280 2145.480 1109.320 ;
        RECT 53.880 1103.880 2145.480 1105.280 ;
        RECT 53.470 1099.160 2145.480 1103.880 ;
        RECT 53.470 1097.760 2145.080 1099.160 ;
        RECT 53.470 1093.720 2145.480 1097.760 ;
        RECT 53.880 1092.320 2145.480 1093.720 ;
        RECT 53.470 1088.280 2145.480 1092.320 ;
        RECT 53.470 1086.880 2145.080 1088.280 ;
        RECT 53.470 1082.840 2145.480 1086.880 ;
        RECT 53.880 1081.440 2145.480 1082.840 ;
        RECT 53.470 1076.720 2145.480 1081.440 ;
        RECT 53.470 1075.320 2145.080 1076.720 ;
        RECT 53.470 1071.280 2145.480 1075.320 ;
        RECT 53.880 1069.880 2145.480 1071.280 ;
        RECT 53.470 1065.840 2145.480 1069.880 ;
        RECT 53.470 1064.440 2145.080 1065.840 ;
        RECT 53.470 1060.400 2145.480 1064.440 ;
        RECT 53.880 1059.000 2145.480 1060.400 ;
        RECT 53.470 1054.280 2145.480 1059.000 ;
        RECT 53.470 1052.880 2145.080 1054.280 ;
        RECT 53.470 1048.840 2145.480 1052.880 ;
        RECT 53.880 1047.440 2145.480 1048.840 ;
        RECT 53.470 1042.720 2145.480 1047.440 ;
        RECT 53.470 1041.320 2145.080 1042.720 ;
        RECT 53.470 1037.960 2145.480 1041.320 ;
        RECT 53.880 1036.560 2145.480 1037.960 ;
        RECT 53.470 1031.840 2145.480 1036.560 ;
        RECT 53.470 1030.440 2145.080 1031.840 ;
        RECT 53.470 1026.400 2145.480 1030.440 ;
        RECT 53.880 1025.000 2145.480 1026.400 ;
        RECT 53.470 1020.280 2145.480 1025.000 ;
        RECT 53.470 1018.880 2145.080 1020.280 ;
        RECT 53.470 1015.520 2145.480 1018.880 ;
        RECT 53.880 1014.120 2145.480 1015.520 ;
        RECT 53.470 1009.400 2145.480 1014.120 ;
        RECT 53.470 1008.000 2145.080 1009.400 ;
        RECT 53.470 1003.960 2145.480 1008.000 ;
        RECT 53.880 1002.560 2145.480 1003.960 ;
        RECT 53.470 997.840 2145.480 1002.560 ;
        RECT 53.470 996.440 2145.080 997.840 ;
        RECT 53.470 993.080 2145.480 996.440 ;
        RECT 53.880 991.680 2145.480 993.080 ;
        RECT 53.470 986.280 2145.480 991.680 ;
        RECT 53.470 984.880 2145.080 986.280 ;
        RECT 53.470 981.520 2145.480 984.880 ;
        RECT 53.880 980.120 2145.480 981.520 ;
        RECT 53.470 975.400 2145.480 980.120 ;
        RECT 53.470 974.000 2145.080 975.400 ;
        RECT 53.470 970.640 2145.480 974.000 ;
        RECT 53.880 969.240 2145.480 970.640 ;
        RECT 53.470 963.840 2145.480 969.240 ;
        RECT 53.470 962.440 2145.080 963.840 ;
        RECT 53.470 959.080 2145.480 962.440 ;
        RECT 53.880 957.680 2145.480 959.080 ;
        RECT 53.470 952.960 2145.480 957.680 ;
        RECT 53.470 951.560 2145.080 952.960 ;
        RECT 53.470 948.200 2145.480 951.560 ;
        RECT 53.880 946.800 2145.480 948.200 ;
        RECT 53.470 941.400 2145.480 946.800 ;
        RECT 53.470 940.000 2145.080 941.400 ;
        RECT 53.470 936.640 2145.480 940.000 ;
        RECT 53.880 935.240 2145.480 936.640 ;
        RECT 53.470 930.520 2145.480 935.240 ;
        RECT 53.470 929.120 2145.080 930.520 ;
        RECT 53.470 925.760 2145.480 929.120 ;
        RECT 53.880 924.360 2145.480 925.760 ;
        RECT 53.470 918.960 2145.480 924.360 ;
        RECT 53.470 917.560 2145.080 918.960 ;
        RECT 53.470 914.200 2145.480 917.560 ;
        RECT 53.880 912.800 2145.480 914.200 ;
        RECT 53.470 907.400 2145.480 912.800 ;
        RECT 53.470 906.000 2145.080 907.400 ;
        RECT 53.470 903.320 2145.480 906.000 ;
        RECT 53.880 901.920 2145.480 903.320 ;
        RECT 53.470 896.520 2145.480 901.920 ;
        RECT 53.470 895.120 2145.080 896.520 ;
        RECT 53.470 891.760 2145.480 895.120 ;
        RECT 53.880 890.360 2145.480 891.760 ;
        RECT 53.470 884.960 2145.480 890.360 ;
        RECT 53.470 883.560 2145.080 884.960 ;
        RECT 53.470 880.880 2145.480 883.560 ;
        RECT 53.880 879.480 2145.480 880.880 ;
        RECT 53.470 874.080 2145.480 879.480 ;
        RECT 53.470 872.680 2145.080 874.080 ;
        RECT 53.470 869.320 2145.480 872.680 ;
        RECT 53.880 867.920 2145.480 869.320 ;
        RECT 53.470 862.520 2145.480 867.920 ;
        RECT 53.470 861.120 2145.080 862.520 ;
        RECT 53.470 858.440 2145.480 861.120 ;
        RECT 53.880 857.040 2145.480 858.440 ;
        RECT 53.470 850.960 2145.480 857.040 ;
        RECT 53.470 849.560 2145.080 850.960 ;
        RECT 53.470 846.880 2145.480 849.560 ;
        RECT 53.880 845.480 2145.480 846.880 ;
        RECT 53.470 840.080 2145.480 845.480 ;
        RECT 53.470 838.680 2145.080 840.080 ;
        RECT 53.470 836.000 2145.480 838.680 ;
        RECT 53.880 834.600 2145.480 836.000 ;
        RECT 53.470 828.520 2145.480 834.600 ;
        RECT 53.470 827.120 2145.080 828.520 ;
        RECT 53.470 824.440 2145.480 827.120 ;
        RECT 53.880 823.040 2145.480 824.440 ;
        RECT 53.470 817.640 2145.480 823.040 ;
        RECT 53.470 816.240 2145.080 817.640 ;
        RECT 53.470 813.560 2145.480 816.240 ;
        RECT 53.880 812.160 2145.480 813.560 ;
        RECT 53.470 806.080 2145.480 812.160 ;
        RECT 53.470 804.680 2145.080 806.080 ;
        RECT 53.470 802.000 2145.480 804.680 ;
        RECT 53.880 800.600 2145.480 802.000 ;
        RECT 53.470 794.520 2145.480 800.600 ;
        RECT 53.470 793.120 2145.080 794.520 ;
        RECT 53.470 791.120 2145.480 793.120 ;
        RECT 53.880 789.720 2145.480 791.120 ;
        RECT 53.470 783.640 2145.480 789.720 ;
        RECT 53.470 782.240 2145.080 783.640 ;
        RECT 53.470 779.560 2145.480 782.240 ;
        RECT 53.880 778.160 2145.480 779.560 ;
        RECT 53.470 772.080 2145.480 778.160 ;
        RECT 53.470 770.680 2145.080 772.080 ;
        RECT 53.470 768.680 2145.480 770.680 ;
        RECT 53.880 767.280 2145.480 768.680 ;
        RECT 53.470 761.200 2145.480 767.280 ;
        RECT 53.470 759.800 2145.080 761.200 ;
        RECT 53.470 757.120 2145.480 759.800 ;
        RECT 53.880 755.720 2145.480 757.120 ;
        RECT 53.470 749.640 2145.480 755.720 ;
        RECT 53.470 748.240 2145.080 749.640 ;
        RECT 53.470 746.240 2145.480 748.240 ;
        RECT 53.880 744.840 2145.480 746.240 ;
        RECT 53.470 738.080 2145.480 744.840 ;
        RECT 53.470 736.680 2145.080 738.080 ;
        RECT 53.470 734.680 2145.480 736.680 ;
        RECT 53.880 733.280 2145.480 734.680 ;
        RECT 53.470 727.200 2145.480 733.280 ;
        RECT 53.470 725.800 2145.080 727.200 ;
        RECT 53.470 723.800 2145.480 725.800 ;
        RECT 53.880 722.400 2145.480 723.800 ;
        RECT 53.470 715.640 2145.480 722.400 ;
        RECT 53.470 714.240 2145.080 715.640 ;
        RECT 53.470 712.240 2145.480 714.240 ;
        RECT 53.880 710.840 2145.480 712.240 ;
        RECT 53.470 704.760 2145.480 710.840 ;
        RECT 53.470 703.360 2145.080 704.760 ;
        RECT 53.470 701.360 2145.480 703.360 ;
        RECT 53.880 699.960 2145.480 701.360 ;
        RECT 53.470 693.200 2145.480 699.960 ;
        RECT 53.470 691.800 2145.080 693.200 ;
        RECT 53.470 689.800 2145.480 691.800 ;
        RECT 53.880 688.400 2145.480 689.800 ;
        RECT 53.470 682.320 2145.480 688.400 ;
        RECT 53.470 680.920 2145.080 682.320 ;
        RECT 53.470 678.920 2145.480 680.920 ;
        RECT 53.880 677.520 2145.480 678.920 ;
        RECT 53.470 670.760 2145.480 677.520 ;
        RECT 53.470 669.360 2145.080 670.760 ;
        RECT 53.470 667.360 2145.480 669.360 ;
        RECT 53.880 665.960 2145.480 667.360 ;
        RECT 53.470 659.200 2145.480 665.960 ;
        RECT 53.470 657.800 2145.080 659.200 ;
        RECT 53.470 656.480 2145.480 657.800 ;
        RECT 53.880 655.080 2145.480 656.480 ;
        RECT 53.470 648.320 2145.480 655.080 ;
        RECT 53.470 646.920 2145.080 648.320 ;
        RECT 53.470 644.920 2145.480 646.920 ;
        RECT 53.880 643.520 2145.480 644.920 ;
        RECT 53.470 636.760 2145.480 643.520 ;
        RECT 53.470 635.360 2145.080 636.760 ;
        RECT 53.470 634.040 2145.480 635.360 ;
        RECT 53.880 632.640 2145.480 634.040 ;
        RECT 53.470 625.880 2145.480 632.640 ;
        RECT 53.470 624.480 2145.080 625.880 ;
        RECT 53.470 622.480 2145.480 624.480 ;
        RECT 53.880 621.080 2145.480 622.480 ;
        RECT 53.470 614.320 2145.480 621.080 ;
        RECT 53.470 612.920 2145.080 614.320 ;
        RECT 53.470 611.600 2145.480 612.920 ;
        RECT 53.880 610.200 2145.480 611.600 ;
        RECT 53.470 602.760 2145.480 610.200 ;
        RECT 53.470 601.360 2145.080 602.760 ;
        RECT 53.470 600.040 2145.480 601.360 ;
        RECT 53.880 598.640 2145.480 600.040 ;
        RECT 53.470 591.880 2145.480 598.640 ;
        RECT 53.470 590.480 2145.080 591.880 ;
        RECT 53.470 589.160 2145.480 590.480 ;
        RECT 53.880 587.760 2145.480 589.160 ;
        RECT 53.470 580.320 2145.480 587.760 ;
        RECT 53.470 578.920 2145.080 580.320 ;
        RECT 53.470 577.600 2145.480 578.920 ;
        RECT 53.880 576.200 2145.480 577.600 ;
        RECT 53.470 569.440 2145.480 576.200 ;
        RECT 53.470 568.040 2145.080 569.440 ;
        RECT 53.470 566.720 2145.480 568.040 ;
        RECT 53.880 565.320 2145.480 566.720 ;
        RECT 53.470 557.880 2145.480 565.320 ;
        RECT 53.470 556.480 2145.080 557.880 ;
        RECT 53.470 555.160 2145.480 556.480 ;
        RECT 53.880 553.760 2145.480 555.160 ;
        RECT 53.470 546.320 2145.480 553.760 ;
        RECT 53.470 544.920 2145.080 546.320 ;
        RECT 53.470 544.280 2145.480 544.920 ;
        RECT 53.880 542.880 2145.480 544.280 ;
        RECT 53.470 535.440 2145.480 542.880 ;
        RECT 53.470 534.040 2145.080 535.440 ;
        RECT 53.470 532.720 2145.480 534.040 ;
        RECT 53.880 531.320 2145.480 532.720 ;
        RECT 53.470 523.880 2145.480 531.320 ;
        RECT 53.470 522.480 2145.080 523.880 ;
        RECT 53.470 521.840 2145.480 522.480 ;
        RECT 53.880 520.440 2145.480 521.840 ;
        RECT 53.470 513.000 2145.480 520.440 ;
        RECT 53.470 511.600 2145.080 513.000 ;
        RECT 53.470 510.280 2145.480 511.600 ;
        RECT 53.880 508.880 2145.480 510.280 ;
        RECT 53.470 501.440 2145.480 508.880 ;
        RECT 53.470 500.040 2145.080 501.440 ;
        RECT 53.470 499.400 2145.480 500.040 ;
        RECT 53.880 498.000 2145.480 499.400 ;
        RECT 53.470 490.560 2145.480 498.000 ;
        RECT 53.470 489.160 2145.080 490.560 ;
        RECT 53.470 487.840 2145.480 489.160 ;
        RECT 53.880 486.440 2145.480 487.840 ;
        RECT 53.470 479.000 2145.480 486.440 ;
        RECT 53.470 477.600 2145.080 479.000 ;
        RECT 53.470 476.960 2145.480 477.600 ;
        RECT 53.880 475.560 2145.480 476.960 ;
        RECT 53.470 467.440 2145.480 475.560 ;
        RECT 53.470 466.040 2145.080 467.440 ;
        RECT 53.470 465.400 2145.480 466.040 ;
        RECT 53.880 464.000 2145.480 465.400 ;
        RECT 53.470 456.560 2145.480 464.000 ;
        RECT 53.470 455.160 2145.080 456.560 ;
        RECT 53.470 454.520 2145.480 455.160 ;
        RECT 53.880 453.120 2145.480 454.520 ;
        RECT 53.470 445.000 2145.480 453.120 ;
        RECT 53.470 443.600 2145.080 445.000 ;
        RECT 53.470 442.960 2145.480 443.600 ;
        RECT 53.880 441.560 2145.480 442.960 ;
        RECT 53.470 434.120 2145.480 441.560 ;
        RECT 53.470 432.720 2145.080 434.120 ;
        RECT 53.470 432.080 2145.480 432.720 ;
        RECT 53.880 430.680 2145.480 432.080 ;
        RECT 53.470 422.560 2145.480 430.680 ;
        RECT 53.470 421.160 2145.080 422.560 ;
        RECT 53.470 420.520 2145.480 421.160 ;
        RECT 53.880 419.120 2145.480 420.520 ;
        RECT 53.470 411.000 2145.480 419.120 ;
        RECT 53.470 409.640 2145.080 411.000 ;
        RECT 53.880 409.600 2145.080 409.640 ;
        RECT 53.880 408.240 2145.480 409.600 ;
        RECT 53.470 400.120 2145.480 408.240 ;
        RECT 53.470 398.720 2145.080 400.120 ;
        RECT 53.470 398.080 2145.480 398.720 ;
        RECT 53.880 396.680 2145.480 398.080 ;
        RECT 53.470 388.560 2145.480 396.680 ;
        RECT 53.470 387.200 2145.080 388.560 ;
        RECT 53.880 387.160 2145.080 387.200 ;
        RECT 53.880 385.800 2145.480 387.160 ;
        RECT 53.470 377.680 2145.480 385.800 ;
        RECT 53.470 376.280 2145.080 377.680 ;
        RECT 53.470 375.640 2145.480 376.280 ;
        RECT 53.880 374.240 2145.480 375.640 ;
        RECT 53.470 366.120 2145.480 374.240 ;
        RECT 53.470 364.760 2145.080 366.120 ;
        RECT 53.880 364.720 2145.080 364.760 ;
        RECT 53.880 363.360 2145.480 364.720 ;
        RECT 53.470 354.560 2145.480 363.360 ;
        RECT 53.470 353.200 2145.080 354.560 ;
        RECT 53.880 353.160 2145.080 353.200 ;
        RECT 53.880 351.800 2145.480 353.160 ;
        RECT 53.470 343.680 2145.480 351.800 ;
        RECT 53.470 342.320 2145.080 343.680 ;
        RECT 53.880 342.280 2145.080 342.320 ;
        RECT 53.880 340.920 2145.480 342.280 ;
        RECT 53.470 332.120 2145.480 340.920 ;
        RECT 53.470 330.760 2145.080 332.120 ;
        RECT 53.880 330.720 2145.080 330.760 ;
        RECT 53.880 329.360 2145.480 330.720 ;
        RECT 53.470 321.240 2145.480 329.360 ;
        RECT 53.470 319.880 2145.080 321.240 ;
        RECT 53.880 319.840 2145.080 319.880 ;
        RECT 53.880 318.480 2145.480 319.840 ;
        RECT 53.470 309.680 2145.480 318.480 ;
        RECT 53.470 308.320 2145.080 309.680 ;
        RECT 53.880 308.280 2145.080 308.320 ;
        RECT 53.880 306.920 2145.480 308.280 ;
        RECT 53.470 298.120 2145.480 306.920 ;
        RECT 53.470 297.440 2145.080 298.120 ;
        RECT 53.880 296.720 2145.080 297.440 ;
        RECT 53.880 296.040 2145.480 296.720 ;
        RECT 53.470 287.240 2145.480 296.040 ;
        RECT 53.470 285.880 2145.080 287.240 ;
        RECT 53.880 285.840 2145.080 285.880 ;
        RECT 53.880 284.480 2145.480 285.840 ;
        RECT 53.470 275.680 2145.480 284.480 ;
        RECT 53.470 275.000 2145.080 275.680 ;
        RECT 53.880 274.280 2145.080 275.000 ;
        RECT 53.880 273.600 2145.480 274.280 ;
        RECT 53.470 264.800 2145.480 273.600 ;
        RECT 53.470 263.440 2145.080 264.800 ;
        RECT 53.880 263.400 2145.080 263.440 ;
        RECT 53.880 262.040 2145.480 263.400 ;
        RECT 53.470 253.240 2145.480 262.040 ;
        RECT 53.470 252.560 2145.080 253.240 ;
        RECT 53.880 251.840 2145.080 252.560 ;
        RECT 53.880 251.160 2145.480 251.840 ;
        RECT 53.470 242.360 2145.480 251.160 ;
        RECT 53.470 241.000 2145.080 242.360 ;
        RECT 53.880 240.960 2145.080 241.000 ;
        RECT 53.880 239.600 2145.480 240.960 ;
        RECT 53.470 230.800 2145.480 239.600 ;
        RECT 53.470 230.120 2145.080 230.800 ;
        RECT 53.880 229.400 2145.080 230.120 ;
        RECT 53.880 228.720 2145.480 229.400 ;
        RECT 53.470 219.240 2145.480 228.720 ;
        RECT 53.470 218.560 2145.080 219.240 ;
        RECT 53.880 217.840 2145.080 218.560 ;
        RECT 53.880 217.160 2145.480 217.840 ;
        RECT 53.470 208.360 2145.480 217.160 ;
        RECT 53.470 207.680 2145.080 208.360 ;
        RECT 53.880 206.960 2145.080 207.680 ;
        RECT 53.880 206.280 2145.480 206.960 ;
        RECT 53.470 196.800 2145.480 206.280 ;
        RECT 53.470 196.120 2145.080 196.800 ;
        RECT 53.880 195.400 2145.080 196.120 ;
        RECT 53.880 194.720 2145.480 195.400 ;
        RECT 53.470 185.920 2145.480 194.720 ;
        RECT 53.470 185.240 2145.080 185.920 ;
        RECT 53.880 184.520 2145.080 185.240 ;
        RECT 53.880 183.840 2145.480 184.520 ;
        RECT 53.470 174.360 2145.480 183.840 ;
        RECT 53.470 173.680 2145.080 174.360 ;
        RECT 53.880 172.960 2145.080 173.680 ;
        RECT 53.880 172.280 2145.480 172.960 ;
        RECT 53.470 162.800 2145.480 172.280 ;
        RECT 53.880 161.400 2145.080 162.800 ;
        RECT 53.470 151.920 2145.480 161.400 ;
        RECT 53.470 151.240 2145.080 151.920 ;
        RECT 53.880 150.520 2145.080 151.240 ;
        RECT 53.880 149.840 2145.480 150.520 ;
        RECT 53.470 140.360 2145.480 149.840 ;
        RECT 53.880 138.960 2145.080 140.360 ;
        RECT 53.470 129.480 2145.480 138.960 ;
        RECT 53.470 128.800 2145.080 129.480 ;
        RECT 53.880 128.080 2145.080 128.800 ;
        RECT 53.880 127.400 2145.480 128.080 ;
        RECT 53.470 117.920 2145.480 127.400 ;
        RECT 53.880 116.520 2145.080 117.920 ;
        RECT 53.470 106.360 2145.480 116.520 ;
        RECT 53.880 104.960 2145.080 106.360 ;
        RECT 53.470 95.480 2145.480 104.960 ;
        RECT 53.880 94.080 2145.080 95.480 ;
        RECT 53.470 83.920 2145.480 94.080 ;
        RECT 53.880 82.520 2145.080 83.920 ;
        RECT 53.470 73.040 2145.480 82.520 ;
        RECT 53.880 71.640 2145.080 73.040 ;
        RECT 53.470 61.480 2145.480 71.640 ;
        RECT 53.880 60.080 2145.080 61.480 ;
        RECT 53.470 50.600 2145.480 60.080 ;
        RECT 53.880 49.200 2145.080 50.600 ;
        RECT 53.470 44.300 2145.480 49.200 ;
      LAYER met4 ;
        RECT 0.000 0.000 2198.860 2286.000 ;
      LAYER met5 ;
        RECT 0.000 70.610 2198.860 2286.000 ;
  END
END mac_tile
END LIBRARY

