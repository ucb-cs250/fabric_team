VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 266.785 BY 277.505 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 273.505 247.850 277.505 ;
    END
  END COUT
  PIN cb_e_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 2.760 266.785 3.360 ;
    END
  END cb_e_clb1_input[0]
  PIN cb_e_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 8.200 266.785 8.800 ;
    END
  END cb_e_clb1_input[1]
  PIN cb_e_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 14.320 266.785 14.920 ;
    END
  END cb_e_clb1_input[2]
  PIN cb_e_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 20.440 266.785 21.040 ;
    END
  END cb_e_clb1_input[3]
  PIN cb_e_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 26.560 266.785 27.160 ;
    END
  END cb_e_clb1_input[4]
  PIN cb_e_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 32.680 266.785 33.280 ;
    END
  END cb_e_clb1_input[5]
  PIN cb_e_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 38.800 266.785 39.400 ;
    END
  END cb_e_clb1_input[6]
  PIN cb_e_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 44.920 266.785 45.520 ;
    END
  END cb_e_clb1_input[7]
  PIN cb_e_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 50.360 266.785 50.960 ;
    END
  END cb_e_clb1_input[8]
  PIN cb_e_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 56.480 266.785 57.080 ;
    END
  END cb_e_clb1_input[9]
  PIN cb_e_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 62.600 266.785 63.200 ;
    END
  END cb_e_clb1_output[0]
  PIN cb_e_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 68.720 266.785 69.320 ;
    END
  END cb_e_clb1_output[1]
  PIN cb_e_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 74.840 266.785 75.440 ;
    END
  END cb_e_clb1_output[2]
  PIN cb_e_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 80.960 266.785 81.560 ;
    END
  END cb_e_clb1_output[3]
  PIN cb_e_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END cb_e_single1_in[0]
  PIN cb_e_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END cb_e_single1_in[10]
  PIN cb_e_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END cb_e_single1_in[11]
  PIN cb_e_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END cb_e_single1_in[12]
  PIN cb_e_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END cb_e_single1_in[13]
  PIN cb_e_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END cb_e_single1_in[14]
  PIN cb_e_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END cb_e_single1_in[15]
  PIN cb_e_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END cb_e_single1_in[1]
  PIN cb_e_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END cb_e_single1_in[2]
  PIN cb_e_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END cb_e_single1_in[3]
  PIN cb_e_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END cb_e_single1_in[4]
  PIN cb_e_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END cb_e_single1_in[5]
  PIN cb_e_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END cb_e_single1_in[6]
  PIN cb_e_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END cb_e_single1_in[7]
  PIN cb_e_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END cb_e_single1_in[8]
  PIN cb_e_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END cb_e_single1_in[9]
  PIN cb_e_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END cb_e_single1_out[0]
  PIN cb_e_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END cb_e_single1_out[10]
  PIN cb_e_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END cb_e_single1_out[11]
  PIN cb_e_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END cb_e_single1_out[12]
  PIN cb_e_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END cb_e_single1_out[13]
  PIN cb_e_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END cb_e_single1_out[14]
  PIN cb_e_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END cb_e_single1_out[15]
  PIN cb_e_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cb_e_single1_out[1]
  PIN cb_e_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END cb_e_single1_out[2]
  PIN cb_e_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cb_e_single1_out[3]
  PIN cb_e_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cb_e_single1_out[4]
  PIN cb_e_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END cb_e_single1_out[5]
  PIN cb_e_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cb_e_single1_out[6]
  PIN cb_e_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END cb_e_single1_out[7]
  PIN cb_e_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END cb_e_single1_out[8]
  PIN cb_e_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END cb_e_single1_out[9]
  PIN cb_n_clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 273.505 2.670 277.505 ;
    END
  END cb_n_clb1_input[0]
  PIN cb_n_clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 273.505 7.730 277.505 ;
    END
  END cb_n_clb1_input[1]
  PIN cb_n_clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 273.505 13.250 277.505 ;
    END
  END cb_n_clb1_input[2]
  PIN cb_n_clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 273.505 18.310 277.505 ;
    END
  END cb_n_clb1_input[3]
  PIN cb_n_clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 273.505 23.830 277.505 ;
    END
  END cb_n_clb1_input[4]
  PIN cb_n_clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 273.505 29.350 277.505 ;
    END
  END cb_n_clb1_input[5]
  PIN cb_n_clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 273.505 34.410 277.505 ;
    END
  END cb_n_clb1_input[6]
  PIN cb_n_clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 273.505 39.930 277.505 ;
    END
  END cb_n_clb1_input[7]
  PIN cb_n_clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 273.505 44.990 277.505 ;
    END
  END cb_n_clb1_input[8]
  PIN cb_n_clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 273.505 50.510 277.505 ;
    END
  END cb_n_clb1_input[9]
  PIN cb_n_clb1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 273.505 56.030 277.505 ;
    END
  END cb_n_clb1_output[0]
  PIN cb_n_clb1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 273.505 61.090 277.505 ;
    END
  END cb_n_clb1_output[1]
  PIN cb_n_clb1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 273.505 66.610 277.505 ;
    END
  END cb_n_clb1_output[2]
  PIN cb_n_clb1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 273.505 71.670 277.505 ;
    END
  END cb_n_clb1_output[3]
  PIN cb_n_single1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END cb_n_single1_in[0]
  PIN cb_n_single1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END cb_n_single1_in[10]
  PIN cb_n_single1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END cb_n_single1_in[11]
  PIN cb_n_single1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END cb_n_single1_in[12]
  PIN cb_n_single1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END cb_n_single1_in[13]
  PIN cb_n_single1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END cb_n_single1_in[14]
  PIN cb_n_single1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END cb_n_single1_in[15]
  PIN cb_n_single1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END cb_n_single1_in[1]
  PIN cb_n_single1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END cb_n_single1_in[2]
  PIN cb_n_single1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END cb_n_single1_in[3]
  PIN cb_n_single1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END cb_n_single1_in[4]
  PIN cb_n_single1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END cb_n_single1_in[5]
  PIN cb_n_single1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END cb_n_single1_in[6]
  PIN cb_n_single1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END cb_n_single1_in[7]
  PIN cb_n_single1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END cb_n_single1_in[8]
  PIN cb_n_single1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END cb_n_single1_in[9]
  PIN cb_n_single1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END cb_n_single1_out[0]
  PIN cb_n_single1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END cb_n_single1_out[10]
  PIN cb_n_single1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END cb_n_single1_out[11]
  PIN cb_n_single1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END cb_n_single1_out[12]
  PIN cb_n_single1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END cb_n_single1_out[13]
  PIN cb_n_single1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END cb_n_single1_out[14]
  PIN cb_n_single1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END cb_n_single1_out[15]
  PIN cb_n_single1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END cb_n_single1_out[1]
  PIN cb_n_single1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END cb_n_single1_out[2]
  PIN cb_n_single1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END cb_n_single1_out[3]
  PIN cb_n_single1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END cb_n_single1_out[4]
  PIN cb_n_single1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END cb_n_single1_out[5]
  PIN cb_n_single1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END cb_n_single1_out[6]
  PIN cb_n_single1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END cb_n_single1_out[7]
  PIN cb_n_single1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END cb_n_single1_out[8]
  PIN cb_n_single1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END cb_n_single1_out[9]
  PIN cfg_bit_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END cfg_bit_in
  PIN cfg_bit_in_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END cfg_bit_in_valid
  PIN cfg_bit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 273.505 258.430 277.505 ;
    END
  END cfg_bit_out
  PIN cfg_bit_out_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 273.505 263.950 277.505 ;
    END
  END cfg_bit_out_valid
  PIN cfg_in_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END cfg_in_start
  PIN cfg_out_start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 273.505 253.370 277.505 ;
    END
  END cfg_out_start
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END clb_south_out[3]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END clb_west_out[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END clk
  PIN crst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END crst
  PIN sb_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 87.080 266.785 87.680 ;
    END
  END sb_east_in[0]
  PIN sb_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 146.920 266.785 147.520 ;
    END
  END sb_east_in[10]
  PIN sb_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 153.040 266.785 153.640 ;
    END
  END sb_east_in[11]
  PIN sb_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 159.160 266.785 159.760 ;
    END
  END sb_east_in[12]
  PIN sb_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 165.280 266.785 165.880 ;
    END
  END sb_east_in[13]
  PIN sb_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 171.400 266.785 172.000 ;
    END
  END sb_east_in[14]
  PIN sb_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 177.520 266.785 178.120 ;
    END
  END sb_east_in[15]
  PIN sb_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 93.200 266.785 93.800 ;
    END
  END sb_east_in[1]
  PIN sb_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 98.640 266.785 99.240 ;
    END
  END sb_east_in[2]
  PIN sb_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 104.760 266.785 105.360 ;
    END
  END sb_east_in[3]
  PIN sb_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 110.880 266.785 111.480 ;
    END
  END sb_east_in[4]
  PIN sb_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 117.000 266.785 117.600 ;
    END
  END sb_east_in[5]
  PIN sb_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 123.120 266.785 123.720 ;
    END
  END sb_east_in[6]
  PIN sb_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 129.240 266.785 129.840 ;
    END
  END sb_east_in[7]
  PIN sb_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 135.360 266.785 135.960 ;
    END
  END sb_east_in[8]
  PIN sb_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 141.480 266.785 142.080 ;
    END
  END sb_east_in[9]
  PIN sb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 183.640 266.785 184.240 ;
    END
  END sb_east_out[0]
  PIN sb_east_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 243.480 266.785 244.080 ;
    END
  END sb_east_out[10]
  PIN sb_east_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 249.600 266.785 250.200 ;
    END
  END sb_east_out[11]
  PIN sb_east_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 255.720 266.785 256.320 ;
    END
  END sb_east_out[12]
  PIN sb_east_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 261.840 266.785 262.440 ;
    END
  END sb_east_out[13]
  PIN sb_east_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 267.960 266.785 268.560 ;
    END
  END sb_east_out[14]
  PIN sb_east_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 274.080 266.785 274.680 ;
    END
  END sb_east_out[15]
  PIN sb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 189.080 266.785 189.680 ;
    END
  END sb_east_out[1]
  PIN sb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 195.200 266.785 195.800 ;
    END
  END sb_east_out[2]
  PIN sb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 201.320 266.785 201.920 ;
    END
  END sb_east_out[3]
  PIN sb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 207.440 266.785 208.040 ;
    END
  END sb_east_out[4]
  PIN sb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 213.560 266.785 214.160 ;
    END
  END sb_east_out[5]
  PIN sb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 219.680 266.785 220.280 ;
    END
  END sb_east_out[6]
  PIN sb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 225.800 266.785 226.400 ;
    END
  END sb_east_out[7]
  PIN sb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 231.920 266.785 232.520 ;
    END
  END sb_east_out[8]
  PIN sb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.785 237.360 266.785 237.960 ;
    END
  END sb_east_out[9]
  PIN sb_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 273.505 77.190 277.505 ;
    END
  END sb_north_in[0]
  PIN sb_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 273.505 130.550 277.505 ;
    END
  END sb_north_in[10]
  PIN sb_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 273.505 136.070 277.505 ;
    END
  END sb_north_in[11]
  PIN sb_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 273.505 141.130 277.505 ;
    END
  END sb_north_in[12]
  PIN sb_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 273.505 146.650 277.505 ;
    END
  END sb_north_in[13]
  PIN sb_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 273.505 151.710 277.505 ;
    END
  END sb_north_in[14]
  PIN sb_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 273.505 157.230 277.505 ;
    END
  END sb_north_in[15]
  PIN sb_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 273.505 82.710 277.505 ;
    END
  END sb_north_in[1]
  PIN sb_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 273.505 87.770 277.505 ;
    END
  END sb_north_in[2]
  PIN sb_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 273.505 93.290 277.505 ;
    END
  END sb_north_in[3]
  PIN sb_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 273.505 98.350 277.505 ;
    END
  END sb_north_in[4]
  PIN sb_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 273.505 103.870 277.505 ;
    END
  END sb_north_in[5]
  PIN sb_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 273.505 109.390 277.505 ;
    END
  END sb_north_in[6]
  PIN sb_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 273.505 114.450 277.505 ;
    END
  END sb_north_in[7]
  PIN sb_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 273.505 119.970 277.505 ;
    END
  END sb_north_in[8]
  PIN sb_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 273.505 125.030 277.505 ;
    END
  END sb_north_in[9]
  PIN sb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 273.505 162.750 277.505 ;
    END
  END sb_north_out[0]
  PIN sb_north_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 273.505 216.110 277.505 ;
    END
  END sb_north_out[10]
  PIN sb_north_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 273.505 221.170 277.505 ;
    END
  END sb_north_out[11]
  PIN sb_north_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 273.505 226.690 277.505 ;
    END
  END sb_north_out[12]
  PIN sb_north_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 273.505 231.750 277.505 ;
    END
  END sb_north_out[13]
  PIN sb_north_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 273.505 237.270 277.505 ;
    END
  END sb_north_out[14]
  PIN sb_north_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 273.505 242.790 277.505 ;
    END
  END sb_north_out[15]
  PIN sb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 273.505 167.810 277.505 ;
    END
  END sb_north_out[1]
  PIN sb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 273.505 173.330 277.505 ;
    END
  END sb_north_out[2]
  PIN sb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 273.505 178.390 277.505 ;
    END
  END sb_north_out[3]
  PIN sb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 273.505 183.910 277.505 ;
    END
  END sb_north_out[4]
  PIN sb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 273.505 189.430 277.505 ;
    END
  END sb_north_out[5]
  PIN sb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 273.505 194.490 277.505 ;
    END
  END sb_north_out[6]
  PIN sb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 273.505 200.010 277.505 ;
    END
  END sb_north_out[7]
  PIN sb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 273.505 205.070 277.505 ;
    END
  END sb_north_out[8]
  PIN sb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 273.505 210.590 277.505 ;
    END
  END sb_north_out[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 266.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 266.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 266.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 266.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 6.885 261.595 268.175 ;
      LAYER met1 ;
        RECT 2.370 6.500 263.970 268.900 ;
      LAYER met2 ;
        RECT 2.950 273.225 7.170 274.565 ;
        RECT 8.010 273.225 12.690 274.565 ;
        RECT 13.530 273.225 17.750 274.565 ;
        RECT 18.590 273.225 23.270 274.565 ;
        RECT 24.110 273.225 28.790 274.565 ;
        RECT 29.630 273.225 33.850 274.565 ;
        RECT 34.690 273.225 39.370 274.565 ;
        RECT 40.210 273.225 44.430 274.565 ;
        RECT 45.270 273.225 49.950 274.565 ;
        RECT 50.790 273.225 55.470 274.565 ;
        RECT 56.310 273.225 60.530 274.565 ;
        RECT 61.370 273.225 66.050 274.565 ;
        RECT 66.890 273.225 71.110 274.565 ;
        RECT 71.950 273.225 76.630 274.565 ;
        RECT 77.470 273.225 82.150 274.565 ;
        RECT 82.990 273.225 87.210 274.565 ;
        RECT 88.050 273.225 92.730 274.565 ;
        RECT 93.570 273.225 97.790 274.565 ;
        RECT 98.630 273.225 103.310 274.565 ;
        RECT 104.150 273.225 108.830 274.565 ;
        RECT 109.670 273.225 113.890 274.565 ;
        RECT 114.730 273.225 119.410 274.565 ;
        RECT 120.250 273.225 124.470 274.565 ;
        RECT 125.310 273.225 129.990 274.565 ;
        RECT 130.830 273.225 135.510 274.565 ;
        RECT 136.350 273.225 140.570 274.565 ;
        RECT 141.410 273.225 146.090 274.565 ;
        RECT 146.930 273.225 151.150 274.565 ;
        RECT 151.990 273.225 156.670 274.565 ;
        RECT 157.510 273.225 162.190 274.565 ;
        RECT 163.030 273.225 167.250 274.565 ;
        RECT 168.090 273.225 172.770 274.565 ;
        RECT 173.610 273.225 177.830 274.565 ;
        RECT 178.670 273.225 183.350 274.565 ;
        RECT 184.190 273.225 188.870 274.565 ;
        RECT 189.710 273.225 193.930 274.565 ;
        RECT 194.770 273.225 199.450 274.565 ;
        RECT 200.290 273.225 204.510 274.565 ;
        RECT 205.350 273.225 210.030 274.565 ;
        RECT 210.870 273.225 215.550 274.565 ;
        RECT 216.390 273.225 220.610 274.565 ;
        RECT 221.450 273.225 226.130 274.565 ;
        RECT 226.970 273.225 231.190 274.565 ;
        RECT 232.030 273.225 236.710 274.565 ;
        RECT 237.550 273.225 242.230 274.565 ;
        RECT 243.070 273.225 247.290 274.565 ;
        RECT 248.130 273.225 252.810 274.565 ;
        RECT 253.650 273.225 257.870 274.565 ;
        RECT 258.710 273.225 263.390 274.565 ;
        RECT 2.400 4.280 263.940 273.225 ;
        RECT 2.950 2.875 7.170 4.280 ;
        RECT 8.010 2.875 12.230 4.280 ;
        RECT 13.070 2.875 17.290 4.280 ;
        RECT 18.130 2.875 22.350 4.280 ;
        RECT 23.190 2.875 27.410 4.280 ;
        RECT 28.250 2.875 32.470 4.280 ;
        RECT 33.310 2.875 37.990 4.280 ;
        RECT 38.830 2.875 43.050 4.280 ;
        RECT 43.890 2.875 48.110 4.280 ;
        RECT 48.950 2.875 53.170 4.280 ;
        RECT 54.010 2.875 58.230 4.280 ;
        RECT 59.070 2.875 63.290 4.280 ;
        RECT 64.130 2.875 68.810 4.280 ;
        RECT 69.650 2.875 73.870 4.280 ;
        RECT 74.710 2.875 78.930 4.280 ;
        RECT 79.770 2.875 83.990 4.280 ;
        RECT 84.830 2.875 89.050 4.280 ;
        RECT 89.890 2.875 94.110 4.280 ;
        RECT 94.950 2.875 99.170 4.280 ;
        RECT 100.010 2.875 104.690 4.280 ;
        RECT 105.530 2.875 109.750 4.280 ;
        RECT 110.590 2.875 114.810 4.280 ;
        RECT 115.650 2.875 119.870 4.280 ;
        RECT 120.710 2.875 124.930 4.280 ;
        RECT 125.770 2.875 129.990 4.280 ;
        RECT 130.830 2.875 135.510 4.280 ;
        RECT 136.350 2.875 140.570 4.280 ;
        RECT 141.410 2.875 145.630 4.280 ;
        RECT 146.470 2.875 150.690 4.280 ;
        RECT 151.530 2.875 155.750 4.280 ;
        RECT 156.590 2.875 160.810 4.280 ;
        RECT 161.650 2.875 165.870 4.280 ;
        RECT 166.710 2.875 171.390 4.280 ;
        RECT 172.230 2.875 176.450 4.280 ;
        RECT 177.290 2.875 181.510 4.280 ;
        RECT 182.350 2.875 186.570 4.280 ;
        RECT 187.410 2.875 191.630 4.280 ;
        RECT 192.470 2.875 196.690 4.280 ;
        RECT 197.530 2.875 202.210 4.280 ;
        RECT 203.050 2.875 207.270 4.280 ;
        RECT 208.110 2.875 212.330 4.280 ;
        RECT 213.170 2.875 217.390 4.280 ;
        RECT 218.230 2.875 222.450 4.280 ;
        RECT 223.290 2.875 227.510 4.280 ;
        RECT 228.350 2.875 232.570 4.280 ;
        RECT 233.410 2.875 238.090 4.280 ;
        RECT 238.930 2.875 243.150 4.280 ;
        RECT 243.990 2.875 248.210 4.280 ;
        RECT 249.050 2.875 253.270 4.280 ;
        RECT 254.110 2.875 258.330 4.280 ;
        RECT 259.170 2.875 263.390 4.280 ;
      LAYER met3 ;
        RECT 4.400 273.680 262.385 274.545 ;
        RECT 4.000 268.960 262.785 273.680 ;
        RECT 4.400 267.560 262.385 268.960 ;
        RECT 4.000 262.840 262.785 267.560 ;
        RECT 4.400 261.440 262.385 262.840 ;
        RECT 4.000 256.720 262.785 261.440 ;
        RECT 4.400 255.320 262.385 256.720 ;
        RECT 4.000 250.600 262.785 255.320 ;
        RECT 4.400 249.200 262.385 250.600 ;
        RECT 4.000 244.480 262.785 249.200 ;
        RECT 4.400 243.080 262.385 244.480 ;
        RECT 4.000 238.360 262.785 243.080 ;
        RECT 4.400 236.960 262.385 238.360 ;
        RECT 4.000 232.920 262.785 236.960 ;
        RECT 4.400 231.520 262.385 232.920 ;
        RECT 4.000 226.800 262.785 231.520 ;
        RECT 4.400 225.400 262.385 226.800 ;
        RECT 4.000 220.680 262.785 225.400 ;
        RECT 4.400 219.280 262.385 220.680 ;
        RECT 4.000 214.560 262.785 219.280 ;
        RECT 4.400 213.160 262.385 214.560 ;
        RECT 4.000 208.440 262.785 213.160 ;
        RECT 4.400 207.040 262.385 208.440 ;
        RECT 4.000 202.320 262.785 207.040 ;
        RECT 4.400 200.920 262.385 202.320 ;
        RECT 4.000 196.200 262.785 200.920 ;
        RECT 4.400 194.800 262.385 196.200 ;
        RECT 4.000 190.080 262.785 194.800 ;
        RECT 4.400 188.680 262.385 190.080 ;
        RECT 4.000 184.640 262.785 188.680 ;
        RECT 4.400 183.240 262.385 184.640 ;
        RECT 4.000 178.520 262.785 183.240 ;
        RECT 4.400 177.120 262.385 178.520 ;
        RECT 4.000 172.400 262.785 177.120 ;
        RECT 4.400 171.000 262.385 172.400 ;
        RECT 4.000 166.280 262.785 171.000 ;
        RECT 4.400 164.880 262.385 166.280 ;
        RECT 4.000 160.160 262.785 164.880 ;
        RECT 4.400 158.760 262.385 160.160 ;
        RECT 4.000 154.040 262.785 158.760 ;
        RECT 4.400 152.640 262.385 154.040 ;
        RECT 4.000 147.920 262.785 152.640 ;
        RECT 4.400 146.520 262.385 147.920 ;
        RECT 4.000 142.480 262.785 146.520 ;
        RECT 4.400 141.080 262.385 142.480 ;
        RECT 4.000 136.360 262.785 141.080 ;
        RECT 4.400 134.960 262.385 136.360 ;
        RECT 4.000 130.240 262.785 134.960 ;
        RECT 4.400 128.840 262.385 130.240 ;
        RECT 4.000 124.120 262.785 128.840 ;
        RECT 4.400 122.720 262.385 124.120 ;
        RECT 4.000 118.000 262.785 122.720 ;
        RECT 4.400 116.600 262.385 118.000 ;
        RECT 4.000 111.880 262.785 116.600 ;
        RECT 4.400 110.480 262.385 111.880 ;
        RECT 4.000 105.760 262.785 110.480 ;
        RECT 4.400 104.360 262.385 105.760 ;
        RECT 4.000 99.640 262.785 104.360 ;
        RECT 4.400 98.240 262.385 99.640 ;
        RECT 4.000 94.200 262.785 98.240 ;
        RECT 4.400 92.800 262.385 94.200 ;
        RECT 4.000 88.080 262.785 92.800 ;
        RECT 4.400 86.680 262.385 88.080 ;
        RECT 4.000 81.960 262.785 86.680 ;
        RECT 4.400 80.560 262.385 81.960 ;
        RECT 4.000 75.840 262.785 80.560 ;
        RECT 4.400 74.440 262.385 75.840 ;
        RECT 4.000 69.720 262.785 74.440 ;
        RECT 4.400 68.320 262.385 69.720 ;
        RECT 4.000 63.600 262.785 68.320 ;
        RECT 4.400 62.200 262.385 63.600 ;
        RECT 4.000 57.480 262.785 62.200 ;
        RECT 4.400 56.080 262.385 57.480 ;
        RECT 4.000 51.360 262.785 56.080 ;
        RECT 4.400 49.960 262.385 51.360 ;
        RECT 4.000 45.920 262.785 49.960 ;
        RECT 4.400 44.520 262.385 45.920 ;
        RECT 4.000 39.800 262.785 44.520 ;
        RECT 4.400 38.400 262.385 39.800 ;
        RECT 4.000 33.680 262.785 38.400 ;
        RECT 4.400 32.280 262.385 33.680 ;
        RECT 4.000 27.560 262.785 32.280 ;
        RECT 4.400 26.160 262.385 27.560 ;
        RECT 4.000 21.440 262.785 26.160 ;
        RECT 4.400 20.040 262.385 21.440 ;
        RECT 4.000 15.320 262.785 20.040 ;
        RECT 4.400 13.920 262.385 15.320 ;
        RECT 4.000 9.200 262.785 13.920 ;
        RECT 4.400 7.800 262.385 9.200 ;
        RECT 4.000 3.760 262.785 7.800 ;
        RECT 4.400 2.895 262.385 3.760 ;
      LAYER met4 ;
        RECT 8.575 11.055 20.640 262.985 ;
        RECT 23.040 11.055 97.440 262.985 ;
        RECT 99.840 11.055 174.240 262.985 ;
        RECT 176.640 11.055 251.040 262.985 ;
        RECT 253.440 11.055 258.650 262.985 ;
      LAYER met5 ;
        RECT 163.420 17.900 258.860 19.500 ;
  END
END clb_tile
END LIBRARY

