VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block_east
  CLASS BLOCK ;
  FOREIGN baked_connection_block_east ;
  ORIGIN 0.000 0.000 ;
  SIZE 254.225 BY 264.945 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.190 260.945 246.470 264.945 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 7.520 254.225 8.120 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 22.480 254.225 23.080 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 38.120 254.225 38.720 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 53.760 254.225 54.360 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 69.400 254.225 70.000 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 85.040 254.225 85.640 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 100.680 254.225 101.280 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 116.320 254.225 116.920 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 131.960 254.225 132.560 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 147.600 254.225 148.200 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 163.240 254.225 163.840 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 250.225 178.880 254.225 179.480 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 194.520 254.225 195.120 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 210.160 254.225 210.760 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 225.800 254.225 226.400 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 241.440 254.225 242.040 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 250.225 257.080 254.225 257.680 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 260.945 119.050 264.945 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 134.870 260.945 135.150 264.945 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 150.970 260.945 151.250 264.945 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 260.945 166.890 264.945 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 182.710 260.945 182.990 264.945 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 198.350 260.945 198.630 264.945 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 214.450 260.945 214.730 264.945 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 230.090 260.945 230.370 264.945 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END double1[7]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 260.945 23.830 264.945 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 260.945 8.190 264.945 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 260.945 39.930 264.945 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 260.945 55.570 264.945 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 260.945 71.670 264.945 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 260.945 87.310 264.945 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 103.130 260.945 103.410 264.945 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 253.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 253.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 249.175 253.045 ;
      LAYER met1 ;
        RECT 5.520 7.860 249.250 253.200 ;
      LAYER met2 ;
        RECT 7.000 260.665 7.630 260.945 ;
        RECT 8.470 260.665 23.270 260.945 ;
        RECT 24.110 260.665 39.370 260.945 ;
        RECT 40.210 260.665 55.010 260.945 ;
        RECT 55.850 260.665 71.110 260.945 ;
        RECT 71.950 260.665 86.750 260.945 ;
        RECT 87.590 260.665 102.850 260.945 ;
        RECT 103.690 260.665 118.490 260.945 ;
        RECT 119.330 260.665 134.590 260.945 ;
        RECT 135.430 260.665 150.690 260.945 ;
        RECT 151.530 260.665 166.330 260.945 ;
        RECT 167.170 260.665 182.430 260.945 ;
        RECT 183.270 260.665 198.070 260.945 ;
        RECT 198.910 260.665 214.170 260.945 ;
        RECT 215.010 260.665 229.810 260.945 ;
        RECT 230.650 260.665 245.910 260.945 ;
        RECT 246.750 260.665 249.230 260.945 ;
        RECT 7.000 4.280 249.230 260.665 ;
        RECT 7.000 4.000 8.550 4.280 ;
        RECT 9.390 4.000 26.490 4.280 ;
        RECT 27.330 4.000 44.890 4.280 ;
        RECT 45.730 4.000 62.830 4.280 ;
        RECT 63.670 4.000 81.230 4.280 ;
        RECT 82.070 4.000 99.170 4.280 ;
        RECT 100.010 4.000 117.570 4.280 ;
        RECT 118.410 4.000 135.510 4.280 ;
        RECT 136.350 4.000 153.910 4.280 ;
        RECT 154.750 4.000 171.850 4.280 ;
        RECT 172.690 4.000 190.250 4.280 ;
        RECT 191.090 4.000 208.190 4.280 ;
        RECT 209.030 4.000 226.590 4.280 ;
        RECT 227.430 4.000 244.530 4.280 ;
        RECT 245.370 4.000 249.230 4.280 ;
      LAYER met3 ;
        RECT 4.400 256.680 249.825 257.545 ;
        RECT 4.000 242.440 250.225 256.680 ;
        RECT 4.400 241.040 249.825 242.440 ;
        RECT 4.000 226.800 250.225 241.040 ;
        RECT 4.400 225.400 249.825 226.800 ;
        RECT 4.000 211.160 250.225 225.400 ;
        RECT 4.400 209.760 249.825 211.160 ;
        RECT 4.000 195.520 250.225 209.760 ;
        RECT 4.400 194.120 249.825 195.520 ;
        RECT 4.000 179.880 250.225 194.120 ;
        RECT 4.400 178.480 249.825 179.880 ;
        RECT 4.000 164.240 250.225 178.480 ;
        RECT 4.400 162.840 249.825 164.240 ;
        RECT 4.000 148.600 250.225 162.840 ;
        RECT 4.400 147.200 249.825 148.600 ;
        RECT 4.000 132.960 250.225 147.200 ;
        RECT 4.400 131.560 249.825 132.960 ;
        RECT 4.000 117.320 250.225 131.560 ;
        RECT 4.400 115.920 249.825 117.320 ;
        RECT 4.000 101.680 250.225 115.920 ;
        RECT 4.400 100.280 249.825 101.680 ;
        RECT 4.000 86.040 250.225 100.280 ;
        RECT 4.400 84.640 249.825 86.040 ;
        RECT 4.000 70.400 250.225 84.640 ;
        RECT 4.400 69.000 249.825 70.400 ;
        RECT 4.000 54.760 250.225 69.000 ;
        RECT 4.400 53.360 249.825 54.760 ;
        RECT 4.000 39.120 250.225 53.360 ;
        RECT 4.400 37.720 249.825 39.120 ;
        RECT 4.000 23.480 250.225 37.720 ;
        RECT 4.400 22.080 249.825 23.480 ;
        RECT 4.000 8.520 250.225 22.080 ;
        RECT 4.400 7.655 249.825 8.520 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 253.200 ;
  END
END baked_connection_block_east
END LIBRARY

