VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_slicel
  CLASS BLOCK ;
  FOREIGN baked_slicel ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.990 BY 236.710 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.550 232.710 207.830 236.710 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.510 232.710 219.790 236.710 ;
    END
  END carry_out
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 8.200 225.990 8.800 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END clk
  PIN higher_order_address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 232.710 5.890 236.710 ;
    END
  END higher_order_address[0]
  PIN higher_order_address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 232.710 17.390 236.710 ;
    END
  END higher_order_address[1]
  PIN lut_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 232.710 124.570 236.710 ;
    END
  END lut_output[0]
  PIN lut_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 232.710 136.530 236.710 ;
    END
  END lut_output[1]
  PIN lut_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END lut_output[2]
  PIN lut_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END lut_output[3]
  PIN lut_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 221.990 176.840 225.990 177.440 ;
    END
  END lut_output[4]
  PIN lut_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 221.990 193.840 225.990 194.440 ;
    END
  END lut_output[5]
  PIN lut_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END lut_output[6]
  PIN lut_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END lut_output[7]
  PIN lut_output_registered[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 232.710 148.490 236.710 ;
    END
  END lut_output_registered[0]
  PIN lut_output_registered[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.710 232.710 159.990 236.710 ;
    END
  END lut_output_registered[1]
  PIN lut_output_registered[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END lut_output_registered[2]
  PIN lut_output_registered[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END lut_output_registered[3]
  PIN lut_output_registered[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 221.990 210.840 225.990 211.440 ;
    END
  END lut_output_registered[4]
  PIN lut_output_registered[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 221.990 227.840 225.990 228.440 ;
    END
  END lut_output_registered[5]
  PIN lut_output_registered[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END lut_output_registered[6]
  PIN lut_output_registered[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END lut_output_registered[7]
  PIN luts_input[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 232.710 29.350 236.710 ;
    END
  END luts_input[0]
  PIN luts_input[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END luts_input[10]
  PIN luts_input[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END luts_input[11]
  PIN luts_input[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END luts_input[12]
  PIN luts_input[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END luts_input[13]
  PIN luts_input[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END luts_input[14]
  PIN luts_input[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END luts_input[15]
  PIN luts_input[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 41.520 225.990 42.120 ;
    END
  END luts_input[16]
  PIN luts_input[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 58.520 225.990 59.120 ;
    END
  END luts_input[17]
  PIN luts_input[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 75.520 225.990 76.120 ;
    END
  END luts_input[18]
  PIN luts_input[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 92.520 225.990 93.120 ;
    END
  END luts_input[19]
  PIN luts_input[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 232.710 41.310 236.710 ;
    END
  END luts_input[1]
  PIN luts_input[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 109.520 225.990 110.120 ;
    END
  END luts_input[20]
  PIN luts_input[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 126.520 225.990 127.120 ;
    END
  END luts_input[21]
  PIN luts_input[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 142.840 225.990 143.440 ;
    END
  END luts_input[22]
  PIN luts_input[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 159.840 225.990 160.440 ;
    END
  END luts_input[23]
  PIN luts_input[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END luts_input[24]
  PIN luts_input[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END luts_input[25]
  PIN luts_input[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END luts_input[26]
  PIN luts_input[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END luts_input[27]
  PIN luts_input[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END luts_input[28]
  PIN luts_input[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END luts_input[29]
  PIN luts_input[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 232.710 53.270 236.710 ;
    END
  END luts_input[2]
  PIN luts_input[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END luts_input[30]
  PIN luts_input[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END luts_input[31]
  PIN luts_input[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 232.710 65.230 236.710 ;
    END
  END luts_input[3]
  PIN luts_input[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 232.710 77.190 236.710 ;
    END
  END luts_input[4]
  PIN luts_input[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.410 232.710 88.690 236.710 ;
    END
  END luts_input[5]
  PIN luts_input[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 232.710 100.650 236.710 ;
    END
  END luts_input[6]
  PIN luts_input[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 232.710 112.610 236.710 ;
    END
  END luts_input[7]
  PIN luts_input[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END luts_input[8]
  PIN luts_input[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END luts_input[9]
  PIN reg_we
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END reg_we
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.590 232.710 195.870 236.710 ;
    END
  END set_in
  PIN set_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END set_in_soft
  PIN set_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END set_out
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.630 232.710 183.910 236.710 ;
    END
  END shift_in
  PIN shift_in_from_tile_bodge
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 221.990 24.520 225.990 25.120 ;
    END
  END shift_in_from_tile_bodge
  PIN shift_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END shift_in_soft
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END shift_out
  PIN shift_out_to_tile_bodge
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 171.670 232.710 171.950 236.710 ;
    END
  END shift_out_to_tile_bodge
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 226.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 226.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 220.340 225.845 ;
      LAYER met1 ;
        RECT 5.520 4.460 220.340 226.000 ;
      LAYER met2 ;
        RECT 6.170 232.430 16.830 232.710 ;
        RECT 17.670 232.430 28.790 232.710 ;
        RECT 29.630 232.430 40.750 232.710 ;
        RECT 41.590 232.430 52.710 232.710 ;
        RECT 53.550 232.430 64.670 232.710 ;
        RECT 65.510 232.430 76.630 232.710 ;
        RECT 77.470 232.430 88.130 232.710 ;
        RECT 88.970 232.430 100.090 232.710 ;
        RECT 100.930 232.430 112.050 232.710 ;
        RECT 112.890 232.430 124.010 232.710 ;
        RECT 124.850 232.430 135.970 232.710 ;
        RECT 136.810 232.430 147.930 232.710 ;
        RECT 148.770 232.430 159.430 232.710 ;
        RECT 160.270 232.430 171.390 232.710 ;
        RECT 172.230 232.430 183.350 232.710 ;
        RECT 184.190 232.430 195.310 232.710 ;
        RECT 196.150 232.430 207.270 232.710 ;
        RECT 208.110 232.430 219.230 232.710 ;
        RECT 5.680 4.280 219.780 232.430 ;
        RECT 5.680 4.000 6.710 4.280 ;
        RECT 7.550 4.000 20.510 4.280 ;
        RECT 21.350 4.000 34.770 4.280 ;
        RECT 35.610 4.000 49.030 4.280 ;
        RECT 49.870 4.000 62.830 4.280 ;
        RECT 63.670 4.000 77.090 4.280 ;
        RECT 77.930 4.000 91.350 4.280 ;
        RECT 92.190 4.000 105.150 4.280 ;
        RECT 105.990 4.000 119.410 4.280 ;
        RECT 120.250 4.000 133.670 4.280 ;
        RECT 134.510 4.000 147.470 4.280 ;
        RECT 148.310 4.000 161.730 4.280 ;
        RECT 162.570 4.000 175.990 4.280 ;
        RECT 176.830 4.000 189.790 4.280 ;
        RECT 190.630 4.000 204.050 4.280 ;
        RECT 204.890 4.000 218.310 4.280 ;
        RECT 219.150 4.000 219.780 4.280 ;
      LAYER met3 ;
        RECT 4.400 227.440 221.590 228.305 ;
        RECT 4.000 213.200 221.990 227.440 ;
        RECT 4.400 211.840 221.990 213.200 ;
        RECT 4.400 211.800 221.590 211.840 ;
        RECT 4.000 210.440 221.590 211.800 ;
        RECT 4.000 197.560 221.990 210.440 ;
        RECT 4.400 196.160 221.990 197.560 ;
        RECT 4.000 194.840 221.990 196.160 ;
        RECT 4.000 193.440 221.590 194.840 ;
        RECT 4.000 181.920 221.990 193.440 ;
        RECT 4.400 180.520 221.990 181.920 ;
        RECT 4.000 177.840 221.990 180.520 ;
        RECT 4.000 176.440 221.590 177.840 ;
        RECT 4.000 166.280 221.990 176.440 ;
        RECT 4.400 164.880 221.990 166.280 ;
        RECT 4.000 160.840 221.990 164.880 ;
        RECT 4.000 159.440 221.590 160.840 ;
        RECT 4.000 149.960 221.990 159.440 ;
        RECT 4.400 148.560 221.990 149.960 ;
        RECT 4.000 143.840 221.990 148.560 ;
        RECT 4.000 142.440 221.590 143.840 ;
        RECT 4.000 134.320 221.990 142.440 ;
        RECT 4.400 132.920 221.990 134.320 ;
        RECT 4.000 127.520 221.990 132.920 ;
        RECT 4.000 126.120 221.590 127.520 ;
        RECT 4.000 118.680 221.990 126.120 ;
        RECT 4.400 117.280 221.990 118.680 ;
        RECT 4.000 110.520 221.990 117.280 ;
        RECT 4.000 109.120 221.590 110.520 ;
        RECT 4.000 103.040 221.990 109.120 ;
        RECT 4.400 101.640 221.990 103.040 ;
        RECT 4.000 93.520 221.990 101.640 ;
        RECT 4.000 92.120 221.590 93.520 ;
        RECT 4.000 87.400 221.990 92.120 ;
        RECT 4.400 86.000 221.990 87.400 ;
        RECT 4.000 76.520 221.990 86.000 ;
        RECT 4.000 75.120 221.590 76.520 ;
        RECT 4.000 71.080 221.990 75.120 ;
        RECT 4.400 69.680 221.990 71.080 ;
        RECT 4.000 59.520 221.990 69.680 ;
        RECT 4.000 58.120 221.590 59.520 ;
        RECT 4.000 55.440 221.990 58.120 ;
        RECT 4.400 54.040 221.990 55.440 ;
        RECT 4.000 42.520 221.990 54.040 ;
        RECT 4.000 41.120 221.590 42.520 ;
        RECT 4.000 39.800 221.990 41.120 ;
        RECT 4.400 38.400 221.990 39.800 ;
        RECT 4.000 25.520 221.990 38.400 ;
        RECT 4.000 24.160 221.590 25.520 ;
        RECT 4.400 24.120 221.590 24.160 ;
        RECT 4.400 22.760 221.990 24.120 ;
        RECT 4.000 9.200 221.990 22.760 ;
        RECT 4.000 8.520 221.590 9.200 ;
        RECT 4.400 7.800 221.590 8.520 ;
        RECT 4.400 7.120 221.990 7.800 ;
        RECT 4.000 4.255 221.990 7.120 ;
      LAYER met4 ;
        RECT 133.695 10.640 210.385 226.000 ;
  END
END baked_slicel
END LIBRARY

