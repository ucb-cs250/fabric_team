VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_connection_block
  CLASS BLOCK ;
  FOREIGN baked_connection_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 242.560 BY 253.280 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 210.160 242.560 210.760 ;
    END
  END cen
  PIN clb0_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END clb0_cin
  PIN clb0_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END clb0_cout
  PIN clb0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END clb0_input[0]
  PIN clb0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END clb0_input[1]
  PIN clb0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END clb0_input[2]
  PIN clb0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END clb0_input[3]
  PIN clb0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END clb0_input[4]
  PIN clb0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END clb0_input[5]
  PIN clb0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END clb0_input[6]
  PIN clb0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END clb0_input[7]
  PIN clb0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END clb0_input[8]
  PIN clb0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END clb0_input[9]
  PIN clb0_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END clb0_output[0]
  PIN clb0_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END clb0_output[1]
  PIN clb0_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END clb0_output[2]
  PIN clb0_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END clb0_output[3]
  PIN clb0_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END clb0_output[4]
  PIN clb1_cin
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 249.280 6.350 253.280 ;
    END
  END clb1_cin
  PIN clb1_cout
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 249.280 18.770 253.280 ;
    END
  END clb1_cout
  PIN clb1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.370 249.280 31.650 253.280 ;
    END
  END clb1_input[0]
  PIN clb1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 249.280 44.530 253.280 ;
    END
  END clb1_input[1]
  PIN clb1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 249.280 56.950 253.280 ;
    END
  END clb1_input[2]
  PIN clb1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 249.280 69.830 253.280 ;
    END
  END clb1_input[3]
  PIN clb1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 249.280 82.710 253.280 ;
    END
  END clb1_input[4]
  PIN clb1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 249.280 95.590 253.280 ;
    END
  END clb1_input[5]
  PIN clb1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 249.280 108.010 253.280 ;
    END
  END clb1_input[6]
  PIN clb1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 249.280 120.890 253.280 ;
    END
  END clb1_input[7]
  PIN clb1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 249.280 133.770 253.280 ;
    END
  END clb1_input[8]
  PIN clb1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.370 249.280 146.650 253.280 ;
    END
  END clb1_input[9]
  PIN clb1_output[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 249.280 159.070 253.280 ;
    END
  END clb1_output[0]
  PIN clb1_output[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.670 249.280 171.950 253.280 ;
    END
  END clb1_output[1]
  PIN clb1_output[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.550 249.280 184.830 253.280 ;
    END
  END clb1_output[2]
  PIN clb1_output[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.430 249.280 197.710 253.280 ;
    END
  END clb1_output[3]
  PIN clb1_output[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.850 249.280 210.130 253.280 ;
    END
  END clb1_output[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.730 249.280 223.010 253.280 ;
    END
  END clk
  PIN double0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END double0[0]
  PIN double0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END double0[1]
  PIN double0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END double0[2]
  PIN double0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END double0[3]
  PIN double0[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END double0[4]
  PIN double0[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END double0[5]
  PIN double0[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END double0[6]
  PIN double0[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END double0[7]
  PIN double1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 75.520 242.560 76.120 ;
    END
  END double1[0]
  PIN double1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 92.520 242.560 93.120 ;
    END
  END double1[1]
  PIN double1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 108.840 242.560 109.440 ;
    END
  END double1[2]
  PIN double1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 125.840 242.560 126.440 ;
    END
  END double1[3]
  PIN double1[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 142.840 242.560 143.440 ;
    END
  END double1[4]
  PIN double1[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 159.840 242.560 160.440 ;
    END
  END double1[5]
  PIN double1[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 176.840 242.560 177.440 ;
    END
  END double1[6]
  PIN double1[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 193.160 242.560 193.760 ;
    END
  END double1[7]
  PIN global[-1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END global[-1]
  PIN global[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 227.160 242.560 227.760 ;
    END
  END global[0]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 244.160 242.560 244.760 ;
    END
  END rst
  PIN set_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.610 249.280 235.890 253.280 ;
    END
  END set_in
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END shift_in
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END shift_out
  PIN single0[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END single0[0]
  PIN single0[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END single0[1]
  PIN single0[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END single0[2]
  PIN single0[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END single0[3]
  PIN single1[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 8.200 242.560 8.800 ;
    END
  END single1[0]
  PIN single1[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 24.520 242.560 25.120 ;
    END
  END single1[1]
  PIN single1[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 41.520 242.560 42.120 ;
    END
  END single1[2]
  PIN single1[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 238.560 58.520 242.560 59.120 ;
    END
  END single1[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 242.320 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 242.320 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 236.900 242.165 ;
      LAYER met1 ;
        RECT 5.520 10.640 236.900 242.320 ;
      LAYER met2 ;
        RECT 6.630 249.000 18.210 249.280 ;
        RECT 19.050 249.000 31.090 249.280 ;
        RECT 31.930 249.000 43.970 249.280 ;
        RECT 44.810 249.000 56.390 249.280 ;
        RECT 57.230 249.000 69.270 249.280 ;
        RECT 70.110 249.000 82.150 249.280 ;
        RECT 82.990 249.000 95.030 249.280 ;
        RECT 95.870 249.000 107.450 249.280 ;
        RECT 108.290 249.000 120.330 249.280 ;
        RECT 121.170 249.000 133.210 249.280 ;
        RECT 134.050 249.000 146.090 249.280 ;
        RECT 146.930 249.000 158.510 249.280 ;
        RECT 159.350 249.000 171.390 249.280 ;
        RECT 172.230 249.000 184.270 249.280 ;
        RECT 185.110 249.000 197.150 249.280 ;
        RECT 197.990 249.000 209.570 249.280 ;
        RECT 210.410 249.000 222.450 249.280 ;
        RECT 223.290 249.000 235.330 249.280 ;
        RECT 6.080 4.280 235.880 249.000 ;
        RECT 6.630 4.000 18.210 4.280 ;
        RECT 19.050 4.000 31.090 4.280 ;
        RECT 31.930 4.000 43.970 4.280 ;
        RECT 44.810 4.000 56.390 4.280 ;
        RECT 57.230 4.000 69.270 4.280 ;
        RECT 70.110 4.000 82.150 4.280 ;
        RECT 82.990 4.000 95.030 4.280 ;
        RECT 95.870 4.000 107.450 4.280 ;
        RECT 108.290 4.000 120.330 4.280 ;
        RECT 121.170 4.000 133.210 4.280 ;
        RECT 134.050 4.000 146.090 4.280 ;
        RECT 146.930 4.000 158.510 4.280 ;
        RECT 159.350 4.000 171.390 4.280 ;
        RECT 172.230 4.000 184.270 4.280 ;
        RECT 185.110 4.000 197.150 4.280 ;
        RECT 197.990 4.000 209.570 4.280 ;
        RECT 210.410 4.000 222.450 4.280 ;
        RECT 223.290 4.000 235.330 4.280 ;
      LAYER met3 ;
        RECT 4.000 243.800 238.160 244.625 ;
        RECT 4.400 243.760 238.160 243.800 ;
        RECT 4.400 242.400 238.560 243.760 ;
        RECT 4.000 228.160 238.560 242.400 ;
        RECT 4.000 226.760 238.160 228.160 ;
        RECT 4.000 224.080 238.560 226.760 ;
        RECT 4.400 222.680 238.560 224.080 ;
        RECT 4.000 211.160 238.560 222.680 ;
        RECT 4.000 209.760 238.160 211.160 ;
        RECT 4.000 205.040 238.560 209.760 ;
        RECT 4.400 203.640 238.560 205.040 ;
        RECT 4.000 194.160 238.560 203.640 ;
        RECT 4.000 192.760 238.160 194.160 ;
        RECT 4.000 185.320 238.560 192.760 ;
        RECT 4.400 183.920 238.560 185.320 ;
        RECT 4.000 177.840 238.560 183.920 ;
        RECT 4.000 176.440 238.160 177.840 ;
        RECT 4.000 165.600 238.560 176.440 ;
        RECT 4.400 164.200 238.560 165.600 ;
        RECT 4.000 160.840 238.560 164.200 ;
        RECT 4.000 159.440 238.160 160.840 ;
        RECT 4.000 146.560 238.560 159.440 ;
        RECT 4.400 145.160 238.560 146.560 ;
        RECT 4.000 143.840 238.560 145.160 ;
        RECT 4.000 142.440 238.160 143.840 ;
        RECT 4.000 126.840 238.560 142.440 ;
        RECT 4.400 125.440 238.160 126.840 ;
        RECT 4.000 109.840 238.560 125.440 ;
        RECT 4.000 108.440 238.160 109.840 ;
        RECT 4.000 107.800 238.560 108.440 ;
        RECT 4.400 106.400 238.560 107.800 ;
        RECT 4.000 93.520 238.560 106.400 ;
        RECT 4.000 92.120 238.160 93.520 ;
        RECT 4.000 88.080 238.560 92.120 ;
        RECT 4.400 86.680 238.560 88.080 ;
        RECT 4.000 76.520 238.560 86.680 ;
        RECT 4.000 75.120 238.160 76.520 ;
        RECT 4.000 68.360 238.560 75.120 ;
        RECT 4.400 66.960 238.560 68.360 ;
        RECT 4.000 59.520 238.560 66.960 ;
        RECT 4.000 58.120 238.160 59.520 ;
        RECT 4.000 49.320 238.560 58.120 ;
        RECT 4.400 47.920 238.560 49.320 ;
        RECT 4.000 42.520 238.560 47.920 ;
        RECT 4.000 41.120 238.160 42.520 ;
        RECT 4.000 29.600 238.560 41.120 ;
        RECT 4.400 28.200 238.560 29.600 ;
        RECT 4.000 25.520 238.560 28.200 ;
        RECT 4.000 24.120 238.160 25.520 ;
        RECT 4.000 10.560 238.560 24.120 ;
        RECT 4.400 9.200 238.560 10.560 ;
        RECT 4.400 9.160 238.160 9.200 ;
        RECT 4.000 8.335 238.160 9.160 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 242.320 ;
  END
END baked_connection_block
END LIBRARY

