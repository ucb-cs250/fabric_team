module fpga #(
)(
);



/* This FPGA lays out tiles in the following fixed configuration (not to
* scale).
* +-----------++-----------++-----------+
* | clb_tile  ||           || clb_tile  |
* +-----------+| sram_tile |+-----------+
* +-----------+|           |+-----------+
* | clb_tile  ||           || clb_tile  |
* +-----------++-----------++-----------+
* +-----------++-----------++-----------+
* | clb_tile  ||           || clb_tile  |
* +-----------+| mac_tile  |+-----------+
* +-----------+|           |+-----------+
* | clb_tile  ||           || clb_tile  |
* +-----------++-----------++-----------+
* +-----------++-----------++-----------+
* | clb_tile  || clb_tile  || clb_tile  |
* +-----------++-----------++-----------+
* +-----------++-----------++-----------+
* | clb_tile  || clb_tile  || clb_tile  |
* +-----------++-----------++-----------+
*/


mac_tile #(

) mac (

);

endmodule
