magic
tech sky130A
magscale 1 2
timestamp 1608061428
<< locali >>
rect 4077 42551 4111 42721
rect 15025 30583 15059 30753
rect 4169 28543 4203 28713
rect 9045 24599 9079 24837
rect 16681 22967 16715 23137
rect 10517 13855 10551 13957
rect 13001 5015 13035 5321
<< viali >>
rect 11161 47141 11195 47175
rect 9781 47073 9815 47107
rect 9965 47073 9999 47107
rect 11345 47073 11379 47107
rect 12633 47073 12667 47107
rect 12817 47073 12851 47107
rect 14013 47073 14047 47107
rect 14197 47073 14231 47107
rect 15669 47073 15703 47107
rect 15761 47073 15795 47107
rect 13093 47005 13127 47039
rect 16221 47005 16255 47039
rect 10057 46869 10091 46903
rect 11437 46869 11471 46903
rect 14289 46869 14323 46903
rect 15485 46869 15519 46903
rect 10241 46665 10275 46699
rect 15209 46665 15243 46699
rect 13829 46529 13863 46563
rect 5549 46461 5583 46495
rect 8677 46461 8711 46495
rect 8953 46461 8987 46495
rect 11161 46461 11195 46495
rect 12633 46461 12667 46495
rect 14105 46461 14139 46495
rect 16313 46461 16347 46495
rect 16589 46461 16623 46495
rect 5365 46393 5399 46427
rect 12449 46393 12483 46427
rect 16497 46393 16531 46427
rect 17049 46393 17083 46427
rect 5641 46325 5675 46359
rect 11345 46325 11379 46359
rect 12725 46325 12759 46359
rect 6285 46121 6319 46155
rect 8217 46053 8251 46087
rect 12357 46053 12391 46087
rect 13829 46053 13863 46087
rect 17785 46053 17819 46087
rect 8401 45985 8435 46019
rect 10701 45985 10735 46019
rect 13921 45985 13955 46019
rect 16129 45985 16163 46019
rect 16405 45985 16439 46019
rect 4905 45917 4939 45951
rect 5181 45917 5215 45951
rect 10977 45917 11011 45951
rect 8493 45781 8527 45815
rect 13645 45781 13679 45815
rect 14105 45781 14139 45815
rect 5457 45577 5491 45611
rect 8769 45577 8803 45611
rect 13829 45577 13863 45611
rect 16313 45577 16347 45611
rect 11253 45509 11287 45543
rect 9873 45441 9907 45475
rect 12449 45441 12483 45475
rect 18521 45441 18555 45475
rect 4997 45373 5031 45407
rect 5273 45373 5307 45407
rect 6837 45373 6871 45407
rect 7021 45373 7055 45407
rect 8309 45373 8343 45407
rect 8493 45373 8527 45407
rect 8585 45373 8619 45407
rect 10149 45373 10183 45407
rect 12725 45373 12759 45407
rect 14933 45373 14967 45407
rect 15209 45373 15243 45407
rect 18245 45373 18279 45407
rect 5181 45305 5215 45339
rect 18061 45305 18095 45339
rect 7113 45237 7147 45271
rect 7573 45033 7607 45067
rect 4813 44965 4847 44999
rect 9873 44965 9907 44999
rect 11437 44965 11471 44999
rect 11989 44965 12023 44999
rect 13001 44965 13035 44999
rect 13553 44965 13587 44999
rect 17785 44965 17819 44999
rect 4721 44897 4755 44931
rect 4905 44897 4939 44931
rect 5365 44897 5399 44931
rect 6469 44897 6503 44931
rect 9965 44897 9999 44931
rect 11345 44897 11379 44931
rect 11529 44897 11563 44931
rect 13093 44897 13127 44931
rect 16405 44897 16439 44931
rect 6193 44829 6227 44863
rect 9689 44829 9723 44863
rect 16129 44829 16163 44863
rect 10149 44693 10183 44727
rect 12817 44693 12851 44727
rect 5641 44489 5675 44523
rect 9229 44489 9263 44523
rect 10793 44489 10827 44523
rect 15301 44489 15335 44523
rect 10333 44421 10367 44455
rect 7665 44353 7699 44387
rect 14473 44353 14507 44387
rect 3065 44285 3099 44319
rect 4261 44285 4295 44319
rect 4537 44285 4571 44319
rect 7941 44285 7975 44319
rect 10609 44285 10643 44319
rect 12725 44285 12759 44319
rect 13921 44285 13955 44319
rect 14105 44285 14139 44319
rect 15485 44285 15519 44319
rect 15577 44285 15611 44319
rect 16865 44285 16899 44319
rect 2881 44217 2915 44251
rect 3433 44217 3467 44251
rect 10517 44217 10551 44251
rect 12541 44217 12575 44251
rect 16037 44217 16071 44251
rect 12817 44149 12851 44183
rect 17049 44149 17083 44183
rect 6561 43945 6595 43979
rect 4905 43877 4939 43911
rect 11713 43877 11747 43911
rect 17693 43877 17727 43911
rect 4997 43809 5031 43843
rect 6377 43809 6411 43843
rect 7665 43809 7699 43843
rect 7757 43809 7791 43843
rect 10149 43809 10183 43843
rect 10333 43809 10367 43843
rect 11805 43809 11839 43843
rect 13553 43809 13587 43843
rect 13645 43809 13679 43843
rect 16313 43809 16347 43843
rect 11529 43741 11563 43775
rect 12265 43741 12299 43775
rect 14105 43741 14139 43775
rect 16037 43741 16071 43775
rect 4721 43673 4755 43707
rect 5181 43605 5215 43639
rect 7481 43605 7515 43639
rect 7941 43605 7975 43639
rect 10425 43605 10459 43639
rect 13369 43605 13403 43639
rect 10333 43401 10367 43435
rect 14013 43401 14047 43435
rect 18337 43401 18371 43435
rect 12725 43265 12759 43299
rect 15209 43265 15243 43299
rect 3709 43197 3743 43231
rect 5365 43197 5399 43231
rect 5549 43197 5583 43231
rect 7757 43197 7791 43231
rect 8953 43197 8987 43231
rect 9137 43197 9171 43231
rect 10609 43197 10643 43231
rect 12449 43197 12483 43231
rect 14933 43197 14967 43231
rect 18245 43197 18279 43231
rect 3525 43129 3559 43163
rect 5917 43129 5951 43163
rect 7573 43129 7607 43163
rect 9505 43129 9539 43163
rect 10517 43129 10551 43163
rect 11069 43129 11103 43163
rect 18061 43129 18095 43163
rect 3801 43061 3835 43095
rect 7849 43061 7883 43095
rect 16313 43061 16347 43095
rect 13553 42857 13587 42891
rect 4169 42789 4203 42823
rect 8217 42789 8251 42823
rect 1777 42721 1811 42755
rect 2881 42721 2915 42755
rect 4077 42721 4111 42755
rect 4353 42721 4387 42755
rect 8401 42721 8435 42755
rect 9689 42721 9723 42755
rect 12173 42721 12207 42755
rect 12449 42721 12483 42755
rect 15393 42721 15427 42755
rect 15577 42721 15611 42755
rect 18429 42721 18463 42755
rect 1961 42585 1995 42619
rect 4721 42653 4755 42687
rect 5549 42653 5583 42687
rect 5825 42653 5859 42687
rect 6929 42653 6963 42687
rect 9965 42653 9999 42687
rect 11345 42653 11379 42687
rect 15945 42653 15979 42687
rect 16773 42653 16807 42687
rect 17049 42653 17083 42687
rect 3065 42517 3099 42551
rect 4077 42517 4111 42551
rect 8493 42517 8527 42551
rect 4261 42313 4295 42347
rect 5181 42313 5215 42347
rect 5641 42313 5675 42347
rect 9137 42313 9171 42347
rect 18245 42313 18279 42347
rect 14381 42245 14415 42279
rect 15945 42245 15979 42279
rect 2697 42177 2731 42211
rect 7573 42177 7607 42211
rect 11161 42177 11195 42211
rect 13553 42177 13587 42211
rect 15117 42177 15151 42211
rect 2973 42109 3007 42143
rect 5365 42109 5399 42143
rect 5457 42109 5491 42143
rect 7849 42109 7883 42143
rect 10793 42109 10827 42143
rect 11345 42109 11379 42143
rect 13001 42109 13035 42143
rect 13185 42109 13219 42143
rect 14657 42109 14691 42143
rect 16221 42109 16255 42143
rect 18061 42109 18095 42143
rect 14565 42041 14599 42075
rect 16129 42041 16163 42075
rect 16681 42041 16715 42075
rect 5641 41769 5675 41803
rect 15669 41769 15703 41803
rect 7757 41701 7791 41735
rect 9873 41701 9907 41735
rect 18429 41701 18463 41735
rect 2605 41633 2639 41667
rect 2789 41633 2823 41667
rect 7849 41633 7883 41667
rect 9965 41633 9999 41667
rect 11805 41633 11839 41667
rect 12173 41633 12207 41667
rect 13461 41633 13495 41667
rect 13921 41633 13955 41667
rect 14381 41633 14415 41667
rect 15393 41633 15427 41667
rect 15577 41633 15611 41667
rect 17049 41633 17083 41667
rect 3157 41565 3191 41599
rect 4261 41565 4295 41599
rect 4537 41565 4571 41599
rect 7573 41565 7607 41599
rect 11989 41565 12023 41599
rect 14013 41565 14047 41599
rect 16773 41565 16807 41599
rect 9689 41497 9723 41531
rect 8033 41429 8067 41463
rect 10149 41429 10183 41463
rect 13277 41429 13311 41463
rect 3433 41225 3467 41259
rect 4537 41225 4571 41259
rect 8401 41225 8435 41259
rect 9873 41225 9907 41259
rect 12909 41225 12943 41259
rect 5273 41089 5307 41123
rect 11161 41089 11195 41123
rect 14749 41089 14783 41123
rect 2973 41021 3007 41055
rect 3157 41021 3191 41055
rect 3249 41021 3283 41055
rect 4813 41021 4847 41055
rect 7021 41021 7055 41055
rect 7297 41021 7331 41055
rect 9689 41021 9723 41055
rect 10977 41021 11011 41055
rect 11529 41021 11563 41055
rect 13093 41021 13127 41055
rect 13553 41021 13587 41055
rect 14381 41021 14415 41055
rect 14933 41021 14967 41055
rect 16037 41021 16071 41055
rect 16221 41021 16255 41055
rect 4721 40953 4755 40987
rect 16129 40953 16163 40987
rect 16681 40953 16715 40987
rect 3065 40681 3099 40715
rect 18153 40681 18187 40715
rect 6653 40613 6687 40647
rect 7205 40613 7239 40647
rect 15393 40613 15427 40647
rect 15945 40613 15979 40647
rect 1777 40545 1811 40579
rect 2881 40545 2915 40579
rect 4445 40545 4479 40579
rect 4813 40545 4847 40579
rect 5181 40545 5215 40579
rect 6745 40545 6779 40579
rect 8217 40545 8251 40579
rect 8769 40545 8803 40579
rect 9873 40545 9907 40579
rect 11161 40545 11195 40579
rect 11529 40545 11563 40579
rect 12541 40545 12575 40579
rect 15577 40545 15611 40579
rect 17049 40545 17083 40579
rect 6469 40477 6503 40511
rect 8401 40477 8435 40511
rect 12817 40477 12851 40511
rect 16773 40477 16807 40511
rect 1961 40341 1995 40375
rect 10057 40341 10091 40375
rect 11069 40341 11103 40375
rect 13921 40341 13955 40375
rect 4905 40137 4939 40171
rect 7757 40137 7791 40171
rect 9321 40137 9355 40171
rect 12909 40137 12943 40171
rect 15117 40137 15151 40171
rect 18337 40137 18371 40171
rect 3525 40001 3559 40035
rect 11161 40001 11195 40035
rect 13921 40001 13955 40035
rect 2145 39933 2179 39967
rect 2421 39933 2455 39967
rect 4813 39933 4847 39967
rect 5365 39933 5399 39967
rect 6561 39933 6595 39967
rect 7941 39933 7975 39967
rect 8401 39933 8435 39967
rect 9229 39933 9263 39967
rect 9873 39933 9907 39967
rect 10977 39933 11011 39967
rect 11437 39933 11471 39967
rect 13461 39933 13495 39967
rect 13553 39933 13587 39967
rect 13829 39933 13863 39967
rect 14933 39933 14967 39967
rect 16129 39933 16163 39967
rect 16221 39933 16255 39967
rect 16313 39933 16347 39967
rect 18061 39933 18095 39967
rect 18245 39933 18279 39967
rect 16773 39865 16807 39899
rect 6377 39797 6411 39831
rect 12081 39593 12115 39627
rect 18337 39593 18371 39627
rect 6745 39525 6779 39559
rect 2881 39457 2915 39491
rect 4629 39457 4663 39491
rect 4813 39457 4847 39491
rect 5181 39457 5215 39491
rect 6285 39457 6319 39491
rect 6469 39457 6503 39491
rect 7757 39457 7791 39491
rect 8217 39457 8251 39491
rect 8401 39457 8435 39491
rect 8769 39457 8803 39491
rect 10517 39457 10551 39491
rect 13185 39457 13219 39491
rect 13921 39457 13955 39491
rect 14381 39457 14415 39491
rect 15301 39457 15335 39491
rect 15485 39457 15519 39491
rect 17049 39457 17083 39491
rect 10793 39389 10827 39423
rect 14013 39389 14047 39423
rect 16773 39389 16807 39423
rect 13001 39321 13035 39355
rect 3065 39253 3099 39287
rect 7573 39253 7607 39287
rect 15577 39253 15611 39287
rect 2513 39049 2547 39083
rect 3709 39049 3743 39083
rect 11437 39049 11471 39083
rect 2053 38913 2087 38947
rect 5549 38913 5583 38947
rect 7481 38913 7515 38947
rect 10149 38913 10183 38947
rect 12633 38913 12667 38947
rect 15485 38913 15519 38947
rect 2329 38845 2363 38879
rect 3709 38845 3743 38879
rect 4353 38845 4387 38879
rect 5457 38845 5491 38879
rect 5917 38845 5951 38879
rect 7113 38845 7147 38879
rect 7665 38845 7699 38879
rect 8677 38845 8711 38879
rect 9781 38845 9815 38879
rect 10333 38845 10367 38879
rect 11337 38845 11371 38879
rect 12909 38845 12943 38879
rect 15393 38845 15427 38879
rect 15853 38845 15887 38879
rect 16681 38845 16715 38879
rect 2237 38777 2271 38811
rect 8861 38709 8895 38743
rect 14013 38709 14047 38743
rect 16865 38709 16899 38743
rect 4353 38505 4387 38539
rect 8677 38505 8711 38539
rect 9873 38505 9907 38539
rect 12633 38437 12667 38471
rect 16865 38437 16899 38471
rect 2881 38369 2915 38403
rect 4077 38369 4111 38403
rect 4261 38369 4295 38403
rect 5825 38369 5859 38403
rect 6101 38369 6135 38403
rect 7113 38369 7147 38403
rect 7481 38369 7515 38403
rect 7665 38369 7699 38403
rect 8861 38369 8895 38403
rect 9689 38369 9723 38403
rect 10977 38369 11011 38403
rect 13921 38369 13955 38403
rect 14013 38369 14047 38403
rect 14381 38369 14415 38403
rect 15577 38369 15611 38403
rect 15853 38369 15887 38403
rect 17049 38369 17083 38403
rect 11253 38301 11287 38335
rect 15669 38301 15703 38335
rect 3065 38233 3099 38267
rect 5641 38233 5675 38267
rect 17141 38165 17175 38199
rect 3985 37961 4019 37995
rect 5825 37961 5859 37995
rect 6929 37961 6963 37995
rect 10977 37961 11011 37995
rect 11437 37961 11471 37995
rect 13001 37961 13035 37995
rect 8493 37825 8527 37859
rect 13461 37825 13495 37859
rect 18153 37825 18187 37859
rect 2881 37757 2915 37791
rect 3893 37757 3927 37791
rect 4537 37757 4571 37791
rect 5641 37757 5675 37791
rect 6837 37757 6871 37791
rect 7573 37757 7607 37791
rect 8769 37757 8803 37791
rect 11161 37757 11195 37791
rect 11253 37757 11287 37791
rect 13553 37757 13587 37791
rect 13921 37757 13955 37791
rect 14105 37757 14139 37791
rect 14933 37757 14967 37791
rect 16037 37757 16071 37791
rect 16313 37757 16347 37791
rect 18061 37757 18095 37791
rect 2973 37689 3007 37723
rect 16221 37689 16255 37723
rect 16773 37689 16807 37723
rect 10057 37621 10091 37655
rect 15117 37621 15151 37655
rect 6101 37417 6135 37451
rect 12081 37417 12115 37451
rect 15485 37417 15519 37451
rect 2605 37349 2639 37383
rect 8677 37349 8711 37383
rect 11069 37349 11103 37383
rect 14105 37349 14139 37383
rect 18153 37349 18187 37383
rect 2421 37281 2455 37315
rect 2697 37281 2731 37315
rect 4721 37281 4755 37315
rect 4997 37281 5031 37315
rect 7573 37281 7607 37315
rect 7665 37281 7699 37315
rect 8033 37281 8067 37315
rect 8125 37281 8159 37315
rect 9781 37281 9815 37315
rect 9965 37281 9999 37315
rect 10517 37281 10551 37315
rect 10701 37281 10735 37315
rect 12449 37281 12483 37315
rect 12633 37281 12667 37315
rect 13001 37281 13035 37315
rect 13185 37281 13219 37315
rect 14013 37281 14047 37315
rect 15301 37281 15335 37315
rect 16497 37281 16531 37315
rect 16773 37281 16807 37315
rect 2881 37077 2915 37111
rect 4353 36873 4387 36907
rect 5549 36873 5583 36907
rect 7113 36873 7147 36907
rect 8401 36873 8435 36907
rect 10793 36873 10827 36907
rect 12909 36873 12943 36907
rect 16129 36873 16163 36907
rect 3065 36737 3099 36771
rect 6837 36737 6871 36771
rect 9689 36737 9723 36771
rect 15117 36737 15151 36771
rect 2789 36669 2823 36703
rect 5273 36669 5307 36703
rect 5457 36669 5491 36703
rect 6929 36669 6963 36703
rect 8217 36669 8251 36703
rect 9505 36669 9539 36703
rect 9781 36669 9815 36703
rect 10333 36669 10367 36703
rect 10517 36669 10551 36703
rect 11989 36669 12023 36703
rect 12817 36669 12851 36703
rect 14657 36669 14691 36703
rect 14749 36669 14783 36703
rect 15025 36669 15059 36703
rect 16037 36669 16071 36703
rect 16589 36669 16623 36703
rect 12633 36601 12667 36635
rect 14013 36601 14047 36635
rect 9321 36533 9355 36567
rect 11805 36533 11839 36567
rect 10609 36329 10643 36363
rect 15761 36329 15795 36363
rect 3065 36261 3099 36295
rect 4629 36261 4663 36295
rect 2973 36193 3007 36227
rect 5181 36193 5215 36227
rect 5273 36193 5307 36227
rect 5457 36193 5491 36227
rect 5733 36193 5767 36227
rect 6101 36193 6135 36227
rect 10977 36193 11011 36227
rect 11345 36193 11379 36227
rect 13001 36193 13035 36227
rect 13369 36193 13403 36227
rect 13553 36193 13587 36227
rect 15301 36193 15335 36227
rect 15577 36193 15611 36227
rect 16865 36193 16899 36227
rect 17049 36193 17083 36227
rect 7113 36125 7147 36159
rect 7389 36125 7423 36159
rect 10793 36125 10827 36159
rect 11253 36125 11287 36159
rect 13093 36125 13127 36159
rect 15393 36057 15427 36091
rect 8677 35989 8711 36023
rect 12449 35989 12483 36023
rect 17141 35989 17175 36023
rect 10425 35785 10459 35819
rect 16313 35785 16347 35819
rect 3617 35717 3651 35751
rect 9137 35717 9171 35751
rect 12725 35649 12759 35683
rect 13829 35649 13863 35683
rect 15209 35649 15243 35683
rect 3525 35581 3559 35615
rect 4537 35581 4571 35615
rect 4721 35581 4755 35615
rect 5181 35581 5215 35615
rect 5273 35581 5307 35615
rect 6837 35581 6871 35615
rect 8033 35581 8067 35615
rect 8217 35581 8251 35615
rect 8677 35581 8711 35615
rect 8769 35581 8803 35615
rect 10333 35581 10367 35615
rect 11345 35581 11379 35615
rect 12449 35581 12483 35615
rect 14933 35581 14967 35615
rect 18061 35581 18095 35615
rect 18245 35581 18279 35615
rect 5825 35513 5859 35547
rect 7021 35445 7055 35479
rect 11437 35445 11471 35479
rect 18337 35445 18371 35479
rect 15393 35241 15427 35275
rect 14381 35173 14415 35207
rect 18245 35173 18279 35207
rect 4261 35105 4295 35139
rect 4813 35105 4847 35139
rect 5641 35105 5675 35139
rect 8217 35105 8251 35139
rect 9965 35105 9999 35139
rect 12547 35105 12581 35139
rect 13645 35105 13679 35139
rect 15301 35105 15335 35139
rect 5917 35037 5951 35071
rect 8125 35037 8159 35071
rect 10241 35037 10275 35071
rect 14013 35037 14047 35071
rect 16589 35037 16623 35071
rect 16865 35037 16899 35071
rect 13921 34969 13955 35003
rect 4169 34901 4203 34935
rect 7021 34901 7055 34935
rect 8401 34901 8435 34935
rect 11529 34901 11563 34935
rect 12725 34901 12759 34935
rect 13810 34901 13844 34935
rect 2789 34697 2823 34731
rect 10241 34697 10275 34731
rect 12587 34697 12621 34731
rect 12725 34697 12759 34731
rect 18061 34697 18095 34731
rect 18521 34697 18555 34731
rect 14105 34629 14139 34663
rect 3249 34561 3283 34595
rect 5825 34561 5859 34595
rect 6929 34561 6963 34595
rect 12817 34561 12851 34595
rect 12909 34561 12943 34595
rect 15577 34561 15611 34595
rect 3157 34493 3191 34527
rect 3525 34493 3559 34527
rect 3709 34493 3743 34527
rect 4537 34493 4571 34527
rect 4721 34493 4755 34527
rect 5181 34493 5215 34527
rect 5273 34493 5307 34527
rect 7021 34493 7055 34527
rect 7481 34493 7515 34527
rect 7573 34493 7607 34527
rect 9229 34493 9263 34527
rect 9321 34493 9355 34527
rect 9689 34493 9723 34527
rect 9781 34493 9815 34527
rect 11345 34493 11379 34527
rect 11437 34493 11471 34527
rect 14013 34493 14047 34527
rect 15485 34493 15519 34527
rect 15761 34493 15795 34527
rect 18337 34493 18371 34527
rect 19809 34493 19843 34527
rect 12449 34425 12483 34459
rect 18245 34425 18279 34459
rect 19625 34425 19659 34459
rect 8033 34357 8067 34391
rect 19901 34357 19935 34391
rect 2237 34153 2271 34187
rect 4905 34153 4939 34187
rect 8493 34153 8527 34187
rect 9965 34153 9999 34187
rect 11069 34153 11103 34187
rect 13001 34153 13035 34187
rect 18245 34085 18279 34119
rect 2605 34017 2639 34051
rect 2973 34017 3007 34051
rect 3157 34017 3191 34051
rect 4813 34017 4847 34051
rect 6101 34017 6135 34051
rect 8309 34017 8343 34051
rect 9781 34017 9815 34051
rect 11621 34017 11655 34051
rect 11989 34017 12023 34051
rect 12173 34017 12207 34051
rect 13185 34017 13219 34051
rect 13921 34017 13955 34051
rect 14381 34017 14415 34051
rect 16589 34017 16623 34051
rect 2697 33949 2731 33983
rect 5825 33949 5859 33983
rect 11437 33949 11471 33983
rect 14013 33949 14047 33983
rect 16865 33949 16899 33983
rect 7205 33813 7239 33847
rect 8861 33609 8895 33643
rect 14013 33609 14047 33643
rect 16037 33609 16071 33643
rect 2237 33473 2271 33507
rect 4721 33473 4755 33507
rect 5641 33473 5675 33507
rect 7757 33473 7791 33507
rect 16773 33473 16807 33507
rect 2513 33405 2547 33439
rect 5181 33405 5215 33439
rect 5365 33405 5399 33439
rect 5733 33405 5767 33439
rect 7481 33405 7515 33439
rect 10149 33405 10183 33439
rect 10241 33405 10275 33439
rect 10609 33405 10643 33439
rect 10701 33405 10735 33439
rect 12449 33405 12483 33439
rect 12725 33405 12759 33439
rect 14933 33405 14967 33439
rect 16313 33405 16347 33439
rect 16221 33337 16255 33371
rect 3801 33269 3835 33303
rect 11161 33269 11195 33303
rect 15025 33269 15059 33303
rect 2053 33065 2087 33099
rect 3065 33065 3099 33099
rect 4169 33065 4203 33099
rect 7389 33065 7423 33099
rect 8677 33065 8711 33099
rect 12357 33065 12391 33099
rect 13645 32997 13679 33031
rect 1961 32929 1995 32963
rect 2973 32929 3007 32963
rect 4077 32929 4111 32963
rect 5917 32929 5951 32963
rect 8585 32929 8619 32963
rect 9689 32929 9723 32963
rect 9873 32929 9907 32963
rect 11161 32929 11195 32963
rect 11345 32929 11379 32963
rect 11897 32929 11931 32963
rect 12081 32929 12115 32963
rect 13553 32929 13587 32963
rect 15945 32929 15979 32963
rect 16313 32929 16347 32963
rect 16497 32929 16531 32963
rect 6009 32861 6043 32895
rect 6285 32861 6319 32895
rect 14013 32861 14047 32895
rect 14105 32861 14139 32895
rect 15853 32861 15887 32895
rect 13921 32793 13955 32827
rect 5733 32725 5767 32759
rect 9965 32725 9999 32759
rect 13369 32725 13403 32759
rect 13810 32725 13844 32759
rect 15393 32725 15427 32759
rect 3985 32453 4019 32487
rect 6193 32453 6227 32487
rect 7665 32385 7699 32419
rect 9229 32385 9263 32419
rect 9505 32385 9539 32419
rect 10609 32385 10643 32419
rect 13645 32385 13679 32419
rect 13921 32385 13955 32419
rect 1501 32317 1535 32351
rect 2881 32317 2915 32351
rect 3065 32317 3099 32351
rect 3617 32317 3651 32351
rect 3801 32317 3835 32351
rect 5089 32317 5123 32351
rect 6377 32317 6411 32351
rect 7849 32317 7883 32351
rect 8217 32317 8251 32351
rect 8401 32317 8435 32351
rect 12449 32317 12483 32351
rect 16313 32317 16347 32351
rect 16129 32249 16163 32283
rect 16681 32249 16715 32283
rect 1593 32181 1627 32215
rect 5273 32181 5307 32215
rect 7481 32181 7515 32215
rect 12633 32181 12667 32215
rect 15209 32181 15243 32215
rect 4997 31977 5031 32011
rect 7297 31977 7331 32011
rect 8677 31977 8711 32011
rect 13369 31977 13403 32011
rect 16681 31977 16715 32011
rect 3065 31909 3099 31943
rect 9689 31909 9723 31943
rect 1961 31841 1995 31875
rect 2973 31841 3007 31875
rect 4813 31841 4847 31875
rect 5917 31841 5951 31875
rect 8493 31841 8527 31875
rect 9873 31841 9907 31875
rect 11345 31841 11379 31875
rect 11897 31841 11931 31875
rect 12081 31841 12115 31875
rect 13553 31841 13587 31875
rect 13645 31841 13679 31875
rect 14381 31841 14415 31875
rect 17785 31841 17819 31875
rect 6193 31773 6227 31807
rect 10149 31773 10183 31807
rect 11161 31773 11195 31807
rect 14013 31773 14047 31807
rect 15301 31773 15335 31807
rect 15577 31773 15611 31807
rect 13810 31705 13844 31739
rect 13921 31705 13955 31739
rect 2053 31637 2087 31671
rect 12357 31637 12391 31671
rect 17877 31637 17911 31671
rect 11989 31433 12023 31467
rect 14013 31433 14047 31467
rect 15209 31433 15243 31467
rect 1501 31297 1535 31331
rect 1777 31297 1811 31331
rect 4077 31297 4111 31331
rect 9689 31297 9723 31331
rect 12725 31297 12759 31331
rect 16221 31297 16255 31331
rect 4169 31229 4203 31263
rect 4721 31229 4755 31263
rect 4905 31229 4939 31263
rect 7113 31229 7147 31263
rect 8125 31229 8159 31263
rect 8401 31229 8435 31263
rect 10609 31229 10643 31263
rect 10793 31229 10827 31263
rect 12173 31229 12207 31263
rect 12449 31229 12483 31263
rect 15761 31229 15795 31263
rect 15853 31229 15887 31263
rect 16129 31229 16163 31263
rect 2881 31093 2915 31127
rect 5181 31093 5215 31127
rect 7205 31093 7239 31127
rect 10885 31093 10919 31127
rect 3065 30889 3099 30923
rect 6193 30889 6227 30923
rect 10977 30889 11011 30923
rect 15945 30889 15979 30923
rect 7481 30821 7515 30855
rect 11989 30821 12023 30855
rect 1861 30753 1895 30787
rect 2881 30753 2915 30787
rect 5181 30753 5215 30787
rect 5641 30753 5675 30787
rect 5733 30753 5767 30787
rect 7389 30753 7423 30787
rect 7665 30753 7699 30787
rect 9965 30753 9999 30787
rect 10517 30753 10551 30787
rect 10701 30753 10735 30787
rect 12449 30753 12483 30787
rect 12633 30753 12667 30787
rect 13001 30753 13035 30787
rect 13185 30753 13219 30787
rect 14013 30753 14047 30787
rect 15025 30753 15059 30787
rect 15301 30753 15335 30787
rect 16865 30753 16899 30787
rect 4997 30685 5031 30719
rect 9873 30685 9907 30719
rect 1961 30617 1995 30651
rect 15669 30685 15703 30719
rect 16957 30617 16991 30651
rect 7205 30549 7239 30583
rect 7757 30549 7791 30583
rect 14105 30549 14139 30583
rect 15025 30549 15059 30583
rect 15439 30549 15473 30583
rect 15577 30549 15611 30583
rect 10609 30277 10643 30311
rect 12633 30209 12667 30243
rect 13553 30209 13587 30243
rect 15853 30209 15887 30243
rect 16405 30209 16439 30243
rect 1961 30141 1995 30175
rect 3157 30141 3191 30175
rect 3249 30141 3283 30175
rect 3617 30141 3651 30175
rect 3709 30141 3743 30175
rect 5365 30141 5399 30175
rect 5549 30141 5583 30175
rect 6837 30141 6871 30175
rect 8033 30141 8067 30175
rect 8125 30141 8159 30175
rect 8217 30141 8251 30175
rect 10793 30141 10827 30175
rect 10977 30141 11011 30175
rect 11345 30141 11379 30175
rect 11529 30141 11563 30175
rect 13001 30141 13035 30175
rect 13277 30141 13311 30175
rect 15945 30141 15979 30175
rect 16313 30141 16347 30175
rect 2053 30073 2087 30107
rect 5917 30073 5951 30107
rect 8677 30073 8711 30107
rect 15301 30073 15335 30107
rect 4169 30005 4203 30039
rect 6929 30005 6963 30039
rect 4905 29801 4939 29835
rect 7205 29801 7239 29835
rect 9873 29733 9907 29767
rect 1409 29665 1443 29699
rect 1685 29665 1719 29699
rect 4721 29665 4755 29699
rect 5825 29665 5859 29699
rect 8493 29665 8527 29699
rect 9689 29665 9723 29699
rect 9965 29665 9999 29699
rect 11713 29665 11747 29699
rect 12173 29665 12207 29699
rect 12265 29665 12299 29699
rect 13737 29665 13771 29699
rect 13921 29665 13955 29699
rect 15301 29665 15335 29699
rect 15577 29665 15611 29699
rect 6101 29597 6135 29631
rect 11529 29597 11563 29631
rect 2789 29461 2823 29495
rect 8677 29461 8711 29495
rect 10149 29461 10183 29495
rect 12725 29461 12759 29495
rect 14013 29461 14047 29495
rect 16681 29461 16715 29495
rect 8033 29257 8067 29291
rect 15374 29257 15408 29291
rect 18153 29257 18187 29291
rect 4997 29189 5031 29223
rect 9229 29189 9263 29223
rect 15485 29189 15519 29223
rect 16865 29189 16899 29223
rect 3985 29121 4019 29155
rect 13001 29121 13035 29155
rect 15577 29121 15611 29155
rect 1409 29053 1443 29087
rect 1685 29053 1719 29087
rect 4077 29053 4111 29087
rect 4537 29053 4571 29087
rect 4629 29053 4663 29087
rect 6837 29053 6871 29087
rect 7021 29053 7055 29087
rect 7481 29053 7515 29087
rect 7573 29053 7607 29087
rect 9045 29053 9079 29087
rect 10149 29053 10183 29087
rect 10333 29053 10367 29087
rect 10885 29053 10919 29087
rect 11069 29053 11103 29087
rect 12725 29053 12759 29087
rect 15945 29053 15979 29087
rect 16773 29053 16807 29087
rect 18061 29053 18095 29087
rect 14381 28985 14415 29019
rect 15209 28985 15243 29019
rect 2789 28917 2823 28951
rect 11345 28917 11379 28951
rect 3065 28713 3099 28747
rect 4169 28713 4203 28747
rect 17601 28713 17635 28747
rect 1869 28577 1903 28611
rect 2881 28577 2915 28611
rect 4261 28645 4295 28679
rect 11713 28645 11747 28679
rect 5825 28577 5859 28611
rect 8309 28577 8343 28611
rect 10333 28577 10367 28611
rect 12725 28577 12759 28611
rect 13277 28577 13311 28611
rect 13461 28577 13495 28611
rect 16129 28577 16163 28611
rect 16497 28577 16531 28611
rect 17509 28577 17543 28611
rect 4169 28509 4203 28543
rect 4408 28509 4442 28543
rect 4629 28509 4663 28543
rect 6101 28509 6135 28543
rect 10057 28509 10091 28543
rect 12541 28509 12575 28543
rect 16221 28509 16255 28543
rect 16589 28509 16623 28543
rect 1961 28441 1995 28475
rect 4537 28441 4571 28475
rect 4721 28373 4755 28407
rect 7205 28373 7239 28407
rect 8493 28373 8527 28407
rect 13737 28373 13771 28407
rect 15577 28373 15611 28407
rect 2789 28169 2823 28203
rect 11069 28169 11103 28203
rect 12633 28169 12667 28203
rect 18153 28169 18187 28203
rect 9137 28101 9171 28135
rect 4629 28033 4663 28067
rect 5457 28033 5491 28067
rect 10609 28033 10643 28067
rect 13921 28033 13955 28067
rect 1409 27965 1443 27999
rect 1685 27965 1719 27999
rect 4997 27965 5031 27999
rect 5181 27965 5215 27999
rect 5549 27965 5583 27999
rect 7573 27965 7607 27999
rect 7757 27965 7791 27999
rect 8217 27965 8251 27999
rect 9045 27965 9079 27999
rect 9321 27965 9355 27999
rect 10885 27965 10919 27999
rect 12449 27965 12483 27999
rect 13645 27965 13679 27999
rect 16221 27965 16255 27999
rect 16405 27965 16439 27999
rect 16773 27965 16807 27999
rect 18061 27965 18095 27999
rect 7665 27897 7699 27931
rect 10793 27897 10827 27931
rect 15301 27897 15335 27931
rect 9505 27829 9539 27863
rect 1685 27625 1719 27659
rect 7573 27557 7607 27591
rect 10425 27557 10459 27591
rect 13185 27557 13219 27591
rect 1593 27489 1627 27523
rect 2605 27489 2639 27523
rect 2789 27489 2823 27523
rect 4261 27489 4295 27523
rect 4813 27489 4847 27523
rect 4997 27489 5031 27523
rect 6469 27489 6503 27523
rect 6929 27489 6963 27523
rect 7021 27489 7055 27523
rect 8493 27489 8527 27523
rect 9689 27489 9723 27523
rect 9781 27489 9815 27523
rect 9965 27489 9999 27523
rect 11253 27489 11287 27523
rect 11437 27489 11471 27523
rect 13829 27489 13863 27523
rect 14197 27489 14231 27523
rect 14381 27489 14415 27523
rect 15577 27489 15611 27523
rect 17785 27489 17819 27523
rect 3157 27421 3191 27455
rect 4169 27421 4203 27455
rect 6285 27421 6319 27455
rect 13921 27421 13955 27455
rect 15301 27421 15335 27455
rect 16681 27421 16715 27455
rect 5273 27285 5307 27319
rect 8677 27285 8711 27319
rect 11529 27285 11563 27319
rect 17877 27285 17911 27319
rect 10057 27081 10091 27115
rect 11437 27081 11471 27115
rect 15301 27081 15335 27115
rect 16497 27081 16531 27115
rect 12633 27013 12667 27047
rect 2881 26945 2915 26979
rect 3157 26945 3191 26979
rect 5917 26945 5951 26979
rect 13737 26945 13771 26979
rect 1777 26877 1811 26911
rect 5549 26877 5583 26911
rect 6837 26877 6871 26911
rect 8033 26877 8067 26911
rect 8329 26877 8363 26911
rect 8769 26877 8803 26911
rect 9597 26877 9631 26911
rect 9781 26877 9815 26911
rect 9873 26877 9907 26911
rect 11253 26877 11287 26911
rect 12449 26877 12483 26911
rect 14013 26877 14047 26911
rect 16221 26877 16255 26911
rect 16313 26877 16347 26911
rect 18061 26877 18095 26911
rect 5365 26809 5399 26843
rect 8217 26809 8251 26843
rect 1961 26741 1995 26775
rect 4261 26741 4295 26775
rect 7021 26741 7055 26775
rect 18153 26741 18187 26775
rect 6009 26537 6043 26571
rect 8401 26537 8435 26571
rect 14013 26537 14047 26571
rect 4629 26469 4663 26503
rect 10425 26469 10459 26503
rect 12909 26469 12943 26503
rect 2421 26401 2455 26435
rect 2789 26401 2823 26435
rect 4077 26401 4111 26435
rect 4169 26401 4203 26435
rect 6377 26401 6411 26435
rect 6561 26401 6595 26435
rect 6929 26401 6963 26435
rect 7941 26401 7975 26435
rect 8217 26401 8251 26435
rect 9689 26401 9723 26435
rect 9965 26401 9999 26435
rect 11253 26401 11287 26435
rect 13737 26401 13771 26435
rect 13921 26401 13955 26435
rect 15301 26401 15335 26435
rect 2329 26333 2363 26367
rect 2881 26333 2915 26367
rect 6837 26333 6871 26367
rect 11529 26333 11563 26367
rect 16405 26333 16439 26367
rect 16681 26333 16715 26367
rect 8033 26265 8067 26299
rect 9781 26265 9815 26299
rect 1869 26197 1903 26231
rect 15485 26197 15519 26231
rect 17969 26197 18003 26231
rect 8033 25993 8067 26027
rect 10609 25993 10643 26027
rect 13645 25993 13679 26027
rect 1685 25857 1719 25891
rect 3985 25857 4019 25891
rect 4445 25857 4479 25891
rect 7573 25857 7607 25891
rect 10149 25857 10183 25891
rect 14657 25857 14691 25891
rect 15393 25857 15427 25891
rect 1409 25789 1443 25823
rect 4629 25789 4663 25823
rect 4997 25789 5031 25823
rect 5181 25789 5215 25823
rect 7849 25789 7883 25823
rect 9137 25789 9171 25823
rect 10425 25789 10459 25823
rect 12449 25789 12483 25823
rect 12633 25789 12667 25823
rect 13185 25789 13219 25823
rect 13369 25789 13403 25823
rect 15301 25789 15335 25823
rect 15669 25789 15703 25823
rect 15761 25789 15795 25823
rect 16681 25789 16715 25823
rect 3065 25721 3099 25755
rect 7757 25721 7791 25755
rect 10333 25721 10367 25755
rect 9229 25653 9263 25687
rect 16773 25653 16807 25687
rect 5825 25449 5859 25483
rect 9965 25449 9999 25483
rect 12265 25449 12299 25483
rect 1409 25381 1443 25415
rect 7665 25381 7699 25415
rect 13277 25381 13311 25415
rect 17693 25381 17727 25415
rect 2053 25313 2087 25347
rect 2421 25313 2455 25347
rect 4445 25313 4479 25347
rect 7113 25313 7147 25347
rect 7205 25313 7239 25347
rect 8493 25313 8527 25347
rect 9689 25313 9723 25347
rect 9873 25313 9907 25347
rect 11253 25313 11287 25347
rect 11345 25313 11379 25347
rect 11805 25313 11839 25347
rect 11989 25313 12023 25347
rect 13461 25313 13495 25347
rect 16037 25313 16071 25347
rect 2145 25245 2179 25279
rect 2513 25245 2547 25279
rect 4721 25245 4755 25279
rect 16313 25245 16347 25279
rect 6929 25177 6963 25211
rect 8677 25109 8711 25143
rect 13553 25109 13587 25143
rect 4721 24905 4755 24939
rect 9045 24837 9079 24871
rect 10609 24837 10643 24871
rect 16773 24837 16807 24871
rect 2697 24769 2731 24803
rect 7757 24769 7791 24803
rect 2329 24701 2363 24735
rect 3525 24701 3559 24735
rect 3709 24701 3743 24735
rect 4261 24701 4295 24735
rect 4445 24701 4479 24735
rect 5733 24701 5767 24735
rect 7297 24701 7331 24735
rect 7481 24701 7515 24735
rect 2145 24633 2179 24667
rect 11437 24769 11471 24803
rect 10974 24701 11008 24735
rect 11161 24701 11195 24735
rect 12633 24701 12667 24735
rect 14105 24701 14139 24735
rect 14381 24701 14415 24735
rect 16589 24701 16623 24735
rect 18061 24701 18095 24735
rect 19165 24701 19199 24735
rect 9139 24633 9173 24667
rect 12449 24633 12483 24667
rect 15761 24633 15795 24667
rect 19257 24633 19291 24667
rect 5825 24565 5859 24599
rect 9045 24565 9079 24599
rect 12725 24565 12759 24599
rect 18245 24565 18279 24599
rect 1501 24361 1535 24395
rect 8677 24361 8711 24395
rect 16497 24361 16531 24395
rect 6285 24293 6319 24327
rect 9873 24293 9907 24327
rect 10517 24293 10551 24327
rect 13645 24293 13679 24327
rect 17509 24293 17543 24327
rect 1409 24225 1443 24259
rect 2421 24225 2455 24259
rect 2605 24225 2639 24259
rect 7113 24225 7147 24259
rect 7297 24225 7331 24259
rect 8493 24225 8527 24259
rect 9965 24225 9999 24259
rect 10701 24225 10735 24259
rect 11989 24225 12023 24259
rect 15485 24225 15519 24259
rect 16037 24225 16071 24259
rect 16221 24225 16255 24259
rect 18153 24225 18187 24259
rect 18521 24225 18555 24259
rect 19533 24225 19567 24259
rect 4629 24157 4663 24191
rect 4905 24157 4939 24191
rect 12259 24157 12293 24191
rect 15301 24157 15335 24191
rect 18061 24157 18095 24191
rect 18613 24157 18647 24191
rect 2697 24021 2731 24055
rect 7389 24021 7423 24055
rect 9689 24021 9723 24055
rect 10149 24021 10183 24055
rect 10793 24021 10827 24055
rect 19625 24021 19659 24055
rect 8677 23817 8711 23851
rect 10793 23817 10827 23851
rect 14657 23749 14691 23783
rect 18245 23749 18279 23783
rect 19349 23749 19383 23783
rect 4261 23681 4295 23715
rect 5089 23681 5123 23715
rect 10333 23681 10367 23715
rect 13645 23681 13679 23715
rect 15761 23681 15795 23715
rect 16221 23681 16255 23715
rect 2145 23613 2179 23647
rect 2237 23613 2271 23647
rect 2513 23613 2547 23647
rect 2605 23613 2639 23647
rect 4629 23613 4663 23647
rect 4813 23613 4847 23647
rect 5181 23613 5215 23647
rect 6837 23613 6871 23647
rect 7021 23613 7055 23647
rect 7113 23613 7147 23647
rect 8585 23613 8619 23647
rect 10609 23613 10643 23647
rect 12449 23613 12483 23647
rect 13737 23613 13771 23647
rect 14289 23613 14323 23647
rect 14473 23613 14507 23647
rect 16405 23613 16439 23647
rect 16773 23613 16807 23647
rect 16957 23613 16991 23647
rect 18061 23613 18095 23647
rect 19153 23613 19187 23647
rect 20269 23613 20303 23647
rect 1501 23545 1535 23579
rect 7573 23545 7607 23579
rect 8401 23545 8435 23579
rect 10517 23545 10551 23579
rect 12633 23477 12667 23511
rect 20361 23477 20395 23511
rect 2789 23273 2823 23307
rect 8493 23273 8527 23307
rect 12541 23273 12575 23307
rect 13829 23273 13863 23307
rect 15577 23273 15611 23307
rect 18429 23273 18463 23307
rect 5365 23205 5399 23239
rect 9965 23205 9999 23239
rect 15301 23205 15335 23239
rect 17417 23205 17451 23239
rect 1685 23137 1719 23171
rect 4261 23137 4295 23171
rect 4813 23137 4847 23171
rect 4997 23137 5031 23171
rect 7389 23137 7423 23171
rect 10149 23137 10183 23171
rect 11529 23137 11563 23171
rect 11621 23137 11655 23171
rect 11995 23137 12029 23171
rect 12081 23137 12115 23171
rect 13553 23137 13587 23171
rect 13737 23137 13771 23171
rect 15485 23137 15519 23171
rect 16681 23137 16715 23171
rect 16865 23137 16899 23171
rect 16957 23137 16991 23171
rect 18245 23137 18279 23171
rect 19349 23137 19383 23171
rect 1409 23069 1443 23103
rect 4169 23069 4203 23103
rect 7113 23069 7147 23103
rect 10241 22933 10275 22967
rect 16681 22933 16715 22967
rect 19533 22933 19567 22967
rect 1869 22729 1903 22763
rect 2927 22729 2961 22763
rect 8493 22729 8527 22763
rect 19533 22729 19567 22763
rect 3065 22661 3099 22695
rect 3157 22593 3191 22627
rect 4905 22593 4939 22627
rect 10793 22593 10827 22627
rect 15393 22593 15427 22627
rect 16313 22593 16347 22627
rect 18613 22593 18647 22627
rect 1685 22525 1719 22559
rect 2789 22525 2823 22559
rect 5457 22525 5491 22559
rect 5733 22525 5767 22559
rect 5917 22525 5951 22559
rect 6837 22525 6871 22559
rect 7021 22525 7055 22559
rect 8217 22525 8251 22559
rect 8401 22525 8435 22559
rect 9597 22525 9631 22559
rect 10701 22525 10735 22559
rect 10977 22525 11011 22559
rect 13369 22525 13403 22559
rect 13461 22525 13495 22559
rect 13921 22525 13955 22559
rect 14105 22525 14139 22559
rect 15853 22525 15887 22559
rect 16037 22525 16071 22559
rect 16405 22525 16439 22559
rect 18245 22525 18279 22559
rect 19441 22525 19475 22559
rect 18061 22457 18095 22491
rect 3433 22389 3467 22423
rect 7113 22389 7147 22423
rect 9781 22389 9815 22423
rect 11161 22389 11195 22423
rect 14381 22389 14415 22423
rect 13737 22185 13771 22219
rect 6837 22117 6871 22151
rect 10793 22117 10827 22151
rect 1777 22049 1811 22083
rect 2881 22049 2915 22083
rect 4905 22049 4939 22083
rect 5273 22049 5307 22083
rect 7021 22049 7055 22083
rect 8217 22049 8251 22083
rect 8401 22049 8435 22083
rect 10609 22049 10643 22083
rect 10885 22049 10919 22083
rect 11345 22049 11379 22083
rect 12449 22049 12483 22083
rect 17877 22049 17911 22083
rect 18705 22049 18739 22083
rect 19801 22049 19835 22083
rect 4445 21981 4479 22015
rect 7297 21981 7331 22015
rect 8769 21981 8803 22015
rect 12173 21981 12207 22015
rect 16221 21981 16255 22015
rect 16497 21981 16531 22015
rect 19901 21981 19935 22015
rect 1961 21913 1995 21947
rect 5181 21913 5215 21947
rect 3065 21845 3099 21879
rect 18889 21845 18923 21879
rect 8401 21641 8435 21675
rect 11437 21641 11471 21675
rect 14197 21641 14231 21675
rect 16313 21641 16347 21675
rect 12449 21573 12483 21607
rect 5365 21505 5399 21539
rect 9965 21505 9999 21539
rect 13185 21505 13219 21539
rect 15117 21505 15151 21539
rect 18613 21505 18647 21539
rect 2053 21437 2087 21471
rect 3157 21437 3191 21471
rect 3341 21437 3375 21471
rect 3893 21437 3927 21471
rect 4077 21437 4111 21471
rect 5457 21437 5491 21471
rect 6837 21437 6871 21471
rect 7941 21437 7975 21471
rect 8217 21437 8251 21471
rect 9505 21437 9539 21471
rect 9597 21437 9631 21471
rect 9781 21437 9815 21471
rect 11259 21437 11293 21471
rect 12725 21437 12759 21471
rect 14013 21437 14047 21471
rect 15301 21437 15335 21471
rect 15853 21437 15887 21471
rect 16037 21437 16071 21471
rect 18705 21437 18739 21471
rect 19073 21437 19107 21471
rect 19165 21437 19199 21471
rect 20085 21437 20119 21471
rect 5917 21369 5951 21403
rect 8125 21369 8159 21403
rect 12633 21369 12667 21403
rect 18061 21369 18095 21403
rect 2237 21301 2271 21335
rect 4353 21301 4387 21335
rect 7021 21301 7055 21335
rect 20177 21301 20211 21335
rect 3065 21029 3099 21063
rect 6561 21029 6595 21063
rect 9873 21029 9907 21063
rect 10425 21029 10459 21063
rect 15853 21029 15887 21063
rect 4353 20961 4387 20995
rect 5733 20961 5767 20995
rect 7113 20961 7147 20995
rect 7297 20961 7331 20995
rect 7389 20961 7423 20995
rect 7941 20961 7975 20995
rect 9689 20961 9723 20995
rect 9965 20961 9999 20995
rect 11253 20961 11287 20995
rect 12449 20961 12483 20995
rect 13001 20961 13035 20995
rect 13185 20961 13219 20995
rect 15301 20961 15335 20995
rect 15485 20961 15519 20995
rect 17049 20961 17083 20995
rect 19257 20961 19291 20995
rect 1409 20893 1443 20927
rect 1685 20893 1719 20927
rect 4077 20893 4111 20927
rect 7665 20893 7699 20927
rect 12357 20893 12391 20927
rect 16773 20893 16807 20927
rect 18245 20893 18279 20927
rect 13369 20825 13403 20859
rect 11345 20757 11379 20791
rect 19349 20757 19383 20791
rect 1685 20553 1719 20587
rect 10149 20553 10183 20587
rect 11437 20553 11471 20587
rect 18337 20553 18371 20587
rect 5365 20485 5399 20519
rect 8769 20485 8803 20519
rect 9689 20485 9723 20519
rect 15669 20417 15703 20451
rect 16589 20417 16623 20451
rect 18208 20417 18242 20451
rect 18429 20417 18463 20451
rect 2237 20349 2271 20383
rect 2329 20349 2363 20383
rect 2605 20349 2639 20383
rect 2697 20349 2731 20383
rect 4721 20349 4755 20383
rect 4905 20349 4939 20383
rect 5457 20349 5491 20383
rect 7021 20349 7055 20383
rect 7113 20349 7147 20383
rect 8585 20349 8619 20383
rect 9965 20349 9999 20383
rect 11253 20349 11287 20383
rect 13185 20349 13219 20383
rect 13461 20349 13495 20383
rect 16129 20349 16163 20383
rect 16313 20349 16347 20383
rect 16681 20349 16715 20383
rect 19625 20349 19659 20383
rect 6837 20281 6871 20315
rect 7205 20281 7239 20315
rect 7573 20281 7607 20315
rect 9873 20281 9907 20315
rect 14841 20281 14875 20315
rect 18061 20281 18095 20315
rect 19717 20281 19751 20315
rect 18705 20213 18739 20247
rect 1501 20009 1535 20043
rect 6837 20009 6871 20043
rect 8493 20009 8527 20043
rect 14105 20009 14139 20043
rect 15485 20009 15519 20043
rect 18889 19941 18923 19975
rect 1409 19873 1443 19907
rect 2421 19873 2455 19907
rect 4353 19873 4387 19907
rect 5733 19873 5767 19907
rect 8033 19873 8067 19907
rect 8309 19873 8343 19907
rect 9689 19873 9723 19907
rect 9873 19873 9907 19907
rect 11345 19873 11379 19907
rect 11621 19873 11655 19907
rect 13829 19873 13863 19907
rect 14013 19873 14047 19907
rect 15301 19873 15335 19907
rect 17417 19873 17451 19907
rect 17509 19873 17543 19907
rect 17785 19873 17819 19907
rect 17969 19873 18003 19907
rect 18797 19873 18831 19907
rect 2568 19805 2602 19839
rect 2789 19805 2823 19839
rect 5457 19805 5491 19839
rect 2881 19737 2915 19771
rect 8125 19737 8159 19771
rect 2697 19669 2731 19703
rect 4537 19669 4571 19703
rect 9965 19669 9999 19703
rect 12725 19669 12759 19703
rect 16865 19669 16899 19703
rect 2973 19465 3007 19499
rect 4721 19465 4755 19499
rect 6469 19465 6503 19499
rect 7941 19465 7975 19499
rect 8401 19465 8435 19499
rect 9597 19465 9631 19499
rect 14381 19465 14415 19499
rect 18337 19465 18371 19499
rect 2835 19397 2869 19431
rect 4537 19397 4571 19431
rect 10517 19397 10551 19431
rect 3065 19329 3099 19363
rect 4629 19329 4663 19363
rect 16129 19329 16163 19363
rect 18208 19329 18242 19363
rect 18429 19329 18463 19363
rect 1685 19261 1719 19295
rect 1777 19261 1811 19295
rect 2697 19261 2731 19295
rect 4408 19261 4442 19295
rect 6653 19261 6687 19295
rect 6837 19261 6871 19295
rect 8217 19261 8251 19295
rect 9497 19261 9531 19295
rect 10793 19261 10827 19295
rect 13369 19261 13403 19295
rect 13461 19261 13495 19295
rect 13921 19261 13955 19295
rect 14105 19261 14139 19295
rect 15393 19261 15427 19295
rect 16037 19261 16071 19295
rect 16405 19261 16439 19295
rect 16497 19261 16531 19295
rect 3433 19193 3467 19227
rect 4261 19193 4295 19227
rect 8125 19193 8159 19227
rect 10701 19193 10735 19227
rect 11253 19193 11287 19227
rect 18061 19193 18095 19227
rect 7021 19125 7055 19159
rect 18705 19125 18739 19159
rect 2789 18921 2823 18955
rect 8493 18921 8527 18955
rect 9965 18921 9999 18955
rect 11989 18921 12023 18955
rect 15485 18921 15519 18955
rect 19165 18921 19199 18955
rect 4261 18785 4295 18819
rect 4721 18785 4755 18819
rect 4813 18785 4847 18819
rect 6929 18785 6963 18819
rect 7297 18785 7331 18819
rect 8309 18785 8343 18819
rect 10333 18785 10367 18819
rect 10701 18785 10735 18819
rect 10793 18785 10827 18819
rect 11713 18785 11747 18819
rect 11897 18785 11931 18819
rect 13829 18785 13863 18819
rect 14197 18785 14231 18819
rect 14381 18785 14415 18819
rect 15301 18785 15335 18819
rect 16865 18785 16899 18819
rect 19073 18785 19107 18819
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 4169 18717 4203 18751
rect 6285 18717 6319 18751
rect 7021 18717 7055 18751
rect 7205 18717 7239 18751
rect 10425 18717 10459 18751
rect 13921 18717 13955 18751
rect 16589 18717 16623 18751
rect 5273 18581 5307 18615
rect 13461 18581 13495 18615
rect 17969 18581 18003 18615
rect 9873 18377 9907 18411
rect 19533 18377 19567 18411
rect 10885 18309 10919 18343
rect 2421 18241 2455 18275
rect 3525 18241 3559 18275
rect 11253 18241 11287 18275
rect 18613 18241 18647 18275
rect 2053 18173 2087 18207
rect 3249 18173 3283 18207
rect 5733 18173 5767 18207
rect 7021 18173 7055 18207
rect 7389 18173 7423 18207
rect 8309 18173 8343 18207
rect 8585 18173 8619 18207
rect 10793 18173 10827 18207
rect 11069 18173 11103 18207
rect 12817 18173 12851 18207
rect 12909 18173 12943 18207
rect 13369 18173 13403 18207
rect 13553 18173 13587 18207
rect 15485 18173 15519 18207
rect 15761 18173 15795 18207
rect 18061 18173 18095 18207
rect 18245 18173 18279 18207
rect 19441 18173 19475 18207
rect 1869 18105 1903 18139
rect 6837 18105 6871 18139
rect 17141 18105 17175 18139
rect 4629 18037 4663 18071
rect 5825 18037 5859 18071
rect 13829 18037 13863 18071
rect 4445 17833 4479 17867
rect 7021 17833 7055 17867
rect 16497 17833 16531 17867
rect 1593 17765 1627 17799
rect 18705 17765 18739 17799
rect 2237 17697 2271 17731
rect 2329 17697 2363 17731
rect 2605 17697 2639 17731
rect 2789 17697 2823 17731
rect 3893 17697 3927 17731
rect 4353 17697 4387 17731
rect 8125 17697 8159 17731
rect 8217 17697 8251 17731
rect 10793 17697 10827 17731
rect 10885 17697 10919 17731
rect 12449 17697 12483 17731
rect 15485 17697 15519 17731
rect 16037 17697 16071 17731
rect 16221 17697 16255 17731
rect 17509 17697 17543 17731
rect 18613 17697 18647 17731
rect 5457 17629 5491 17663
rect 5733 17629 5767 17663
rect 7941 17629 7975 17663
rect 10609 17629 10643 17663
rect 12180 17629 12214 17663
rect 15301 17629 15335 17663
rect 13737 17561 13771 17595
rect 3709 17493 3743 17527
rect 8401 17493 8435 17527
rect 11069 17493 11103 17527
rect 17693 17493 17727 17527
rect 1685 17289 1719 17323
rect 11069 17289 11103 17323
rect 12725 17289 12759 17323
rect 17049 17289 17083 17323
rect 2697 17221 2731 17255
rect 4261 17221 4295 17255
rect 3065 17153 3099 17187
rect 5733 17153 5767 17187
rect 7757 17153 7791 17187
rect 8677 17153 8711 17187
rect 14657 17153 14691 17187
rect 1593 17085 1627 17119
rect 2605 17085 2639 17119
rect 2881 17085 2915 17119
rect 4169 17085 4203 17119
rect 5457 17085 5491 17119
rect 5641 17085 5675 17119
rect 7389 17085 7423 17119
rect 8769 17085 8803 17119
rect 9321 17085 9355 17119
rect 9505 17085 9539 17119
rect 10793 17085 10827 17119
rect 10977 17085 11011 17119
rect 12633 17085 12667 17119
rect 14013 17085 14047 17119
rect 14841 17085 14875 17119
rect 15393 17085 15427 17119
rect 15577 17085 15611 17119
rect 16865 17085 16899 17119
rect 18061 17085 18095 17119
rect 19165 17085 19199 17119
rect 7205 17017 7239 17051
rect 9873 17017 9907 17051
rect 12449 17017 12483 17051
rect 15945 17017 15979 17051
rect 13829 16949 13863 16983
rect 18245 16949 18279 16983
rect 19257 16949 19291 16983
rect 6469 16745 6503 16779
rect 9965 16745 9999 16779
rect 19349 16745 19383 16779
rect 11713 16677 11747 16711
rect 1409 16609 1443 16643
rect 4261 16609 4295 16643
rect 4353 16609 4387 16643
rect 4721 16609 4755 16643
rect 4813 16609 4847 16643
rect 6285 16609 6319 16643
rect 7573 16609 7607 16643
rect 8125 16609 8159 16643
rect 8309 16609 8343 16643
rect 10149 16609 10183 16643
rect 10333 16609 10367 16643
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 11897 16609 11931 16643
rect 13093 16609 13127 16643
rect 13277 16609 13311 16643
rect 14657 16609 14691 16643
rect 15761 16609 15795 16643
rect 16037 16609 16071 16643
rect 18245 16609 18279 16643
rect 19257 16609 19291 16643
rect 1685 16541 1719 16575
rect 3065 16541 3099 16575
rect 7389 16541 7423 16575
rect 8585 16541 8619 16575
rect 18337 16541 18371 16575
rect 14473 16473 14507 16507
rect 5273 16405 5307 16439
rect 11989 16405 12023 16439
rect 13369 16405 13403 16439
rect 17325 16405 17359 16439
rect 6193 16201 6227 16235
rect 8493 16201 8527 16235
rect 11253 16201 11287 16235
rect 17049 16201 17083 16235
rect 18337 16201 18371 16235
rect 18705 16201 18739 16235
rect 2421 16133 2455 16167
rect 3985 16065 4019 16099
rect 5089 16065 5123 16099
rect 7389 16065 7423 16099
rect 9965 16065 9999 16099
rect 12449 16065 12483 16099
rect 15025 16065 15059 16099
rect 18208 16065 18242 16099
rect 18429 16065 18463 16099
rect 2292 15997 2326 16031
rect 2484 15997 2518 16031
rect 3709 15997 3743 16031
rect 6377 15997 6411 16031
rect 7021 15997 7055 16031
rect 8217 15997 8251 16031
rect 8401 15997 8435 16031
rect 9689 15997 9723 16031
rect 12725 15997 12759 16031
rect 15393 15997 15427 16031
rect 15577 15997 15611 16031
rect 15945 15997 15979 16031
rect 16129 15997 16163 16031
rect 16957 15997 16991 16031
rect 18061 15997 18095 16031
rect 2145 15929 2179 15963
rect 2881 15929 2915 15963
rect 6837 15929 6871 15963
rect 14105 15929 14139 15963
rect 9781 15657 9815 15691
rect 13461 15657 13495 15691
rect 17969 15657 18003 15691
rect 1593 15589 1627 15623
rect 4721 15589 4755 15623
rect 6745 15589 6779 15623
rect 15301 15589 15335 15623
rect 18981 15589 19015 15623
rect 2237 15521 2271 15555
rect 2605 15521 2639 15555
rect 2789 15521 2823 15555
rect 5549 15521 5583 15555
rect 7389 15521 7423 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 9137 15521 9171 15555
rect 9689 15521 9723 15555
rect 10701 15521 10735 15555
rect 13829 15521 13863 15555
rect 14197 15521 14231 15555
rect 14381 15521 14415 15555
rect 15945 15521 15979 15555
rect 16313 15521 16347 15555
rect 17325 15521 17359 15555
rect 18889 15521 18923 15555
rect 2329 15453 2363 15487
rect 5273 15453 5307 15487
rect 5733 15453 5767 15487
rect 7481 15453 7515 15487
rect 10977 15453 11011 15487
rect 13921 15453 13955 15487
rect 15761 15453 15795 15487
rect 16221 15453 16255 15487
rect 17693 15453 17727 15487
rect 17490 15385 17524 15419
rect 8953 15317 8987 15351
rect 12265 15317 12299 15351
rect 17601 15317 17635 15351
rect 19165 15113 19199 15147
rect 9597 15045 9631 15079
rect 13553 15045 13587 15079
rect 16957 15045 16991 15079
rect 2237 14977 2271 15011
rect 3157 14977 3191 15011
rect 14657 14977 14691 15011
rect 1869 14909 1903 14943
rect 3249 14909 3283 14943
rect 3709 14909 3743 14943
rect 3801 14909 3835 14943
rect 5273 14909 5307 14943
rect 5457 14909 5491 14943
rect 6837 14909 6871 14943
rect 7113 14909 7147 14943
rect 9781 14909 9815 14943
rect 9965 14909 9999 14943
rect 10333 14909 10367 14943
rect 10517 14909 10551 14943
rect 11345 14909 11379 14943
rect 12587 14909 12621 14943
rect 12725 14909 12759 14943
rect 13185 14909 13219 14943
rect 13369 14909 13403 14943
rect 14841 14909 14875 14943
rect 15393 14909 15427 14943
rect 15577 14909 15611 14943
rect 16865 14909 16899 14943
rect 18061 14909 18095 14943
rect 19073 14909 19107 14943
rect 1685 14841 1719 14875
rect 8493 14841 8527 14875
rect 4261 14773 4295 14807
rect 5549 14773 5583 14807
rect 11437 14773 11471 14807
rect 15853 14773 15887 14807
rect 18153 14773 18187 14807
rect 15853 14569 15887 14603
rect 8585 14501 8619 14535
rect 2145 14433 2179 14467
rect 2513 14433 2547 14467
rect 7481 14433 7515 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 9689 14433 9723 14467
rect 11253 14433 11287 14467
rect 11483 14433 11517 14467
rect 11621 14433 11655 14467
rect 12081 14433 12115 14467
rect 12265 14433 12299 14467
rect 13553 14433 13587 14467
rect 15761 14433 15795 14467
rect 2237 14365 2271 14399
rect 2605 14365 2639 14399
rect 4813 14365 4847 14399
rect 5089 14365 5123 14399
rect 7297 14365 7331 14399
rect 12541 14365 12575 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 11069 14297 11103 14331
rect 1593 14229 1627 14263
rect 6193 14229 6227 14263
rect 9873 14229 9907 14263
rect 13645 14229 13679 14263
rect 18153 14229 18187 14263
rect 2053 14025 2087 14059
rect 7113 14025 7147 14059
rect 10609 14025 10643 14059
rect 11437 14025 11471 14059
rect 12725 14025 12759 14059
rect 19165 14025 19199 14059
rect 5825 13957 5859 13991
rect 10517 13957 10551 13991
rect 13829 13957 13863 13991
rect 18153 13957 18187 13991
rect 2973 13889 3007 13923
rect 3249 13889 3283 13923
rect 4353 13889 4387 13923
rect 6837 13889 6871 13923
rect 15577 13889 15611 13923
rect 1869 13821 1903 13855
rect 5641 13821 5675 13855
rect 6929 13821 6963 13855
rect 8309 13821 8343 13855
rect 8493 13821 8527 13855
rect 9045 13821 9079 13855
rect 9229 13821 9263 13855
rect 10517 13821 10551 13855
rect 10793 13821 10827 13855
rect 11253 13821 11287 13855
rect 12541 13821 12575 13855
rect 13645 13821 13679 13855
rect 15301 13821 15335 13855
rect 16957 13821 16991 13855
rect 18061 13821 18095 13855
rect 19073 13821 19107 13855
rect 9597 13753 9631 13787
rect 2789 13481 2823 13515
rect 6101 13481 6135 13515
rect 4629 13413 4663 13447
rect 5181 13413 5215 13447
rect 11345 13413 11379 13447
rect 15301 13413 15335 13447
rect 16957 13413 16991 13447
rect 1685 13345 1719 13379
rect 4721 13345 4755 13379
rect 6653 13345 6687 13379
rect 6992 13345 7026 13379
rect 7205 13345 7239 13379
rect 8033 13345 8067 13379
rect 9965 13345 9999 13379
rect 12173 13345 12207 13379
rect 15448 13345 15482 13379
rect 17601 13345 17635 13379
rect 17693 13345 17727 13379
rect 17969 13345 18003 13379
rect 18153 13345 18187 13379
rect 1409 13277 1443 13311
rect 4445 13277 4479 13311
rect 6469 13277 6503 13311
rect 8401 13277 8435 13311
rect 9689 13277 9723 13311
rect 12449 13277 12483 13311
rect 15669 13277 15703 13311
rect 13737 13209 13771 13243
rect 8171 13141 8205 13175
rect 8309 13141 8343 13175
rect 8677 13141 8711 13175
rect 15577 13141 15611 13175
rect 15761 13141 15795 13175
rect 6469 12937 6503 12971
rect 7021 12937 7055 12971
rect 11437 12937 11471 12971
rect 14381 12869 14415 12903
rect 18153 12869 18187 12903
rect 3341 12801 3375 12835
rect 4169 12801 4203 12835
rect 4721 12801 4755 12835
rect 5181 12801 5215 12835
rect 8493 12801 8527 12835
rect 8861 12801 8895 12835
rect 15669 12801 15703 12835
rect 19165 12801 19199 12835
rect 1409 12733 1443 12767
rect 1593 12733 1627 12767
rect 2973 12733 3007 12767
rect 4997 12733 5031 12767
rect 6653 12733 6687 12767
rect 6837 12733 6871 12767
rect 9045 12733 9079 12767
rect 9413 12733 9447 12767
rect 9597 12733 9631 12767
rect 11253 12733 11287 12767
rect 13001 12733 13035 12767
rect 13277 12733 13311 12767
rect 16037 12733 16071 12767
rect 16313 12733 16347 12767
rect 16589 12733 16623 12767
rect 18061 12733 18095 12767
rect 19073 12733 19107 12767
rect 1961 12665 1995 12699
rect 2789 12665 2823 12699
rect 1501 12393 1535 12427
rect 4261 12393 4295 12427
rect 13737 12393 13771 12427
rect 2421 12325 2455 12359
rect 5365 12325 5399 12359
rect 19073 12325 19107 12359
rect 1409 12257 1443 12291
rect 2605 12257 2639 12291
rect 4077 12257 4111 12291
rect 6009 12257 6043 12291
rect 6377 12257 6411 12291
rect 7573 12257 7607 12291
rect 8125 12257 8159 12291
rect 8309 12257 8343 12291
rect 10333 12257 10367 12291
rect 10885 12257 10919 12291
rect 11253 12257 11287 12291
rect 12449 12257 12483 12291
rect 12725 12257 12759 12291
rect 13277 12257 13311 12291
rect 13461 12257 13495 12291
rect 15853 12257 15887 12291
rect 17601 12257 17635 12291
rect 17969 12257 18003 12291
rect 18981 12257 19015 12291
rect 5825 12189 5859 12223
rect 6285 12189 6319 12223
rect 7481 12189 7515 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 17509 12189 17543 12223
rect 18061 12189 18095 12223
rect 8493 12121 8527 12155
rect 16037 12121 16071 12155
rect 2697 12053 2731 12087
rect 12265 12053 12299 12087
rect 17049 12053 17083 12087
rect 10977 11849 11011 11883
rect 11161 11849 11195 11883
rect 19717 11849 19751 11883
rect 4353 11781 4387 11815
rect 16497 11781 16531 11815
rect 2605 11713 2639 11747
rect 8217 11713 8251 11747
rect 8493 11713 8527 11747
rect 10848 11713 10882 11747
rect 11069 11713 11103 11747
rect 15577 11713 15611 11747
rect 2145 11645 2179 11679
rect 2237 11645 2271 11679
rect 2513 11645 2547 11679
rect 4629 11645 4663 11679
rect 6469 11645 6503 11679
rect 6837 11645 6871 11679
rect 9873 11645 9907 11679
rect 12449 11645 12483 11679
rect 13921 11645 13955 11679
rect 14197 11645 14231 11679
rect 16405 11645 16439 11679
rect 16681 11645 16715 11679
rect 18245 11645 18279 11679
rect 19625 11645 19659 11679
rect 1501 11577 1535 11611
rect 4537 11577 4571 11611
rect 5089 11577 5123 11611
rect 10701 11577 10735 11611
rect 17141 11577 17175 11611
rect 18061 11577 18095 11611
rect 18613 11577 18647 11611
rect 19441 11577 19475 11611
rect 6285 11509 6319 11543
rect 7021 11509 7055 11543
rect 12633 11509 12667 11543
rect 2789 11305 2823 11339
rect 6745 11305 6779 11339
rect 9781 11305 9815 11339
rect 19165 11305 19199 11339
rect 16957 11237 16991 11271
rect 1685 11169 1719 11203
rect 4629 11169 4663 11203
rect 4905 11169 4939 11203
rect 7297 11169 7331 11203
rect 7665 11169 7699 11203
rect 7849 11169 7883 11203
rect 9689 11169 9723 11203
rect 13277 11169 13311 11203
rect 13461 11169 13495 11203
rect 15577 11169 15611 11203
rect 18061 11169 18095 11203
rect 1409 11101 1443 11135
rect 4077 11101 4111 11135
rect 5089 11101 5123 11135
rect 7389 11101 7423 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 13737 11101 13771 11135
rect 15301 11101 15335 11135
rect 17785 11101 17819 11135
rect 12173 11033 12207 11067
rect 5457 10761 5491 10795
rect 6929 10761 6963 10795
rect 10425 10761 10459 10795
rect 15485 10761 15519 10795
rect 14381 10693 14415 10727
rect 4169 10625 4203 10659
rect 11069 10625 11103 10659
rect 13185 10625 13219 10659
rect 2605 10557 2639 10591
rect 2881 10557 2915 10591
rect 3893 10557 3927 10591
rect 6561 10557 6595 10591
rect 6837 10557 6871 10591
rect 7849 10557 7883 10591
rect 8033 10557 8067 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 10977 10557 11011 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 13369 10557 13403 10591
rect 13921 10557 13955 10591
rect 14105 10557 14139 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 16405 10557 16439 10591
rect 16497 10557 16531 10591
rect 18061 10557 18095 10591
rect 19165 10557 19199 10591
rect 20177 10557 20211 10591
rect 19257 10489 19291 10523
rect 20269 10489 20303 10523
rect 2605 10421 2639 10455
rect 6377 10421 6411 10455
rect 9045 10421 9079 10455
rect 18245 10421 18279 10455
rect 19165 10217 19199 10251
rect 7021 10149 7055 10183
rect 16497 10149 16531 10183
rect 17233 10149 17267 10183
rect 2605 10081 2639 10115
rect 2973 10081 3007 10115
rect 3157 10081 3191 10115
rect 4077 10081 4111 10115
rect 5365 10081 5399 10115
rect 7849 10081 7883 10115
rect 9689 10081 9723 10115
rect 9965 10081 9999 10115
rect 12725 10081 12759 10115
rect 13185 10081 13219 10115
rect 13737 10081 13771 10115
rect 13921 10081 13955 10115
rect 15307 10081 15341 10115
rect 16644 10081 16678 10115
rect 18061 10081 18095 10115
rect 19073 10081 19107 10115
rect 20913 10081 20947 10115
rect 2697 10013 2731 10047
rect 5641 10013 5675 10047
rect 13001 10013 13035 10047
rect 16865 10013 16899 10047
rect 2053 9945 2087 9979
rect 4261 9945 4295 9979
rect 16773 9945 16807 9979
rect 8033 9877 8067 9911
rect 11253 9877 11287 9911
rect 12541 9877 12575 9911
rect 14197 9877 14231 9911
rect 15485 9877 15519 9911
rect 18153 9877 18187 9911
rect 21005 9877 21039 9911
rect 5733 9673 5767 9707
rect 3433 9605 3467 9639
rect 4629 9537 4663 9571
rect 8769 9537 8803 9571
rect 9965 9537 9999 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 1869 9469 1903 9503
rect 2145 9469 2179 9503
rect 4721 9469 4755 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 7619 9469 7653 9503
rect 7757 9469 7791 9503
rect 8125 9469 8159 9503
rect 8217 9469 8251 9503
rect 9689 9469 9723 9503
rect 12449 9469 12483 9503
rect 13645 9469 13679 9503
rect 14197 9469 14231 9503
rect 14381 9469 14415 9503
rect 16209 9469 16243 9503
rect 18061 9469 18095 9503
rect 19073 9469 19107 9503
rect 20085 9469 20119 9503
rect 1777 9401 1811 9435
rect 19165 9401 19199 9435
rect 11253 9333 11287 9367
rect 16405 9333 16439 9367
rect 18153 9333 18187 9367
rect 20177 9333 20211 9367
rect 1501 9129 1535 9163
rect 19625 9129 19659 9163
rect 3157 9061 3191 9095
rect 5641 9061 5675 9095
rect 8217 9061 8251 9095
rect 9781 9061 9815 9095
rect 14289 9061 14323 9095
rect 1409 8993 1443 9027
rect 2421 8993 2455 9027
rect 2697 8993 2731 9027
rect 4537 8993 4571 9027
rect 5089 8993 5123 9027
rect 5273 8993 5307 9027
rect 6837 8993 6871 9027
rect 9697 8993 9731 9027
rect 10885 8993 10919 9027
rect 11253 8993 11287 9027
rect 12909 8993 12943 9027
rect 13737 8993 13771 9027
rect 13921 8993 13955 9027
rect 18521 8993 18555 9027
rect 19533 8993 19567 9027
rect 4445 8925 4479 8959
rect 6561 8925 6595 8959
rect 11529 8925 11563 8959
rect 16037 8925 16071 8959
rect 16313 8925 16347 8959
rect 17417 8925 17451 8959
rect 2513 8857 2547 8891
rect 10701 8789 10735 8823
rect 18613 8789 18647 8823
rect 4353 8585 4387 8619
rect 16957 8585 16991 8619
rect 19165 8585 19199 8619
rect 5641 8517 5675 8551
rect 10977 8517 11011 8551
rect 12890 8517 12924 8551
rect 13001 8517 13035 8551
rect 15945 8517 15979 8551
rect 3893 8449 3927 8483
rect 11069 8449 11103 8483
rect 14657 8449 14691 8483
rect 2513 8381 2547 8415
rect 2789 8381 2823 8415
rect 2973 8381 3007 8415
rect 4077 8381 4111 8415
rect 4169 8381 4203 8415
rect 5457 8381 5491 8415
rect 6837 8381 6871 8415
rect 8401 8381 8435 8415
rect 8585 8381 8619 8415
rect 9137 8381 9171 8415
rect 9321 8381 9355 8415
rect 10701 8381 10735 8415
rect 10848 8381 10882 8415
rect 13064 8381 13098 8415
rect 13461 8381 13495 8415
rect 14381 8381 14415 8415
rect 16865 8381 16899 8415
rect 18061 8381 18095 8415
rect 19073 8381 19107 8415
rect 1961 8313 1995 8347
rect 12725 8313 12759 8347
rect 7021 8245 7055 8279
rect 9597 8245 9631 8279
rect 11345 8245 11379 8279
rect 18153 8245 18187 8279
rect 4261 8041 4295 8075
rect 11253 8041 11287 8075
rect 15393 8041 15427 8075
rect 6101 7973 6135 8007
rect 12173 7973 12207 8007
rect 16313 7973 16347 8007
rect 1685 7905 1719 7939
rect 4077 7905 4111 7939
rect 5549 7905 5583 7939
rect 5641 7905 5675 7939
rect 7113 7905 7147 7939
rect 7389 7905 7423 7939
rect 7941 7905 7975 7939
rect 8125 7905 8159 7939
rect 9965 7905 9999 7939
rect 12817 7905 12851 7939
rect 13185 7905 13219 7939
rect 14197 7905 14231 7939
rect 14289 7905 14323 7939
rect 15301 7905 15335 7939
rect 16957 7905 16991 7939
rect 17325 7905 17359 7939
rect 17509 7905 17543 7939
rect 18337 7905 18371 7939
rect 1409 7837 1443 7871
rect 5365 7837 5399 7871
rect 7205 7837 7239 7871
rect 9689 7837 9723 7871
rect 12909 7837 12943 7871
rect 13277 7837 13311 7871
rect 17049 7837 17083 7871
rect 8309 7769 8343 7803
rect 2973 7701 3007 7735
rect 6929 7701 6963 7735
rect 18429 7701 18463 7735
rect 7021 7497 7055 7531
rect 11069 7429 11103 7463
rect 12587 7429 12621 7463
rect 12725 7429 12759 7463
rect 16865 7429 16899 7463
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 10940 7361 10974 7395
rect 12817 7361 12851 7395
rect 14565 7361 14599 7395
rect 2243 7293 2277 7327
rect 3617 7293 3651 7327
rect 3893 7293 3927 7327
rect 4905 7293 4939 7327
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 11132 7293 11166 7327
rect 11529 7293 11563 7327
rect 14289 7293 14323 7327
rect 16773 7293 16807 7327
rect 18061 7293 18095 7327
rect 5089 7225 5123 7259
rect 10793 7225 10827 7259
rect 12449 7225 12483 7259
rect 2421 7157 2455 7191
rect 3433 7157 3467 7191
rect 9597 7157 9631 7191
rect 13093 7157 13127 7191
rect 15853 7157 15887 7191
rect 18153 7157 18187 7191
rect 17601 6953 17635 6987
rect 4445 6885 4479 6919
rect 4813 6885 4847 6919
rect 11897 6885 11931 6919
rect 2697 6817 2731 6851
rect 4261 6817 4295 6851
rect 4353 6817 4387 6851
rect 5641 6817 5675 6851
rect 6745 6817 6779 6851
rect 9873 6817 9907 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 15945 6817 15979 6851
rect 16313 6817 16347 6851
rect 16497 6817 16531 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 1869 6749 1903 6783
rect 2421 6749 2455 6783
rect 2881 6749 2915 6783
rect 4077 6749 4111 6783
rect 7021 6749 7055 6783
rect 9781 6749 9815 6783
rect 10333 6749 10367 6783
rect 12725 6749 12759 6783
rect 13001 6749 13035 6783
rect 16037 6749 16071 6783
rect 8309 6681 8343 6715
rect 11253 6681 11287 6715
rect 5825 6613 5859 6647
rect 14105 6613 14139 6647
rect 15393 6613 15427 6647
rect 13001 6409 13035 6443
rect 16589 6409 16623 6443
rect 2973 6341 3007 6375
rect 7941 6341 7975 6375
rect 1685 6273 1719 6307
rect 4353 6273 4387 6307
rect 6929 6273 6963 6307
rect 10149 6273 10183 6307
rect 13461 6273 13495 6307
rect 14013 6273 14047 6307
rect 15025 6273 15059 6307
rect 15301 6273 15335 6307
rect 1409 6205 1443 6239
rect 4537 6205 4571 6239
rect 4905 6205 4939 6239
rect 5089 6205 5123 6239
rect 7021 6205 7055 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 10241 6205 10275 6239
rect 10609 6205 10643 6239
rect 10793 6205 10827 6239
rect 13553 6205 13587 6239
rect 13921 6205 13955 6239
rect 18061 6205 18095 6239
rect 9597 6137 9631 6171
rect 4169 6069 4203 6103
rect 18153 6069 18187 6103
rect 3065 5865 3099 5899
rect 4261 5865 4295 5899
rect 4445 5797 4479 5831
rect 4813 5797 4847 5831
rect 5825 5797 5859 5831
rect 6377 5797 6411 5831
rect 11345 5797 11379 5831
rect 16405 5797 16439 5831
rect 1501 5729 1535 5763
rect 2881 5729 2915 5763
rect 4353 5729 4387 5763
rect 5917 5729 5951 5763
rect 7389 5729 7423 5763
rect 7481 5729 7515 5763
rect 7941 5729 7975 5763
rect 9965 5729 9999 5763
rect 13645 5729 13679 5763
rect 14013 5729 14047 5763
rect 14197 5729 14231 5763
rect 15301 5729 15335 5763
rect 15393 5729 15427 5763
rect 16313 5729 16347 5763
rect 4077 5661 4111 5695
rect 9689 5661 9723 5695
rect 13553 5661 13587 5695
rect 7205 5593 7239 5627
rect 1593 5525 1627 5559
rect 5641 5525 5675 5559
rect 13093 5525 13127 5559
rect 3433 5321 3467 5355
rect 7021 5321 7055 5355
rect 13001 5321 13035 5355
rect 15669 5321 15703 5355
rect 2237 5253 2271 5287
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 5917 5185 5951 5219
rect 9137 5185 9171 5219
rect 11069 5185 11103 5219
rect 2041 5117 2075 5151
rect 3801 5117 3835 5151
rect 4169 5117 4203 5151
rect 5181 5117 5215 5151
rect 5365 5117 5399 5151
rect 5457 5117 5491 5151
rect 6837 5117 6871 5151
rect 8769 5117 8803 5151
rect 10609 5117 10643 5151
rect 10701 5117 10735 5151
rect 10977 5117 11011 5151
rect 8585 5049 8619 5083
rect 9965 5049 9999 5083
rect 14473 5253 14507 5287
rect 13369 5185 13403 5219
rect 13093 5117 13127 5151
rect 15577 5117 15611 5151
rect 13001 4981 13035 5015
rect 9873 4777 9907 4811
rect 12357 4777 12391 4811
rect 15577 4777 15611 4811
rect 4721 4709 4755 4743
rect 5273 4709 5307 4743
rect 13461 4709 13495 4743
rect 15301 4709 15335 4743
rect 2973 4641 3007 4675
rect 3157 4641 3191 4675
rect 4813 4641 4847 4675
rect 6653 4641 6687 4675
rect 6837 4641 6871 4675
rect 7389 4641 7423 4675
rect 7573 4641 7607 4675
rect 9689 4641 9723 4675
rect 13645 4641 13679 4675
rect 15485 4641 15519 4675
rect 23029 4641 23063 4675
rect 2145 4573 2179 4607
rect 2697 4573 2731 4607
rect 4537 4573 4571 4607
rect 10977 4573 11011 4607
rect 11253 4573 11287 4607
rect 14013 4573 14047 4607
rect 23397 4573 23431 4607
rect 23194 4505 23228 4539
rect 7849 4437 7883 4471
rect 23305 4437 23339 4471
rect 23489 4437 23523 4471
rect 3433 4233 3467 4267
rect 18613 4233 18647 4267
rect 22293 4165 22327 4199
rect 2145 4097 2179 4131
rect 7573 4097 7607 4131
rect 7849 4097 7883 4131
rect 9229 4097 9263 4131
rect 12449 4097 12483 4131
rect 13001 4097 13035 4131
rect 14620 4097 14654 4131
rect 14841 4097 14875 4131
rect 15117 4097 15151 4131
rect 22164 4097 22198 4131
rect 22385 4097 22419 4131
rect 22477 4097 22511 4131
rect 1869 4029 1903 4063
rect 4721 4029 4755 4063
rect 4813 4029 4847 4063
rect 5273 4029 5307 4063
rect 5457 4029 5491 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 10793 4029 10827 4063
rect 10977 4029 11011 4063
rect 13093 4029 13127 4063
rect 13461 4029 13495 4063
rect 13645 4029 13679 4063
rect 14703 4029 14737 4063
rect 16037 4029 16071 4063
rect 18521 4029 18555 4063
rect 14473 3961 14507 3995
rect 18337 3961 18371 3995
rect 22017 3961 22051 3995
rect 5733 3893 5767 3927
rect 11253 3893 11287 3927
rect 16129 3893 16163 3927
rect 4537 3689 4571 3723
rect 8125 3689 8159 3723
rect 11253 3689 11287 3723
rect 14289 3689 14323 3723
rect 22845 3689 22879 3723
rect 7113 3621 7147 3655
rect 22201 3621 22235 3655
rect 2697 3553 2731 3587
rect 2973 3553 3007 3587
rect 3157 3553 3191 3587
rect 4353 3553 4387 3587
rect 5733 3553 5767 3587
rect 7941 3553 7975 3587
rect 9965 3553 9999 3587
rect 12817 3553 12851 3587
rect 12909 3553 12943 3587
rect 13185 3553 13219 3587
rect 14197 3553 14231 3587
rect 15301 3553 15335 3587
rect 16681 3553 16715 3587
rect 18245 3553 18279 3587
rect 2145 3485 2179 3519
rect 5457 3485 5491 3519
rect 9689 3485 9723 3519
rect 13277 3485 13311 3519
rect 17049 3485 17083 3519
rect 18392 3485 18426 3519
rect 18613 3485 18647 3519
rect 22569 3485 22603 3519
rect 16846 3417 16880 3451
rect 22477 3417 22511 3451
rect 12265 3349 12299 3383
rect 15393 3349 15427 3383
rect 16957 3349 16991 3383
rect 17325 3349 17359 3383
rect 18521 3349 18555 3383
rect 18705 3349 18739 3383
rect 22366 3349 22400 3383
rect 4077 3145 4111 3179
rect 5181 3145 5215 3179
rect 10057 3145 10091 3179
rect 15098 3145 15132 3179
rect 19349 3145 19383 3179
rect 21557 3145 21591 3179
rect 13829 3077 13863 3111
rect 15209 3077 15243 3111
rect 19238 3077 19272 3111
rect 21189 3077 21223 3111
rect 2973 3009 3007 3043
rect 5917 3009 5951 3043
rect 9137 3009 9171 3043
rect 12725 3009 12759 3043
rect 15301 3009 15335 3043
rect 15393 3009 15427 3043
rect 19441 3009 19475 3043
rect 21281 3009 21315 3043
rect 1501 2941 1535 2975
rect 2697 2941 2731 2975
rect 5457 2941 5491 2975
rect 7481 2941 7515 2975
rect 7757 2941 7791 2975
rect 9965 2941 9999 2975
rect 10977 2941 11011 2975
rect 12449 2941 12483 2975
rect 21060 2941 21094 2975
rect 22569 2941 22603 2975
rect 5365 2873 5399 2907
rect 14933 2873 14967 2907
rect 19073 2873 19107 2907
rect 20913 2873 20947 2907
rect 1593 2805 1627 2839
rect 11069 2805 11103 2839
rect 19717 2805 19751 2839
rect 22661 2805 22695 2839
rect 8125 2601 8159 2635
rect 11253 2601 11287 2635
rect 12725 2601 12759 2635
rect 15577 2601 15611 2635
rect 18981 2601 19015 2635
rect 23029 2601 23063 2635
rect 1869 2533 1903 2567
rect 4445 2533 4479 2567
rect 13829 2533 13863 2567
rect 18337 2533 18371 2567
rect 22385 2533 22419 2567
rect 2016 2465 2050 2499
rect 4261 2465 4295 2499
rect 4537 2465 4571 2499
rect 5825 2465 5859 2499
rect 7113 2465 7147 2499
rect 7665 2465 7699 2499
rect 7849 2465 7883 2499
rect 9873 2465 9907 2499
rect 10149 2465 10183 2499
rect 12633 2465 12667 2499
rect 13976 2465 14010 2499
rect 15485 2465 15519 2499
rect 18484 2465 18518 2499
rect 21373 2465 21407 2499
rect 22532 2465 22566 2499
rect 2237 2397 2271 2431
rect 5917 2397 5951 2431
rect 6929 2397 6963 2431
rect 14197 2397 14231 2431
rect 18705 2397 18739 2431
rect 22753 2397 22787 2431
rect 2145 2329 2179 2363
rect 14105 2329 14139 2363
rect 21465 2329 21499 2363
rect 22661 2329 22695 2363
rect 2513 2261 2547 2295
rect 4721 2261 4755 2295
rect 14289 2261 14323 2295
rect 18613 2261 18647 2295
<< metal1 >>
rect 22094 49104 22100 49156
rect 22152 49144 22158 49156
rect 23198 49144 23204 49156
rect 22152 49116 23204 49144
rect 22152 49104 22158 49116
rect 23198 49104 23204 49116
rect 23256 49104 23262 49156
rect 1104 47354 24840 47376
rect 1104 47302 8912 47354
rect 8964 47302 8976 47354
rect 9028 47302 9040 47354
rect 9092 47302 9104 47354
rect 9156 47302 16843 47354
rect 16895 47302 16907 47354
rect 16959 47302 16971 47354
rect 17023 47302 17035 47354
rect 17087 47302 24840 47354
rect 1104 47280 24840 47302
rect 11238 47240 11244 47252
rect 9968 47212 11244 47240
rect 8202 47064 8208 47116
rect 8260 47104 8266 47116
rect 9968 47113 9996 47212
rect 11238 47200 11244 47212
rect 11296 47240 11302 47252
rect 12158 47240 12164 47252
rect 11296 47212 12164 47240
rect 11296 47200 11302 47212
rect 12158 47200 12164 47212
rect 12216 47200 12222 47252
rect 21174 47200 21180 47252
rect 21232 47240 21238 47252
rect 21634 47240 21640 47252
rect 21232 47212 21640 47240
rect 21232 47200 21238 47212
rect 21634 47200 21640 47212
rect 21692 47200 21698 47252
rect 11149 47175 11207 47181
rect 11149 47141 11161 47175
rect 11195 47172 11207 47175
rect 13814 47172 13820 47184
rect 11195 47144 12572 47172
rect 11195 47141 11207 47144
rect 11149 47135 11207 47141
rect 12544 47116 12572 47144
rect 12820 47144 13820 47172
rect 9769 47107 9827 47113
rect 9769 47104 9781 47107
rect 8260 47076 9781 47104
rect 8260 47064 8266 47076
rect 9769 47073 9781 47076
rect 9815 47073 9827 47107
rect 9769 47067 9827 47073
rect 9953 47107 10011 47113
rect 9953 47073 9965 47107
rect 9999 47073 10011 47107
rect 9953 47067 10011 47073
rect 11333 47107 11391 47113
rect 11333 47073 11345 47107
rect 11379 47104 11391 47107
rect 11379 47076 12388 47104
rect 11379 47073 11391 47076
rect 11333 47067 11391 47073
rect 3050 46928 3056 46980
rect 3108 46968 3114 46980
rect 6270 46968 6276 46980
rect 3108 46940 6276 46968
rect 3108 46928 3114 46940
rect 6270 46928 6276 46940
rect 6328 46928 6334 46980
rect 12360 46912 12388 47076
rect 12526 47064 12532 47116
rect 12584 47104 12590 47116
rect 12820 47113 12848 47144
rect 13814 47132 13820 47144
rect 13872 47172 13878 47184
rect 14550 47172 14556 47184
rect 13872 47144 14556 47172
rect 13872 47132 13878 47144
rect 14550 47132 14556 47144
rect 14608 47132 14614 47184
rect 12621 47107 12679 47113
rect 12621 47104 12633 47107
rect 12584 47076 12633 47104
rect 12584 47064 12590 47076
rect 12621 47073 12633 47076
rect 12667 47073 12679 47107
rect 12621 47067 12679 47073
rect 12805 47107 12863 47113
rect 12805 47073 12817 47107
rect 12851 47073 12863 47107
rect 13998 47104 14004 47116
rect 13959 47076 14004 47104
rect 12805 47067 12863 47073
rect 13998 47064 14004 47076
rect 14056 47064 14062 47116
rect 14182 47104 14188 47116
rect 14143 47076 14188 47104
rect 14182 47064 14188 47076
rect 14240 47064 14246 47116
rect 15654 47104 15660 47116
rect 15615 47076 15660 47104
rect 15654 47064 15660 47076
rect 15712 47064 15718 47116
rect 15746 47064 15752 47116
rect 15804 47104 15810 47116
rect 15804 47076 15849 47104
rect 15804 47064 15810 47076
rect 12434 46996 12440 47048
rect 12492 47036 12498 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12492 47008 13093 47036
rect 12492 46996 12498 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 16206 47036 16212 47048
rect 16167 47008 16212 47036
rect 13081 46999 13139 47005
rect 16206 46996 16212 47008
rect 16264 46996 16270 47048
rect 2682 46860 2688 46912
rect 2740 46900 2746 46912
rect 3326 46900 3332 46912
rect 2740 46872 3332 46900
rect 2740 46860 2746 46872
rect 3326 46860 3332 46872
rect 3384 46860 3390 46912
rect 10042 46900 10048 46912
rect 10003 46872 10048 46900
rect 10042 46860 10048 46872
rect 10100 46860 10106 46912
rect 11422 46900 11428 46912
rect 11383 46872 11428 46900
rect 11422 46860 11428 46872
rect 11480 46860 11486 46912
rect 12342 46900 12348 46912
rect 12255 46872 12348 46900
rect 12342 46860 12348 46872
rect 12400 46900 12406 46912
rect 13722 46900 13728 46912
rect 12400 46872 13728 46900
rect 12400 46860 12406 46872
rect 13722 46860 13728 46872
rect 13780 46860 13786 46912
rect 14274 46900 14280 46912
rect 14235 46872 14280 46900
rect 14274 46860 14280 46872
rect 14332 46860 14338 46912
rect 15470 46900 15476 46912
rect 15431 46872 15476 46900
rect 15470 46860 15476 46872
rect 15528 46860 15534 46912
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 24026 46900 24032 46912
rect 20036 46872 24032 46900
rect 20036 46860 20042 46872
rect 24026 46860 24032 46872
rect 24084 46860 24090 46912
rect 1104 46810 24840 46832
rect 1104 46758 4947 46810
rect 4999 46758 5011 46810
rect 5063 46758 5075 46810
rect 5127 46758 5139 46810
rect 5191 46758 12878 46810
rect 12930 46758 12942 46810
rect 12994 46758 13006 46810
rect 13058 46758 13070 46810
rect 13122 46758 20808 46810
rect 20860 46758 20872 46810
rect 20924 46758 20936 46810
rect 20988 46758 21000 46810
rect 21052 46758 24840 46810
rect 1104 46736 24840 46758
rect 1946 46656 1952 46708
rect 2004 46696 2010 46708
rect 4338 46696 4344 46708
rect 2004 46668 4344 46696
rect 2004 46656 2010 46668
rect 4338 46656 4344 46668
rect 4396 46656 4402 46708
rect 10229 46699 10287 46705
rect 10229 46665 10241 46699
rect 10275 46696 10287 46699
rect 10594 46696 10600 46708
rect 10275 46668 10600 46696
rect 10275 46665 10287 46668
rect 10229 46659 10287 46665
rect 10594 46656 10600 46668
rect 10652 46656 10658 46708
rect 14182 46656 14188 46708
rect 14240 46696 14246 46708
rect 15197 46699 15255 46705
rect 15197 46696 15209 46699
rect 14240 46668 15209 46696
rect 14240 46656 14246 46668
rect 15197 46665 15209 46668
rect 15243 46696 15255 46699
rect 17678 46696 17684 46708
rect 15243 46668 17684 46696
rect 15243 46665 15255 46668
rect 15197 46659 15255 46665
rect 17678 46656 17684 46668
rect 17736 46656 17742 46708
rect 18414 46656 18420 46708
rect 18472 46696 18478 46708
rect 25590 46696 25596 46708
rect 18472 46668 25596 46696
rect 18472 46656 18478 46668
rect 25590 46656 25596 46668
rect 25648 46656 25654 46708
rect 1118 46588 1124 46640
rect 1176 46628 1182 46640
rect 5718 46628 5724 46640
rect 1176 46600 5724 46628
rect 1176 46588 1182 46600
rect 5718 46588 5724 46600
rect 5776 46588 5782 46640
rect 13817 46563 13875 46569
rect 13817 46529 13829 46563
rect 13863 46560 13875 46563
rect 14826 46560 14832 46572
rect 13863 46532 14832 46560
rect 13863 46529 13875 46532
rect 13817 46523 13875 46529
rect 14826 46520 14832 46532
rect 14884 46520 14890 46572
rect 5537 46495 5595 46501
rect 5537 46461 5549 46495
rect 5583 46492 5595 46495
rect 5902 46492 5908 46504
rect 5583 46464 5908 46492
rect 5583 46461 5595 46464
rect 5537 46455 5595 46461
rect 5902 46452 5908 46464
rect 5960 46452 5966 46504
rect 7650 46452 7656 46504
rect 7708 46492 7714 46504
rect 8665 46495 8723 46501
rect 8665 46492 8677 46495
rect 7708 46464 8677 46492
rect 7708 46452 7714 46464
rect 8665 46461 8677 46464
rect 8711 46461 8723 46495
rect 8665 46455 8723 46461
rect 8754 46452 8760 46504
rect 8812 46492 8818 46504
rect 8941 46495 8999 46501
rect 8941 46492 8953 46495
rect 8812 46464 8953 46492
rect 8812 46452 8818 46464
rect 8941 46461 8953 46464
rect 8987 46461 8999 46495
rect 11146 46492 11152 46504
rect 11107 46464 11152 46492
rect 8941 46455 8999 46461
rect 11146 46452 11152 46464
rect 11204 46452 11210 46504
rect 12621 46495 12679 46501
rect 12621 46461 12633 46495
rect 12667 46492 12679 46495
rect 14090 46492 14096 46504
rect 12667 46464 13952 46492
rect 14051 46464 14096 46492
rect 12667 46461 12679 46464
rect 12621 46455 12679 46461
rect 5353 46427 5411 46433
rect 5353 46393 5365 46427
rect 5399 46424 5411 46427
rect 5442 46424 5448 46436
rect 5399 46396 5448 46424
rect 5399 46393 5411 46396
rect 5353 46387 5411 46393
rect 5442 46384 5448 46396
rect 5500 46384 5506 46436
rect 12437 46427 12495 46433
rect 12437 46393 12449 46427
rect 12483 46424 12495 46427
rect 12526 46424 12532 46436
rect 12483 46396 12532 46424
rect 12483 46393 12495 46396
rect 12437 46387 12495 46393
rect 12526 46384 12532 46396
rect 12584 46424 12590 46436
rect 13170 46424 13176 46436
rect 12584 46396 13176 46424
rect 12584 46384 12590 46396
rect 13170 46384 13176 46396
rect 13228 46384 13234 46436
rect 5626 46356 5632 46368
rect 5587 46328 5632 46356
rect 5626 46316 5632 46328
rect 5684 46316 5690 46368
rect 11330 46356 11336 46368
rect 11291 46328 11336 46356
rect 11330 46316 11336 46328
rect 11388 46316 11394 46368
rect 12710 46356 12716 46368
rect 12671 46328 12716 46356
rect 12710 46316 12716 46328
rect 12768 46316 12774 46368
rect 13924 46356 13952 46464
rect 14090 46452 14096 46464
rect 14148 46452 14154 46504
rect 15470 46452 15476 46504
rect 15528 46492 15534 46504
rect 16301 46495 16359 46501
rect 16301 46492 16313 46495
rect 15528 46464 16313 46492
rect 15528 46452 15534 46464
rect 16301 46461 16313 46464
rect 16347 46461 16359 46495
rect 16301 46455 16359 46461
rect 16577 46495 16635 46501
rect 16577 46461 16589 46495
rect 16623 46492 16635 46495
rect 17126 46492 17132 46504
rect 16623 46464 17132 46492
rect 16623 46461 16635 46464
rect 16577 46455 16635 46461
rect 17126 46452 17132 46464
rect 17184 46452 17190 46504
rect 15378 46384 15384 46436
rect 15436 46424 15442 46436
rect 16485 46427 16543 46433
rect 16485 46424 16497 46427
rect 15436 46396 16497 46424
rect 15436 46384 15442 46396
rect 16485 46393 16497 46396
rect 16531 46393 16543 46427
rect 16485 46387 16543 46393
rect 16666 46384 16672 46436
rect 16724 46424 16730 46436
rect 17037 46427 17095 46433
rect 17037 46424 17049 46427
rect 16724 46396 17049 46424
rect 16724 46384 16730 46396
rect 17037 46393 17049 46396
rect 17083 46393 17095 46427
rect 17037 46387 17095 46393
rect 17954 46384 17960 46436
rect 18012 46424 18018 46436
rect 20070 46424 20076 46436
rect 18012 46396 20076 46424
rect 18012 46384 18018 46396
rect 20070 46384 20076 46396
rect 20128 46384 20134 46436
rect 21358 46384 21364 46436
rect 21416 46424 21422 46436
rect 24762 46424 24768 46436
rect 21416 46396 24768 46424
rect 21416 46384 21422 46396
rect 24762 46384 24768 46396
rect 24820 46384 24826 46436
rect 16114 46356 16120 46368
rect 13924 46328 16120 46356
rect 16114 46316 16120 46328
rect 16172 46316 16178 46368
rect 1104 46266 24840 46288
rect 1104 46214 8912 46266
rect 8964 46214 8976 46266
rect 9028 46214 9040 46266
rect 9092 46214 9104 46266
rect 9156 46214 16843 46266
rect 16895 46214 16907 46266
rect 16959 46214 16971 46266
rect 17023 46214 17035 46266
rect 17087 46214 24840 46266
rect 1104 46192 24840 46214
rect 5902 46112 5908 46164
rect 5960 46152 5966 46164
rect 6273 46155 6331 46161
rect 6273 46152 6285 46155
rect 5960 46124 6285 46152
rect 5960 46112 5966 46124
rect 6273 46121 6285 46124
rect 6319 46121 6331 46155
rect 6273 46115 6331 46121
rect 18506 46112 18512 46164
rect 18564 46152 18570 46164
rect 22462 46152 22468 46164
rect 18564 46124 22468 46152
rect 18564 46112 18570 46124
rect 22462 46112 22468 46124
rect 22520 46112 22526 46164
rect 8202 46084 8208 46096
rect 8163 46056 8208 46084
rect 8202 46044 8208 46056
rect 8260 46044 8266 46096
rect 12342 46084 12348 46096
rect 12303 46056 12348 46084
rect 12342 46044 12348 46056
rect 12400 46044 12406 46096
rect 13817 46087 13875 46093
rect 13817 46053 13829 46087
rect 13863 46084 13875 46087
rect 14274 46084 14280 46096
rect 13863 46056 14280 46084
rect 13863 46053 13875 46056
rect 13817 46047 13875 46053
rect 14274 46044 14280 46056
rect 14332 46044 14338 46096
rect 17773 46087 17831 46093
rect 17773 46053 17785 46087
rect 17819 46084 17831 46087
rect 18230 46084 18236 46096
rect 17819 46056 18236 46084
rect 17819 46053 17831 46056
rect 17773 46047 17831 46053
rect 8389 46019 8447 46025
rect 8389 45985 8401 46019
rect 8435 46016 8447 46019
rect 10594 46016 10600 46028
rect 8435 45988 10600 46016
rect 8435 45985 8447 45988
rect 8389 45979 8447 45985
rect 10594 45976 10600 45988
rect 10652 45976 10658 46028
rect 10689 46019 10747 46025
rect 10689 45985 10701 46019
rect 10735 46016 10747 46019
rect 10778 46016 10784 46028
rect 10735 45988 10784 46016
rect 10735 45985 10747 45988
rect 10689 45979 10747 45985
rect 10778 45976 10784 45988
rect 10836 45976 10842 46028
rect 13906 45976 13912 46028
rect 13964 46016 13970 46028
rect 13964 45988 14009 46016
rect 13964 45976 13970 45988
rect 14826 45976 14832 46028
rect 14884 46016 14890 46028
rect 16117 46019 16175 46025
rect 16117 46016 16129 46019
rect 14884 45988 16129 46016
rect 14884 45976 14890 45988
rect 16117 45985 16129 45988
rect 16163 45985 16175 46019
rect 16117 45979 16175 45985
rect 16393 46019 16451 46025
rect 16393 45985 16405 46019
rect 16439 46016 16451 46019
rect 16666 46016 16672 46028
rect 16439 45988 16672 46016
rect 16439 45985 16451 45988
rect 16393 45979 16451 45985
rect 16666 45976 16672 45988
rect 16724 45976 16730 46028
rect 382 45908 388 45960
rect 440 45948 446 45960
rect 2682 45948 2688 45960
rect 440 45920 2688 45948
rect 440 45908 446 45920
rect 2682 45908 2688 45920
rect 2740 45908 2746 45960
rect 4798 45908 4804 45960
rect 4856 45948 4862 45960
rect 4893 45951 4951 45957
rect 4893 45948 4905 45951
rect 4856 45920 4905 45948
rect 4856 45908 4862 45920
rect 4893 45917 4905 45920
rect 4939 45917 4951 45951
rect 4893 45911 4951 45917
rect 5169 45951 5227 45957
rect 5169 45917 5181 45951
rect 5215 45948 5227 45951
rect 5350 45948 5356 45960
rect 5215 45920 5356 45948
rect 5215 45917 5227 45920
rect 5169 45911 5227 45917
rect 5350 45908 5356 45920
rect 5408 45908 5414 45960
rect 10962 45948 10968 45960
rect 10923 45920 10968 45948
rect 10962 45908 10968 45920
rect 11020 45908 11026 45960
rect 15470 45880 15476 45892
rect 13648 45852 15476 45880
rect 13648 45824 13676 45852
rect 15470 45840 15476 45852
rect 15528 45840 15534 45892
rect 8478 45812 8484 45824
rect 8439 45784 8484 45812
rect 8478 45772 8484 45784
rect 8536 45772 8542 45824
rect 13630 45812 13636 45824
rect 13591 45784 13636 45812
rect 13630 45772 13636 45784
rect 13688 45772 13694 45824
rect 14090 45812 14096 45824
rect 14051 45784 14096 45812
rect 14090 45772 14096 45784
rect 14148 45772 14154 45824
rect 15930 45772 15936 45824
rect 15988 45812 15994 45824
rect 17788 45812 17816 46047
rect 18230 46044 18236 46056
rect 18288 46044 18294 46096
rect 15988 45784 17816 45812
rect 15988 45772 15994 45784
rect 1104 45722 24840 45744
rect 1104 45670 4947 45722
rect 4999 45670 5011 45722
rect 5063 45670 5075 45722
rect 5127 45670 5139 45722
rect 5191 45670 12878 45722
rect 12930 45670 12942 45722
rect 12994 45670 13006 45722
rect 13058 45670 13070 45722
rect 13122 45670 20808 45722
rect 20860 45670 20872 45722
rect 20924 45670 20936 45722
rect 20988 45670 21000 45722
rect 21052 45670 24840 45722
rect 1104 45648 24840 45670
rect 5350 45568 5356 45620
rect 5408 45608 5414 45620
rect 5445 45611 5503 45617
rect 5445 45608 5457 45611
rect 5408 45580 5457 45608
rect 5408 45568 5414 45580
rect 5445 45577 5457 45580
rect 5491 45577 5503 45611
rect 8754 45608 8760 45620
rect 8715 45580 8760 45608
rect 5445 45571 5503 45577
rect 8754 45568 8760 45580
rect 8812 45568 8818 45620
rect 13814 45608 13820 45620
rect 13775 45580 13820 45608
rect 13814 45568 13820 45580
rect 13872 45568 13878 45620
rect 16114 45568 16120 45620
rect 16172 45608 16178 45620
rect 16301 45611 16359 45617
rect 16301 45608 16313 45611
rect 16172 45580 16313 45608
rect 16172 45568 16178 45580
rect 16301 45577 16313 45580
rect 16347 45577 16359 45611
rect 16301 45571 16359 45577
rect 11238 45540 11244 45552
rect 11199 45512 11244 45540
rect 11238 45500 11244 45512
rect 11296 45500 11302 45552
rect 9861 45475 9919 45481
rect 9861 45441 9873 45475
rect 9907 45472 9919 45475
rect 10778 45472 10784 45484
rect 9907 45444 10784 45472
rect 9907 45441 9919 45444
rect 9861 45435 9919 45441
rect 10778 45432 10784 45444
rect 10836 45472 10842 45484
rect 12437 45475 12495 45481
rect 12437 45472 12449 45475
rect 10836 45444 12449 45472
rect 10836 45432 10842 45444
rect 12437 45441 12449 45444
rect 12483 45472 12495 45475
rect 13354 45472 13360 45484
rect 12483 45444 13360 45472
rect 12483 45441 12495 45444
rect 12437 45435 12495 45441
rect 13354 45432 13360 45444
rect 13412 45432 13418 45484
rect 15654 45432 15660 45484
rect 15712 45472 15718 45484
rect 18509 45475 18567 45481
rect 18509 45472 18521 45475
rect 15712 45444 18521 45472
rect 15712 45432 15718 45444
rect 18509 45441 18521 45444
rect 18555 45441 18567 45475
rect 18509 45435 18567 45441
rect 4706 45364 4712 45416
rect 4764 45404 4770 45416
rect 4985 45407 5043 45413
rect 4985 45404 4997 45407
rect 4764 45376 4997 45404
rect 4764 45364 4770 45376
rect 4985 45373 4997 45376
rect 5031 45373 5043 45407
rect 5258 45404 5264 45416
rect 5219 45376 5264 45404
rect 4985 45367 5043 45373
rect 5258 45364 5264 45376
rect 5316 45364 5322 45416
rect 5442 45364 5448 45416
rect 5500 45404 5506 45416
rect 6825 45407 6883 45413
rect 6825 45404 6837 45407
rect 5500 45376 6837 45404
rect 5500 45364 5506 45376
rect 6825 45373 6837 45376
rect 6871 45373 6883 45407
rect 6825 45367 6883 45373
rect 7009 45407 7067 45413
rect 7009 45373 7021 45407
rect 7055 45404 7067 45407
rect 7466 45404 7472 45416
rect 7055 45376 7472 45404
rect 7055 45373 7067 45376
rect 7009 45367 7067 45373
rect 7466 45364 7472 45376
rect 7524 45364 7530 45416
rect 7742 45364 7748 45416
rect 7800 45404 7806 45416
rect 8297 45407 8355 45413
rect 8297 45404 8309 45407
rect 7800 45376 8309 45404
rect 7800 45364 7806 45376
rect 8297 45373 8309 45376
rect 8343 45373 8355 45407
rect 8478 45404 8484 45416
rect 8439 45376 8484 45404
rect 8297 45367 8355 45373
rect 8478 45364 8484 45376
rect 8536 45364 8542 45416
rect 8573 45407 8631 45413
rect 8573 45373 8585 45407
rect 8619 45373 8631 45407
rect 10134 45404 10140 45416
rect 10095 45376 10140 45404
rect 8573 45367 8631 45373
rect 5169 45339 5227 45345
rect 5169 45305 5181 45339
rect 5215 45336 5227 45339
rect 5626 45336 5632 45348
rect 5215 45308 5632 45336
rect 5215 45305 5227 45308
rect 5169 45299 5227 45305
rect 5626 45296 5632 45308
rect 5684 45296 5690 45348
rect 8386 45296 8392 45348
rect 8444 45336 8450 45348
rect 8588 45336 8616 45367
rect 10134 45364 10140 45376
rect 10192 45364 10198 45416
rect 12526 45364 12532 45416
rect 12584 45404 12590 45416
rect 12713 45407 12771 45413
rect 12713 45404 12725 45407
rect 12584 45376 12725 45404
rect 12584 45364 12590 45376
rect 12713 45373 12725 45376
rect 12759 45373 12771 45407
rect 12713 45367 12771 45373
rect 14826 45364 14832 45416
rect 14884 45404 14890 45416
rect 14921 45407 14979 45413
rect 14921 45404 14933 45407
rect 14884 45376 14933 45404
rect 14884 45364 14890 45376
rect 14921 45373 14933 45376
rect 14967 45373 14979 45407
rect 15194 45404 15200 45416
rect 15155 45376 15200 45404
rect 14921 45367 14979 45373
rect 15194 45364 15200 45376
rect 15252 45364 15258 45416
rect 18138 45364 18144 45416
rect 18196 45404 18202 45416
rect 18233 45407 18291 45413
rect 18233 45404 18245 45407
rect 18196 45376 18245 45404
rect 18196 45364 18202 45376
rect 18233 45373 18245 45376
rect 18279 45404 18291 45407
rect 18322 45404 18328 45416
rect 18279 45376 18328 45404
rect 18279 45373 18291 45376
rect 18233 45367 18291 45373
rect 18322 45364 18328 45376
rect 18380 45364 18386 45416
rect 18046 45336 18052 45348
rect 8444 45308 8616 45336
rect 18007 45308 18052 45336
rect 8444 45296 8450 45308
rect 18046 45296 18052 45308
rect 18104 45296 18110 45348
rect 4798 45228 4804 45280
rect 4856 45268 4862 45280
rect 7101 45271 7159 45277
rect 7101 45268 7113 45271
rect 4856 45240 7113 45268
rect 4856 45228 4862 45240
rect 7101 45237 7113 45240
rect 7147 45237 7159 45271
rect 7101 45231 7159 45237
rect 1104 45178 24840 45200
rect 1104 45126 8912 45178
rect 8964 45126 8976 45178
rect 9028 45126 9040 45178
rect 9092 45126 9104 45178
rect 9156 45126 16843 45178
rect 16895 45126 16907 45178
rect 16959 45126 16971 45178
rect 17023 45126 17035 45178
rect 17087 45126 24840 45178
rect 1104 45104 24840 45126
rect 7466 45024 7472 45076
rect 7524 45064 7530 45076
rect 7561 45067 7619 45073
rect 7561 45064 7573 45067
rect 7524 45036 7573 45064
rect 7524 45024 7530 45036
rect 7561 45033 7573 45036
rect 7607 45033 7619 45067
rect 12434 45064 12440 45076
rect 7561 45027 7619 45033
rect 11440 45036 12440 45064
rect 4798 44996 4804 45008
rect 4759 44968 4804 44996
rect 4798 44956 4804 44968
rect 4856 44956 4862 45008
rect 9861 44999 9919 45005
rect 9861 44965 9873 44999
rect 9907 44996 9919 44999
rect 10042 44996 10048 45008
rect 9907 44968 10048 44996
rect 9907 44965 9919 44968
rect 9861 44959 9919 44965
rect 10042 44956 10048 44968
rect 10100 44956 10106 45008
rect 11440 45005 11468 45036
rect 12434 45024 12440 45036
rect 12492 45024 12498 45076
rect 11425 44999 11483 45005
rect 11425 44965 11437 44999
rect 11471 44965 11483 44999
rect 11425 44959 11483 44965
rect 11977 44999 12035 45005
rect 11977 44965 11989 44999
rect 12023 44996 12035 44999
rect 12526 44996 12532 45008
rect 12023 44968 12532 44996
rect 12023 44965 12035 44968
rect 11977 44959 12035 44965
rect 12526 44956 12532 44968
rect 12584 44956 12590 45008
rect 12710 44956 12716 45008
rect 12768 44996 12774 45008
rect 12989 44999 13047 45005
rect 12989 44996 13001 44999
rect 12768 44968 13001 44996
rect 12768 44956 12774 44968
rect 12989 44965 13001 44968
rect 13035 44965 13047 44999
rect 12989 44959 13047 44965
rect 13541 44999 13599 45005
rect 13541 44965 13553 44999
rect 13587 44996 13599 44999
rect 15194 44996 15200 45008
rect 13587 44968 15200 44996
rect 13587 44965 13599 44968
rect 13541 44959 13599 44965
rect 15194 44956 15200 44968
rect 15252 44956 15258 45008
rect 17773 44999 17831 45005
rect 17773 44965 17785 44999
rect 17819 44996 17831 44999
rect 18138 44996 18144 45008
rect 17819 44968 18144 44996
rect 17819 44965 17831 44968
rect 17773 44959 17831 44965
rect 18138 44956 18144 44968
rect 18196 44956 18202 45008
rect 4706 44928 4712 44940
rect 4667 44900 4712 44928
rect 4706 44888 4712 44900
rect 4764 44888 4770 44940
rect 4893 44931 4951 44937
rect 4893 44897 4905 44931
rect 4939 44897 4951 44931
rect 4893 44891 4951 44897
rect 5353 44931 5411 44937
rect 5353 44897 5365 44931
rect 5399 44928 5411 44931
rect 6457 44931 6515 44937
rect 6457 44928 6469 44931
rect 5399 44900 6469 44928
rect 5399 44897 5411 44900
rect 5353 44891 5411 44897
rect 6457 44897 6469 44900
rect 6503 44897 6515 44931
rect 6457 44891 6515 44897
rect 4908 44860 4936 44891
rect 9214 44888 9220 44940
rect 9272 44928 9278 44940
rect 9953 44931 10011 44937
rect 9953 44928 9965 44931
rect 9272 44900 9965 44928
rect 9272 44888 9278 44900
rect 9953 44897 9965 44900
rect 9999 44897 10011 44931
rect 11330 44928 11336 44940
rect 11291 44900 11336 44928
rect 9953 44891 10011 44897
rect 11330 44888 11336 44900
rect 11388 44888 11394 44940
rect 11514 44928 11520 44940
rect 11475 44900 11520 44928
rect 11514 44888 11520 44900
rect 11572 44888 11578 44940
rect 12618 44888 12624 44940
rect 12676 44928 12682 44940
rect 13081 44931 13139 44937
rect 13081 44928 13093 44931
rect 12676 44900 13093 44928
rect 12676 44888 12682 44900
rect 13081 44897 13093 44900
rect 13127 44897 13139 44931
rect 13081 44891 13139 44897
rect 16206 44888 16212 44940
rect 16264 44928 16270 44940
rect 16393 44931 16451 44937
rect 16393 44928 16405 44931
rect 16264 44900 16405 44928
rect 16264 44888 16270 44900
rect 16393 44897 16405 44900
rect 16439 44897 16451 44931
rect 16393 44891 16451 44897
rect 5442 44860 5448 44872
rect 4908 44832 5448 44860
rect 5442 44820 5448 44832
rect 5500 44820 5506 44872
rect 6181 44863 6239 44869
rect 6181 44829 6193 44863
rect 6227 44829 6239 44863
rect 6181 44823 6239 44829
rect 9677 44863 9735 44869
rect 9677 44829 9689 44863
rect 9723 44860 9735 44863
rect 11348 44860 11376 44888
rect 9723 44832 11376 44860
rect 9723 44829 9735 44832
rect 9677 44823 9735 44829
rect 4154 44752 4160 44804
rect 4212 44792 4218 44804
rect 4890 44792 4896 44804
rect 4212 44764 4896 44792
rect 4212 44752 4218 44764
rect 4890 44752 4896 44764
rect 4948 44792 4954 44804
rect 6196 44792 6224 44823
rect 14826 44820 14832 44872
rect 14884 44860 14890 44872
rect 16117 44863 16175 44869
rect 16117 44860 16129 44863
rect 14884 44832 16129 44860
rect 14884 44820 14890 44832
rect 16117 44829 16129 44832
rect 16163 44829 16175 44863
rect 16117 44823 16175 44829
rect 4948 44764 6224 44792
rect 4948 44752 4954 44764
rect 10134 44724 10140 44736
rect 10095 44696 10140 44724
rect 10134 44684 10140 44696
rect 10192 44684 10198 44736
rect 12710 44684 12716 44736
rect 12768 44724 12774 44736
rect 12805 44727 12863 44733
rect 12805 44724 12817 44727
rect 12768 44696 12817 44724
rect 12768 44684 12774 44696
rect 12805 44693 12817 44696
rect 12851 44724 12863 44727
rect 13630 44724 13636 44736
rect 12851 44696 13636 44724
rect 12851 44693 12863 44696
rect 12805 44687 12863 44693
rect 13630 44684 13636 44696
rect 13688 44684 13694 44736
rect 1104 44634 24840 44656
rect 1104 44582 4947 44634
rect 4999 44582 5011 44634
rect 5063 44582 5075 44634
rect 5127 44582 5139 44634
rect 5191 44582 12878 44634
rect 12930 44582 12942 44634
rect 12994 44582 13006 44634
rect 13058 44582 13070 44634
rect 13122 44582 20808 44634
rect 20860 44582 20872 44634
rect 20924 44582 20936 44634
rect 20988 44582 21000 44634
rect 21052 44582 24840 44634
rect 1104 44560 24840 44582
rect 5350 44480 5356 44532
rect 5408 44520 5414 44532
rect 5629 44523 5687 44529
rect 5629 44520 5641 44523
rect 5408 44492 5641 44520
rect 5408 44480 5414 44492
rect 5629 44489 5641 44492
rect 5675 44489 5687 44523
rect 5629 44483 5687 44489
rect 9217 44523 9275 44529
rect 9217 44489 9229 44523
rect 9263 44520 9275 44523
rect 9766 44520 9772 44532
rect 9263 44492 9772 44520
rect 9263 44489 9275 44492
rect 9217 44483 9275 44489
rect 9766 44480 9772 44492
rect 9824 44480 9830 44532
rect 10781 44523 10839 44529
rect 10781 44489 10793 44523
rect 10827 44520 10839 44523
rect 10962 44520 10968 44532
rect 10827 44492 10968 44520
rect 10827 44489 10839 44492
rect 10781 44483 10839 44489
rect 10962 44480 10968 44492
rect 11020 44480 11026 44532
rect 15194 44520 15200 44532
rect 12728 44492 15200 44520
rect 5368 44384 5396 44480
rect 10321 44455 10379 44461
rect 10321 44421 10333 44455
rect 10367 44452 10379 44455
rect 11330 44452 11336 44464
rect 10367 44424 11336 44452
rect 10367 44421 10379 44424
rect 10321 44415 10379 44421
rect 11330 44412 11336 44424
rect 11388 44412 11394 44464
rect 7650 44384 7656 44396
rect 3068 44356 5396 44384
rect 7611 44356 7656 44384
rect 3068 44325 3096 44356
rect 7650 44344 7656 44356
rect 7708 44344 7714 44396
rect 3053 44319 3111 44325
rect 3053 44285 3065 44319
rect 3099 44285 3111 44319
rect 3053 44279 3111 44285
rect 4154 44276 4160 44328
rect 4212 44316 4218 44328
rect 4249 44319 4307 44325
rect 4249 44316 4261 44319
rect 4212 44288 4261 44316
rect 4212 44276 4218 44288
rect 4249 44285 4261 44288
rect 4295 44285 4307 44319
rect 4249 44279 4307 44285
rect 4525 44319 4583 44325
rect 4525 44285 4537 44319
rect 4571 44316 4583 44319
rect 4798 44316 4804 44328
rect 4571 44288 4804 44316
rect 4571 44285 4583 44288
rect 4525 44279 4583 44285
rect 4798 44276 4804 44288
rect 4856 44276 4862 44328
rect 5350 44276 5356 44328
rect 5408 44316 5414 44328
rect 5534 44316 5540 44328
rect 5408 44288 5540 44316
rect 5408 44276 5414 44288
rect 5534 44276 5540 44288
rect 5592 44276 5598 44328
rect 7926 44316 7932 44328
rect 7887 44288 7932 44316
rect 7926 44276 7932 44288
rect 7984 44276 7990 44328
rect 10410 44276 10416 44328
rect 10468 44316 10474 44328
rect 12728 44325 12756 44492
rect 15194 44480 15200 44492
rect 15252 44480 15258 44532
rect 15289 44523 15347 44529
rect 15289 44489 15301 44523
rect 15335 44520 15347 44523
rect 15470 44520 15476 44532
rect 15335 44492 15476 44520
rect 15335 44489 15347 44492
rect 15289 44483 15347 44489
rect 15470 44480 15476 44492
rect 15528 44480 15534 44532
rect 15930 44452 15936 44464
rect 14384 44424 15936 44452
rect 10597 44319 10655 44325
rect 10597 44316 10609 44319
rect 10468 44288 10609 44316
rect 10468 44276 10474 44288
rect 10597 44285 10609 44288
rect 10643 44285 10655 44319
rect 10597 44279 10655 44285
rect 12713 44319 12771 44325
rect 12713 44285 12725 44319
rect 12759 44285 12771 44319
rect 12713 44279 12771 44285
rect 13906 44276 13912 44328
rect 13964 44316 13970 44328
rect 14093 44319 14151 44325
rect 13964 44288 14009 44316
rect 13964 44276 13970 44288
rect 14093 44285 14105 44319
rect 14139 44316 14151 44319
rect 14384 44316 14412 44424
rect 15930 44412 15936 44424
rect 15988 44412 15994 44464
rect 14461 44387 14519 44393
rect 14461 44353 14473 44387
rect 14507 44384 14519 44387
rect 15378 44384 15384 44396
rect 14507 44356 15384 44384
rect 14507 44353 14519 44356
rect 14461 44347 14519 44353
rect 15378 44344 15384 44356
rect 15436 44344 15442 44396
rect 18322 44384 18328 44396
rect 15488 44356 18328 44384
rect 15488 44325 15516 44356
rect 18322 44344 18328 44356
rect 18380 44344 18386 44396
rect 14139 44288 14412 44316
rect 15473 44319 15531 44325
rect 14139 44285 14151 44288
rect 14093 44279 14151 44285
rect 15473 44285 15485 44319
rect 15519 44285 15531 44319
rect 15473 44279 15531 44285
rect 15565 44319 15623 44325
rect 15565 44285 15577 44319
rect 15611 44316 15623 44319
rect 15654 44316 15660 44328
rect 15611 44288 15660 44316
rect 15611 44285 15623 44288
rect 15565 44279 15623 44285
rect 15654 44276 15660 44288
rect 15712 44276 15718 44328
rect 16853 44319 16911 44325
rect 16853 44285 16865 44319
rect 16899 44316 16911 44319
rect 17862 44316 17868 44328
rect 16899 44288 17868 44316
rect 16899 44285 16911 44288
rect 16853 44279 16911 44285
rect 17862 44276 17868 44288
rect 17920 44276 17926 44328
rect 2869 44251 2927 44257
rect 2869 44217 2881 44251
rect 2915 44217 2927 44251
rect 3418 44248 3424 44260
rect 3379 44220 3424 44248
rect 2869 44211 2927 44217
rect 2884 44180 2912 44211
rect 3418 44208 3424 44220
rect 3476 44208 3482 44260
rect 10505 44251 10563 44257
rect 10505 44217 10517 44251
rect 10551 44248 10563 44251
rect 11422 44248 11428 44260
rect 10551 44220 11428 44248
rect 10551 44217 10563 44220
rect 10505 44211 10563 44217
rect 11422 44208 11428 44220
rect 11480 44208 11486 44260
rect 12434 44208 12440 44260
rect 12492 44248 12498 44260
rect 12529 44251 12587 44257
rect 12529 44248 12541 44251
rect 12492 44220 12541 44248
rect 12492 44208 12498 44220
rect 12529 44217 12541 44220
rect 12575 44248 12587 44251
rect 13170 44248 13176 44260
rect 12575 44220 13176 44248
rect 12575 44217 12587 44220
rect 12529 44211 12587 44217
rect 13170 44208 13176 44220
rect 13228 44248 13234 44260
rect 16025 44251 16083 44257
rect 13228 44220 15424 44248
rect 13228 44208 13234 44220
rect 5350 44180 5356 44192
rect 2884 44152 5356 44180
rect 5350 44140 5356 44152
rect 5408 44140 5414 44192
rect 12802 44180 12808 44192
rect 12763 44152 12808 44180
rect 12802 44140 12808 44152
rect 12860 44140 12866 44192
rect 15396 44180 15424 44220
rect 16025 44217 16037 44251
rect 16071 44248 16083 44251
rect 16298 44248 16304 44260
rect 16071 44220 16304 44248
rect 16071 44217 16083 44220
rect 16025 44211 16083 44217
rect 16298 44208 16304 44220
rect 16356 44208 16362 44260
rect 17037 44183 17095 44189
rect 17037 44180 17049 44183
rect 15396 44152 17049 44180
rect 17037 44149 17049 44152
rect 17083 44149 17095 44183
rect 17037 44143 17095 44149
rect 1104 44090 24840 44112
rect 1104 44038 8912 44090
rect 8964 44038 8976 44090
rect 9028 44038 9040 44090
rect 9092 44038 9104 44090
rect 9156 44038 16843 44090
rect 16895 44038 16907 44090
rect 16959 44038 16971 44090
rect 17023 44038 17035 44090
rect 17087 44038 24840 44090
rect 1104 44016 24840 44038
rect 6549 43979 6607 43985
rect 6549 43945 6561 43979
rect 6595 43976 6607 43979
rect 8202 43976 8208 43988
rect 6595 43948 8208 43976
rect 6595 43945 6607 43948
rect 6549 43939 6607 43945
rect 8202 43936 8208 43948
rect 8260 43936 8266 43988
rect 13538 43976 13544 43988
rect 10336 43948 13544 43976
rect 3418 43868 3424 43920
rect 3476 43908 3482 43920
rect 4893 43911 4951 43917
rect 4893 43908 4905 43911
rect 3476 43880 4905 43908
rect 3476 43868 3482 43880
rect 4893 43877 4905 43880
rect 4939 43877 4951 43911
rect 4893 43871 4951 43877
rect 7374 43868 7380 43920
rect 7432 43908 7438 43920
rect 8110 43908 8116 43920
rect 7432 43880 8116 43908
rect 7432 43868 7438 43880
rect 8110 43868 8116 43880
rect 8168 43868 8174 43920
rect 4706 43800 4712 43852
rect 4764 43840 4770 43852
rect 4985 43843 5043 43849
rect 4985 43840 4997 43843
rect 4764 43812 4997 43840
rect 4764 43800 4770 43812
rect 4985 43809 4997 43812
rect 5031 43809 5043 43843
rect 6362 43840 6368 43852
rect 6323 43812 6368 43840
rect 4985 43803 5043 43809
rect 6362 43800 6368 43812
rect 6420 43800 6426 43852
rect 7650 43840 7656 43852
rect 7611 43812 7656 43840
rect 7650 43800 7656 43812
rect 7708 43800 7714 43852
rect 10336 43849 10364 43948
rect 13538 43936 13544 43948
rect 13596 43936 13602 43988
rect 11701 43911 11759 43917
rect 11701 43877 11713 43911
rect 11747 43908 11759 43911
rect 12802 43908 12808 43920
rect 11747 43880 12808 43908
rect 11747 43877 11759 43880
rect 11701 43871 11759 43877
rect 12802 43868 12808 43880
rect 12860 43868 12866 43920
rect 17681 43911 17739 43917
rect 17681 43877 17693 43911
rect 17727 43908 17739 43911
rect 17954 43908 17960 43920
rect 17727 43880 17960 43908
rect 17727 43877 17739 43880
rect 17681 43871 17739 43877
rect 17954 43868 17960 43880
rect 18012 43868 18018 43920
rect 7745 43843 7803 43849
rect 7745 43809 7757 43843
rect 7791 43809 7803 43843
rect 7745 43803 7803 43809
rect 10137 43843 10195 43849
rect 10137 43809 10149 43843
rect 10183 43809 10195 43843
rect 10137 43803 10195 43809
rect 10321 43843 10379 43849
rect 10321 43809 10333 43843
rect 10367 43809 10379 43843
rect 10321 43803 10379 43809
rect 7558 43732 7564 43784
rect 7616 43772 7622 43784
rect 7760 43772 7788 43803
rect 7616 43744 7788 43772
rect 7616 43732 7622 43744
rect 4614 43664 4620 43716
rect 4672 43704 4678 43716
rect 4709 43707 4767 43713
rect 4709 43704 4721 43707
rect 4672 43676 4721 43704
rect 4672 43664 4678 43676
rect 4709 43673 4721 43676
rect 4755 43673 4767 43707
rect 10152 43704 10180 43803
rect 11422 43800 11428 43852
rect 11480 43840 11486 43852
rect 11793 43843 11851 43849
rect 11793 43840 11805 43843
rect 11480 43812 11805 43840
rect 11480 43800 11486 43812
rect 11793 43809 11805 43812
rect 11839 43809 11851 43843
rect 13538 43840 13544 43852
rect 13499 43812 13544 43840
rect 11793 43803 11851 43809
rect 13538 43800 13544 43812
rect 13596 43800 13602 43852
rect 13633 43843 13691 43849
rect 13633 43809 13645 43843
rect 13679 43809 13691 43843
rect 16298 43840 16304 43852
rect 16259 43812 16304 43840
rect 13633 43803 13691 43809
rect 11330 43732 11336 43784
rect 11388 43772 11394 43784
rect 11517 43775 11575 43781
rect 11517 43772 11529 43775
rect 11388 43744 11529 43772
rect 11388 43732 11394 43744
rect 11517 43741 11529 43744
rect 11563 43741 11575 43775
rect 12250 43772 12256 43784
rect 12211 43744 12256 43772
rect 11517 43735 11575 43741
rect 12250 43732 12256 43744
rect 12308 43732 12314 43784
rect 12526 43732 12532 43784
rect 12584 43772 12590 43784
rect 13648 43772 13676 43803
rect 16298 43800 16304 43812
rect 16356 43800 16362 43852
rect 14090 43772 14096 43784
rect 12584 43744 13676 43772
rect 14051 43744 14096 43772
rect 12584 43732 12590 43744
rect 14090 43732 14096 43744
rect 14148 43732 14154 43784
rect 14826 43732 14832 43784
rect 14884 43772 14890 43784
rect 16025 43775 16083 43781
rect 16025 43772 16037 43775
rect 14884 43744 16037 43772
rect 14884 43732 14890 43744
rect 16025 43741 16037 43744
rect 16071 43741 16083 43775
rect 16025 43735 16083 43741
rect 12434 43704 12440 43716
rect 10152 43676 12440 43704
rect 4709 43667 4767 43673
rect 12434 43664 12440 43676
rect 12492 43664 12498 43716
rect 4798 43596 4804 43648
rect 4856 43636 4862 43648
rect 5169 43639 5227 43645
rect 5169 43636 5181 43639
rect 4856 43608 5181 43636
rect 4856 43596 4862 43608
rect 5169 43605 5181 43608
rect 5215 43605 5227 43639
rect 5169 43599 5227 43605
rect 6914 43596 6920 43648
rect 6972 43636 6978 43648
rect 7469 43639 7527 43645
rect 7469 43636 7481 43639
rect 6972 43608 7481 43636
rect 6972 43596 6978 43608
rect 7469 43605 7481 43608
rect 7515 43636 7527 43639
rect 7742 43636 7748 43648
rect 7515 43608 7748 43636
rect 7515 43605 7527 43608
rect 7469 43599 7527 43605
rect 7742 43596 7748 43608
rect 7800 43596 7806 43648
rect 7926 43636 7932 43648
rect 7887 43608 7932 43636
rect 7926 43596 7932 43608
rect 7984 43596 7990 43648
rect 10413 43639 10471 43645
rect 10413 43605 10425 43639
rect 10459 43636 10471 43639
rect 10502 43636 10508 43648
rect 10459 43608 10508 43636
rect 10459 43605 10471 43608
rect 10413 43599 10471 43605
rect 10502 43596 10508 43608
rect 10560 43596 10566 43648
rect 12710 43596 12716 43648
rect 12768 43636 12774 43648
rect 13357 43639 13415 43645
rect 13357 43636 13369 43639
rect 12768 43608 13369 43636
rect 12768 43596 12774 43608
rect 13357 43605 13369 43608
rect 13403 43605 13415 43639
rect 13357 43599 13415 43605
rect 1104 43546 24840 43568
rect 1104 43494 4947 43546
rect 4999 43494 5011 43546
rect 5063 43494 5075 43546
rect 5127 43494 5139 43546
rect 5191 43494 12878 43546
rect 12930 43494 12942 43546
rect 12994 43494 13006 43546
rect 13058 43494 13070 43546
rect 13122 43494 20808 43546
rect 20860 43494 20872 43546
rect 20924 43494 20936 43546
rect 20988 43494 21000 43546
rect 21052 43494 24840 43546
rect 1104 43472 24840 43494
rect 10321 43435 10379 43441
rect 10321 43401 10333 43435
rect 10367 43432 10379 43435
rect 11330 43432 11336 43444
rect 10367 43404 11336 43432
rect 10367 43401 10379 43404
rect 10321 43395 10379 43401
rect 11330 43392 11336 43404
rect 11388 43392 11394 43444
rect 14001 43435 14059 43441
rect 14001 43401 14013 43435
rect 14047 43432 14059 43435
rect 15286 43432 15292 43444
rect 14047 43404 15292 43432
rect 14047 43401 14059 43404
rect 14001 43395 14059 43401
rect 15286 43392 15292 43404
rect 15344 43392 15350 43444
rect 18322 43432 18328 43444
rect 18283 43404 18328 43432
rect 18322 43392 18328 43404
rect 18380 43392 18386 43444
rect 3510 43256 3516 43308
rect 3568 43296 3574 43308
rect 9306 43296 9312 43308
rect 3568 43268 3740 43296
rect 3568 43256 3574 43268
rect 3712 43240 3740 43268
rect 7760 43268 9312 43296
rect 3694 43228 3700 43240
rect 3607 43200 3700 43228
rect 3694 43188 3700 43200
rect 3752 43188 3758 43240
rect 5350 43228 5356 43240
rect 5311 43200 5356 43228
rect 5350 43188 5356 43200
rect 5408 43188 5414 43240
rect 5537 43231 5595 43237
rect 5537 43197 5549 43231
rect 5583 43228 5595 43231
rect 7374 43228 7380 43240
rect 5583 43200 7380 43228
rect 5583 43197 5595 43200
rect 5537 43191 5595 43197
rect 7374 43188 7380 43200
rect 7432 43188 7438 43240
rect 7760 43237 7788 43268
rect 9306 43256 9312 43268
rect 9364 43256 9370 43308
rect 11606 43296 11612 43308
rect 10428 43268 11612 43296
rect 7745 43231 7803 43237
rect 7745 43197 7757 43231
rect 7791 43197 7803 43231
rect 7745 43191 7803 43197
rect 8202 43188 8208 43240
rect 8260 43228 8266 43240
rect 8941 43231 8999 43237
rect 8941 43228 8953 43231
rect 8260 43200 8953 43228
rect 8260 43188 8266 43200
rect 8941 43197 8953 43200
rect 8987 43197 8999 43231
rect 8941 43191 8999 43197
rect 9125 43231 9183 43237
rect 9125 43197 9137 43231
rect 9171 43228 9183 43231
rect 10428 43228 10456 43268
rect 11606 43256 11612 43268
rect 11664 43256 11670 43308
rect 12250 43256 12256 43308
rect 12308 43296 12314 43308
rect 12713 43299 12771 43305
rect 12713 43296 12725 43299
rect 12308 43268 12725 43296
rect 12308 43256 12314 43268
rect 12713 43265 12725 43268
rect 12759 43265 12771 43299
rect 12713 43259 12771 43265
rect 14090 43256 14096 43308
rect 14148 43296 14154 43308
rect 15197 43299 15255 43305
rect 15197 43296 15209 43299
rect 14148 43268 15209 43296
rect 14148 43256 14154 43268
rect 15197 43265 15209 43268
rect 15243 43265 15255 43299
rect 15197 43259 15255 43265
rect 10594 43228 10600 43240
rect 9171 43200 10456 43228
rect 10555 43200 10600 43228
rect 9171 43197 9183 43200
rect 9125 43191 9183 43197
rect 10594 43188 10600 43200
rect 10652 43188 10658 43240
rect 12437 43231 12495 43237
rect 12437 43197 12449 43231
rect 12483 43228 12495 43231
rect 12802 43228 12808 43240
rect 12483 43200 12808 43228
rect 12483 43197 12495 43200
rect 12437 43191 12495 43197
rect 12802 43188 12808 43200
rect 12860 43228 12866 43240
rect 13354 43228 13360 43240
rect 12860 43200 13360 43228
rect 12860 43188 12866 43200
rect 13354 43188 13360 43200
rect 13412 43188 13418 43240
rect 14826 43188 14832 43240
rect 14884 43228 14890 43240
rect 14921 43231 14979 43237
rect 14921 43228 14933 43231
rect 14884 43200 14933 43228
rect 14884 43188 14890 43200
rect 14921 43197 14933 43200
rect 14967 43197 14979 43231
rect 14921 43191 14979 43197
rect 17954 43188 17960 43240
rect 18012 43228 18018 43240
rect 18233 43231 18291 43237
rect 18233 43228 18245 43231
rect 18012 43200 18245 43228
rect 18012 43188 18018 43200
rect 18233 43197 18245 43200
rect 18279 43197 18291 43231
rect 18233 43191 18291 43197
rect 2590 43120 2596 43172
rect 2648 43160 2654 43172
rect 3513 43163 3571 43169
rect 3513 43160 3525 43163
rect 2648 43132 3525 43160
rect 2648 43120 2654 43132
rect 3513 43129 3525 43132
rect 3559 43129 3571 43163
rect 5902 43160 5908 43172
rect 5863 43132 5908 43160
rect 3513 43123 3571 43129
rect 5902 43120 5908 43132
rect 5960 43120 5966 43172
rect 7561 43163 7619 43169
rect 7561 43129 7573 43163
rect 7607 43160 7619 43163
rect 8220 43160 8248 43188
rect 9490 43160 9496 43172
rect 7607 43132 8248 43160
rect 9451 43132 9496 43160
rect 7607 43129 7619 43132
rect 7561 43123 7619 43129
rect 9490 43120 9496 43132
rect 9548 43120 9554 43172
rect 10502 43160 10508 43172
rect 10463 43132 10508 43160
rect 10502 43120 10508 43132
rect 10560 43120 10566 43172
rect 11057 43163 11115 43169
rect 11057 43129 11069 43163
rect 11103 43129 11115 43163
rect 18046 43160 18052 43172
rect 18007 43132 18052 43160
rect 11057 43123 11115 43129
rect 3142 43052 3148 43104
rect 3200 43092 3206 43104
rect 3789 43095 3847 43101
rect 3789 43092 3801 43095
rect 3200 43064 3801 43092
rect 3200 43052 3206 43064
rect 3789 43061 3801 43064
rect 3835 43061 3847 43095
rect 3789 43055 3847 43061
rect 7742 43052 7748 43104
rect 7800 43092 7806 43104
rect 7837 43095 7895 43101
rect 7837 43092 7849 43095
rect 7800 43064 7849 43092
rect 7800 43052 7806 43064
rect 7837 43061 7849 43064
rect 7883 43061 7895 43095
rect 11072 43092 11100 43123
rect 18046 43120 18052 43132
rect 18104 43120 18110 43172
rect 12434 43092 12440 43104
rect 11072 43064 12440 43092
rect 7837 43055 7895 43061
rect 12434 43052 12440 43064
rect 12492 43052 12498 43104
rect 14274 43052 14280 43104
rect 14332 43092 14338 43104
rect 16301 43095 16359 43101
rect 16301 43092 16313 43095
rect 14332 43064 16313 43092
rect 14332 43052 14338 43064
rect 16301 43061 16313 43064
rect 16347 43092 16359 43095
rect 16482 43092 16488 43104
rect 16347 43064 16488 43092
rect 16347 43061 16359 43064
rect 16301 43055 16359 43061
rect 16482 43052 16488 43064
rect 16540 43052 16546 43104
rect 1104 43002 24840 43024
rect 1104 42950 8912 43002
rect 8964 42950 8976 43002
rect 9028 42950 9040 43002
rect 9092 42950 9104 43002
rect 9156 42950 16843 43002
rect 16895 42950 16907 43002
rect 16959 42950 16971 43002
rect 17023 42950 17035 43002
rect 17087 42950 24840 43002
rect 1104 42928 24840 42950
rect 13446 42848 13452 42900
rect 13504 42888 13510 42900
rect 13541 42891 13599 42897
rect 13541 42888 13553 42891
rect 13504 42860 13553 42888
rect 13504 42848 13510 42860
rect 13541 42857 13553 42860
rect 13587 42857 13599 42891
rect 13541 42851 13599 42857
rect 4157 42823 4215 42829
rect 4157 42789 4169 42823
rect 4203 42820 4215 42823
rect 4430 42820 4436 42832
rect 4203 42792 4436 42820
rect 4203 42789 4215 42792
rect 4157 42783 4215 42789
rect 4430 42780 4436 42792
rect 4488 42820 4494 42832
rect 5350 42820 5356 42832
rect 4488 42792 5356 42820
rect 4488 42780 4494 42792
rect 5350 42780 5356 42792
rect 5408 42780 5414 42832
rect 8202 42820 8208 42832
rect 8163 42792 8208 42820
rect 8202 42780 8208 42792
rect 8260 42780 8266 42832
rect 1765 42755 1823 42761
rect 1765 42721 1777 42755
rect 1811 42752 1823 42755
rect 2869 42755 2927 42761
rect 2869 42752 2881 42755
rect 1811 42724 2881 42752
rect 1811 42721 1823 42724
rect 1765 42715 1823 42721
rect 2869 42721 2881 42724
rect 2915 42752 2927 42755
rect 4065 42755 4123 42761
rect 4065 42752 4077 42755
rect 2915 42724 4077 42752
rect 2915 42721 2927 42724
rect 2869 42715 2927 42721
rect 4065 42721 4077 42724
rect 4111 42721 4123 42755
rect 4065 42715 4123 42721
rect 4341 42755 4399 42761
rect 4341 42721 4353 42755
rect 4387 42752 4399 42755
rect 8389 42755 8447 42761
rect 4387 42724 6684 42752
rect 4387 42721 4399 42724
rect 4341 42715 4399 42721
rect 6656 42696 6684 42724
rect 8389 42721 8401 42755
rect 8435 42752 8447 42755
rect 9582 42752 9588 42764
rect 8435 42724 9588 42752
rect 8435 42721 8447 42724
rect 8389 42715 8447 42721
rect 9582 42712 9588 42724
rect 9640 42712 9646 42764
rect 9677 42755 9735 42761
rect 9677 42721 9689 42755
rect 9723 42752 9735 42755
rect 12161 42755 12219 42761
rect 12161 42752 12173 42755
rect 9723 42724 12173 42752
rect 9723 42721 9735 42724
rect 9677 42715 9735 42721
rect 12161 42721 12173 42724
rect 12207 42721 12219 42755
rect 12434 42752 12440 42764
rect 12395 42724 12440 42752
rect 12161 42715 12219 42721
rect 4709 42687 4767 42693
rect 4709 42653 4721 42687
rect 4755 42684 4767 42687
rect 5350 42684 5356 42696
rect 4755 42656 5356 42684
rect 4755 42653 4767 42656
rect 4709 42647 4767 42653
rect 5350 42644 5356 42656
rect 5408 42644 5414 42696
rect 5537 42687 5595 42693
rect 5537 42653 5549 42687
rect 5583 42653 5595 42687
rect 5810 42684 5816 42696
rect 5771 42656 5816 42684
rect 5537 42647 5595 42653
rect 1949 42619 2007 42625
rect 1949 42585 1961 42619
rect 1995 42616 2007 42619
rect 4614 42616 4620 42628
rect 1995 42588 4620 42616
rect 1995 42585 2007 42588
rect 1949 42579 2007 42585
rect 4614 42576 4620 42588
rect 4672 42576 4678 42628
rect 4798 42576 4804 42628
rect 4856 42616 4862 42628
rect 5552 42616 5580 42647
rect 5810 42644 5816 42656
rect 5868 42644 5874 42696
rect 6638 42644 6644 42696
rect 6696 42684 6702 42696
rect 6917 42687 6975 42693
rect 6917 42684 6929 42687
rect 6696 42656 6929 42684
rect 6696 42644 6702 42656
rect 6917 42653 6929 42656
rect 6963 42653 6975 42687
rect 9950 42684 9956 42696
rect 9911 42656 9956 42684
rect 6917 42647 6975 42653
rect 9950 42644 9956 42656
rect 10008 42644 10014 42696
rect 11333 42687 11391 42693
rect 11333 42653 11345 42687
rect 11379 42684 11391 42687
rect 11606 42684 11612 42696
rect 11379 42656 11612 42684
rect 11379 42653 11391 42656
rect 11333 42647 11391 42653
rect 11606 42644 11612 42656
rect 11664 42644 11670 42696
rect 12176 42684 12204 42715
rect 12434 42712 12440 42724
rect 12492 42712 12498 42764
rect 15378 42752 15384 42764
rect 15339 42724 15384 42752
rect 15378 42712 15384 42724
rect 15436 42712 15442 42764
rect 15565 42755 15623 42761
rect 15565 42721 15577 42755
rect 15611 42752 15623 42755
rect 18322 42752 18328 42764
rect 15611 42724 18328 42752
rect 15611 42721 15623 42724
rect 15565 42715 15623 42721
rect 18322 42712 18328 42724
rect 18380 42712 18386 42764
rect 18417 42755 18475 42761
rect 18417 42721 18429 42755
rect 18463 42752 18475 42755
rect 21266 42752 21272 42764
rect 18463 42724 21272 42752
rect 18463 42721 18475 42724
rect 18417 42715 18475 42721
rect 12802 42684 12808 42696
rect 12176 42656 12808 42684
rect 4856 42588 5580 42616
rect 4856 42576 4862 42588
rect 3053 42551 3111 42557
rect 3053 42517 3065 42551
rect 3099 42548 3111 42551
rect 3970 42548 3976 42560
rect 3099 42520 3976 42548
rect 3099 42517 3111 42520
rect 3053 42511 3111 42517
rect 3970 42508 3976 42520
rect 4028 42508 4034 42560
rect 4065 42551 4123 42557
rect 4065 42517 4077 42551
rect 4111 42548 4123 42551
rect 6822 42548 6828 42560
rect 4111 42520 6828 42548
rect 4111 42517 4123 42520
rect 4065 42511 4123 42517
rect 6822 42508 6828 42520
rect 6880 42508 6886 42560
rect 7650 42508 7656 42560
rect 7708 42548 7714 42560
rect 8481 42551 8539 42557
rect 8481 42548 8493 42551
rect 7708 42520 8493 42548
rect 7708 42508 7714 42520
rect 8481 42517 8493 42520
rect 8527 42517 8539 42551
rect 12176 42548 12204 42656
rect 12802 42644 12808 42656
rect 12860 42644 12866 42696
rect 15933 42687 15991 42693
rect 15933 42653 15945 42687
rect 15979 42684 15991 42687
rect 16114 42684 16120 42696
rect 15979 42656 16120 42684
rect 15979 42653 15991 42656
rect 15933 42647 15991 42653
rect 16114 42644 16120 42656
rect 16172 42644 16178 42696
rect 16761 42687 16819 42693
rect 16761 42653 16773 42687
rect 16807 42653 16819 42687
rect 17034 42684 17040 42696
rect 16995 42656 17040 42684
rect 16761 42647 16819 42653
rect 14826 42576 14832 42628
rect 14884 42616 14890 42628
rect 16574 42616 16580 42628
rect 14884 42588 16580 42616
rect 14884 42576 14890 42588
rect 16574 42576 16580 42588
rect 16632 42616 16638 42628
rect 16776 42616 16804 42647
rect 17034 42644 17040 42656
rect 17092 42644 17098 42696
rect 16632 42588 16804 42616
rect 16632 42576 16638 42588
rect 12434 42548 12440 42560
rect 12176 42520 12440 42548
rect 8481 42511 8539 42517
rect 12434 42508 12440 42520
rect 12492 42508 12498 42560
rect 15562 42508 15568 42560
rect 15620 42548 15626 42560
rect 18432 42548 18460 42715
rect 21266 42712 21272 42724
rect 21324 42712 21330 42764
rect 15620 42520 18460 42548
rect 15620 42508 15626 42520
rect 1104 42458 24840 42480
rect 1104 42406 4947 42458
rect 4999 42406 5011 42458
rect 5063 42406 5075 42458
rect 5127 42406 5139 42458
rect 5191 42406 12878 42458
rect 12930 42406 12942 42458
rect 12994 42406 13006 42458
rect 13058 42406 13070 42458
rect 13122 42406 20808 42458
rect 20860 42406 20872 42458
rect 20924 42406 20936 42458
rect 20988 42406 21000 42458
rect 21052 42406 24840 42458
rect 1104 42384 24840 42406
rect 3694 42304 3700 42356
rect 3752 42344 3758 42356
rect 4249 42347 4307 42353
rect 4249 42344 4261 42347
rect 3752 42316 4261 42344
rect 3752 42304 3758 42316
rect 4249 42313 4261 42316
rect 4295 42313 4307 42347
rect 4249 42307 4307 42313
rect 4614 42304 4620 42356
rect 4672 42344 4678 42356
rect 5169 42347 5227 42353
rect 5169 42344 5181 42347
rect 4672 42316 5181 42344
rect 4672 42304 4678 42316
rect 5169 42313 5181 42316
rect 5215 42313 5227 42347
rect 5169 42307 5227 42313
rect 5629 42347 5687 42353
rect 5629 42313 5641 42347
rect 5675 42344 5687 42347
rect 5810 42344 5816 42356
rect 5675 42316 5816 42344
rect 5675 42313 5687 42316
rect 5629 42307 5687 42313
rect 5810 42304 5816 42316
rect 5868 42304 5874 42356
rect 9125 42347 9183 42353
rect 9125 42313 9137 42347
rect 9171 42344 9183 42347
rect 9306 42344 9312 42356
rect 9171 42316 9312 42344
rect 9171 42313 9183 42316
rect 9125 42307 9183 42313
rect 9306 42304 9312 42316
rect 9364 42304 9370 42356
rect 13906 42344 13912 42356
rect 13096 42316 13912 42344
rect 4154 42236 4160 42288
rect 4212 42276 4218 42288
rect 4798 42276 4804 42288
rect 4212 42248 4804 42276
rect 4212 42236 4218 42248
rect 4798 42236 4804 42248
rect 4856 42236 4862 42288
rect 2685 42211 2743 42217
rect 2685 42177 2697 42211
rect 2731 42208 2743 42211
rect 4172 42208 4200 42236
rect 6914 42208 6920 42220
rect 2731 42180 4200 42208
rect 5184 42180 6920 42208
rect 2731 42177 2743 42180
rect 2685 42171 2743 42177
rect 2961 42143 3019 42149
rect 2961 42109 2973 42143
rect 3007 42140 3019 42143
rect 3418 42140 3424 42152
rect 3007 42112 3424 42140
rect 3007 42109 3019 42112
rect 2961 42103 3019 42109
rect 3418 42100 3424 42112
rect 3476 42100 3482 42152
rect 3970 42100 3976 42152
rect 4028 42140 4034 42152
rect 5184 42140 5212 42180
rect 6914 42168 6920 42180
rect 6972 42168 6978 42220
rect 7006 42168 7012 42220
rect 7064 42208 7070 42220
rect 7466 42208 7472 42220
rect 7064 42180 7472 42208
rect 7064 42168 7070 42180
rect 7466 42168 7472 42180
rect 7524 42208 7530 42220
rect 7561 42211 7619 42217
rect 7561 42208 7573 42211
rect 7524 42180 7573 42208
rect 7524 42168 7530 42180
rect 7561 42177 7573 42180
rect 7607 42177 7619 42211
rect 7561 42171 7619 42177
rect 11149 42211 11207 42217
rect 11149 42177 11161 42211
rect 11195 42208 11207 42211
rect 11514 42208 11520 42220
rect 11195 42180 11520 42208
rect 11195 42177 11207 42180
rect 11149 42171 11207 42177
rect 11514 42168 11520 42180
rect 11572 42168 11578 42220
rect 5350 42140 5356 42152
rect 4028 42112 5212 42140
rect 5311 42112 5356 42140
rect 4028 42100 4034 42112
rect 5350 42100 5356 42112
rect 5408 42100 5414 42152
rect 5445 42143 5503 42149
rect 5445 42109 5457 42143
rect 5491 42140 5503 42143
rect 5534 42140 5540 42152
rect 5491 42112 5540 42140
rect 5491 42109 5503 42112
rect 5445 42103 5503 42109
rect 5534 42100 5540 42112
rect 5592 42100 5598 42152
rect 7834 42140 7840 42152
rect 7795 42112 7840 42140
rect 7834 42100 7840 42112
rect 7892 42100 7898 42152
rect 10686 42100 10692 42152
rect 10744 42140 10750 42152
rect 10781 42143 10839 42149
rect 10781 42140 10793 42143
rect 10744 42112 10793 42140
rect 10744 42100 10750 42112
rect 10781 42109 10793 42112
rect 10827 42109 10839 42143
rect 11330 42140 11336 42152
rect 11291 42112 11336 42140
rect 10781 42103 10839 42109
rect 11330 42100 11336 42112
rect 11388 42100 11394 42152
rect 12989 42143 13047 42149
rect 12989 42109 13001 42143
rect 13035 42140 13047 42143
rect 13096 42140 13124 42316
rect 13906 42304 13912 42316
rect 13964 42344 13970 42356
rect 18046 42344 18052 42356
rect 13964 42316 18052 42344
rect 13964 42304 13970 42316
rect 18046 42304 18052 42316
rect 18104 42344 18110 42356
rect 18233 42347 18291 42353
rect 18233 42344 18245 42347
rect 18104 42316 18245 42344
rect 18104 42304 18110 42316
rect 18233 42313 18245 42316
rect 18279 42313 18291 42347
rect 18233 42307 18291 42313
rect 14369 42279 14427 42285
rect 14369 42245 14381 42279
rect 14415 42276 14427 42279
rect 15470 42276 15476 42288
rect 14415 42248 15476 42276
rect 14415 42245 14427 42248
rect 14369 42239 14427 42245
rect 15470 42236 15476 42248
rect 15528 42276 15534 42288
rect 15933 42279 15991 42285
rect 15933 42276 15945 42279
rect 15528 42248 15945 42276
rect 15528 42236 15534 42248
rect 15933 42245 15945 42248
rect 15979 42276 15991 42279
rect 16022 42276 16028 42288
rect 15979 42248 16028 42276
rect 15979 42245 15991 42248
rect 15933 42239 15991 42245
rect 16022 42236 16028 42248
rect 16080 42236 16086 42288
rect 13538 42208 13544 42220
rect 13499 42180 13544 42208
rect 13538 42168 13544 42180
rect 13596 42168 13602 42220
rect 15105 42211 15163 42217
rect 15105 42177 15117 42211
rect 15151 42208 15163 42211
rect 17034 42208 17040 42220
rect 15151 42180 17040 42208
rect 15151 42177 15163 42180
rect 15105 42171 15163 42177
rect 17034 42168 17040 42180
rect 17092 42168 17098 42220
rect 13035 42112 13124 42140
rect 13173 42143 13231 42149
rect 13035 42109 13047 42112
rect 12989 42103 13047 42109
rect 13173 42109 13185 42143
rect 13219 42140 13231 42143
rect 14274 42140 14280 42152
rect 13219 42112 14280 42140
rect 13219 42109 13231 42112
rect 13173 42103 13231 42109
rect 14274 42100 14280 42112
rect 14332 42100 14338 42152
rect 14642 42140 14648 42152
rect 14603 42112 14648 42140
rect 14642 42100 14648 42112
rect 14700 42100 14706 42152
rect 16206 42140 16212 42152
rect 16167 42112 16212 42140
rect 16206 42100 16212 42112
rect 16264 42100 16270 42152
rect 17862 42100 17868 42152
rect 17920 42140 17926 42152
rect 18049 42143 18107 42149
rect 18049 42140 18061 42143
rect 17920 42112 18061 42140
rect 17920 42100 17926 42112
rect 18049 42109 18061 42112
rect 18095 42109 18107 42143
rect 18049 42103 18107 42109
rect 14550 42072 14556 42084
rect 14511 42044 14556 42072
rect 14550 42032 14556 42044
rect 14608 42032 14614 42084
rect 16114 42072 16120 42084
rect 16075 42044 16120 42072
rect 16114 42032 16120 42044
rect 16172 42032 16178 42084
rect 16666 42072 16672 42084
rect 16627 42044 16672 42072
rect 16666 42032 16672 42044
rect 16724 42032 16730 42084
rect 1104 41914 24840 41936
rect 1104 41862 8912 41914
rect 8964 41862 8976 41914
rect 9028 41862 9040 41914
rect 9092 41862 9104 41914
rect 9156 41862 16843 41914
rect 16895 41862 16907 41914
rect 16959 41862 16971 41914
rect 17023 41862 17035 41914
rect 17087 41862 24840 41914
rect 1104 41840 24840 41862
rect 4246 41760 4252 41812
rect 4304 41800 4310 41812
rect 5629 41803 5687 41809
rect 5629 41800 5641 41803
rect 4304 41772 5641 41800
rect 4304 41760 4310 41772
rect 5629 41769 5641 41772
rect 5675 41769 5687 41803
rect 5629 41763 5687 41769
rect 14550 41760 14556 41812
rect 14608 41800 14614 41812
rect 15657 41803 15715 41809
rect 15657 41800 15669 41803
rect 14608 41772 15669 41800
rect 14608 41760 14614 41772
rect 15657 41769 15669 41772
rect 15703 41769 15715 41803
rect 15657 41763 15715 41769
rect 1946 41624 1952 41676
rect 2004 41664 2010 41676
rect 2590 41664 2596 41676
rect 2004 41636 2596 41664
rect 2004 41624 2010 41636
rect 2590 41624 2596 41636
rect 2648 41624 2654 41676
rect 2777 41667 2835 41673
rect 2777 41633 2789 41667
rect 2823 41664 2835 41667
rect 4264 41664 4292 41760
rect 7742 41732 7748 41744
rect 7703 41704 7748 41732
rect 7742 41692 7748 41704
rect 7800 41692 7806 41744
rect 9490 41692 9496 41744
rect 9548 41732 9554 41744
rect 9861 41735 9919 41741
rect 9861 41732 9873 41735
rect 9548 41704 9873 41732
rect 9548 41692 9554 41704
rect 9861 41701 9873 41704
rect 9907 41701 9919 41735
rect 9861 41695 9919 41701
rect 11330 41692 11336 41744
rect 11388 41732 11394 41744
rect 11388 41704 12204 41732
rect 11388 41692 11394 41704
rect 2823 41636 4292 41664
rect 2823 41633 2835 41636
rect 2777 41627 2835 41633
rect 7466 41624 7472 41676
rect 7524 41664 7530 41676
rect 7837 41667 7895 41673
rect 7837 41664 7849 41667
rect 7524 41636 7849 41664
rect 7524 41624 7530 41636
rect 7837 41633 7849 41636
rect 7883 41633 7895 41667
rect 7837 41627 7895 41633
rect 9674 41624 9680 41676
rect 9732 41664 9738 41676
rect 9953 41667 10011 41673
rect 9953 41664 9965 41667
rect 9732 41636 9965 41664
rect 9732 41624 9738 41636
rect 9953 41633 9965 41636
rect 9999 41633 10011 41667
rect 11790 41664 11796 41676
rect 11751 41636 11796 41664
rect 9953 41627 10011 41633
rect 11790 41624 11796 41636
rect 11848 41624 11854 41676
rect 12176 41673 12204 41704
rect 18322 41692 18328 41744
rect 18380 41732 18386 41744
rect 18417 41735 18475 41741
rect 18417 41732 18429 41735
rect 18380 41704 18429 41732
rect 18380 41692 18386 41704
rect 18417 41701 18429 41704
rect 18463 41732 18475 41735
rect 21174 41732 21180 41744
rect 18463 41704 21180 41732
rect 18463 41701 18475 41704
rect 18417 41695 18475 41701
rect 21174 41692 21180 41704
rect 21232 41692 21238 41744
rect 12161 41667 12219 41673
rect 12161 41633 12173 41667
rect 12207 41633 12219 41667
rect 12161 41627 12219 41633
rect 13170 41624 13176 41676
rect 13228 41664 13234 41676
rect 13449 41667 13507 41673
rect 13449 41664 13461 41667
rect 13228 41636 13461 41664
rect 13228 41624 13234 41636
rect 13449 41633 13461 41636
rect 13495 41633 13507 41667
rect 13449 41627 13507 41633
rect 13909 41667 13967 41673
rect 13909 41633 13921 41667
rect 13955 41633 13967 41667
rect 13909 41627 13967 41633
rect 14369 41667 14427 41673
rect 14369 41633 14381 41667
rect 14415 41664 14427 41667
rect 14458 41664 14464 41676
rect 14415 41636 14464 41664
rect 14415 41633 14427 41636
rect 14369 41627 14427 41633
rect 3145 41599 3203 41605
rect 3145 41565 3157 41599
rect 3191 41596 3203 41599
rect 4062 41596 4068 41608
rect 3191 41568 4068 41596
rect 3191 41565 3203 41568
rect 3145 41559 3203 41565
rect 4062 41556 4068 41568
rect 4120 41556 4126 41608
rect 4154 41556 4160 41608
rect 4212 41596 4218 41608
rect 4249 41599 4307 41605
rect 4249 41596 4261 41599
rect 4212 41568 4261 41596
rect 4212 41556 4218 41568
rect 4249 41565 4261 41568
rect 4295 41565 4307 41599
rect 4522 41596 4528 41608
rect 4483 41568 4528 41596
rect 4249 41559 4307 41565
rect 4522 41556 4528 41568
rect 4580 41556 4586 41608
rect 6914 41556 6920 41608
rect 6972 41596 6978 41608
rect 7190 41596 7196 41608
rect 6972 41568 7196 41596
rect 6972 41556 6978 41568
rect 7190 41556 7196 41568
rect 7248 41596 7254 41608
rect 7561 41599 7619 41605
rect 7561 41596 7573 41599
rect 7248 41568 7573 41596
rect 7248 41556 7254 41568
rect 7561 41565 7573 41568
rect 7607 41596 7619 41599
rect 11977 41599 12035 41605
rect 7607 41568 9720 41596
rect 7607 41565 7619 41568
rect 7561 41559 7619 41565
rect 9692 41537 9720 41568
rect 11977 41565 11989 41599
rect 12023 41596 12035 41599
rect 12526 41596 12532 41608
rect 12023 41568 12532 41596
rect 12023 41565 12035 41568
rect 11977 41559 12035 41565
rect 12526 41556 12532 41568
rect 12584 41556 12590 41608
rect 9677 41531 9735 41537
rect 9677 41497 9689 41531
rect 9723 41497 9735 41531
rect 13924 41528 13952 41627
rect 14458 41624 14464 41636
rect 14516 41624 14522 41676
rect 15378 41664 15384 41676
rect 15339 41636 15384 41664
rect 15378 41624 15384 41636
rect 15436 41624 15442 41676
rect 15562 41664 15568 41676
rect 15523 41636 15568 41664
rect 15562 41624 15568 41636
rect 15620 41624 15626 41676
rect 16666 41624 16672 41676
rect 16724 41664 16730 41676
rect 17037 41667 17095 41673
rect 17037 41664 17049 41667
rect 16724 41636 17049 41664
rect 16724 41624 16730 41636
rect 17037 41633 17049 41636
rect 17083 41633 17095 41667
rect 17037 41627 17095 41633
rect 14001 41599 14059 41605
rect 14001 41565 14013 41599
rect 14047 41596 14059 41599
rect 14642 41596 14648 41608
rect 14047 41568 14648 41596
rect 14047 41565 14059 41568
rect 14001 41559 14059 41565
rect 14642 41556 14648 41568
rect 14700 41556 14706 41608
rect 16574 41556 16580 41608
rect 16632 41596 16638 41608
rect 16761 41599 16819 41605
rect 16761 41596 16773 41599
rect 16632 41568 16773 41596
rect 16632 41556 16638 41568
rect 16761 41565 16773 41568
rect 16807 41565 16819 41599
rect 16761 41559 16819 41565
rect 14274 41528 14280 41540
rect 13924 41500 14280 41528
rect 9677 41491 9735 41497
rect 14274 41488 14280 41500
rect 14332 41488 14338 41540
rect 14826 41488 14832 41540
rect 14884 41488 14890 41540
rect 4154 41420 4160 41472
rect 4212 41460 4218 41472
rect 4430 41460 4436 41472
rect 4212 41432 4436 41460
rect 4212 41420 4218 41432
rect 4430 41420 4436 41432
rect 4488 41420 4494 41472
rect 7834 41420 7840 41472
rect 7892 41460 7898 41472
rect 8021 41463 8079 41469
rect 8021 41460 8033 41463
rect 7892 41432 8033 41460
rect 7892 41420 7898 41432
rect 8021 41429 8033 41432
rect 8067 41429 8079 41463
rect 8021 41423 8079 41429
rect 9950 41420 9956 41472
rect 10008 41460 10014 41472
rect 10137 41463 10195 41469
rect 10137 41460 10149 41463
rect 10008 41432 10149 41460
rect 10008 41420 10014 41432
rect 10137 41429 10149 41432
rect 10183 41429 10195 41463
rect 10137 41423 10195 41429
rect 13265 41463 13323 41469
rect 13265 41429 13277 41463
rect 13311 41460 13323 41463
rect 14844 41460 14872 41488
rect 13311 41432 14872 41460
rect 13311 41429 13323 41432
rect 13265 41423 13323 41429
rect 1104 41370 24840 41392
rect 1104 41318 4947 41370
rect 4999 41318 5011 41370
rect 5063 41318 5075 41370
rect 5127 41318 5139 41370
rect 5191 41318 12878 41370
rect 12930 41318 12942 41370
rect 12994 41318 13006 41370
rect 13058 41318 13070 41370
rect 13122 41318 20808 41370
rect 20860 41318 20872 41370
rect 20924 41318 20936 41370
rect 20988 41318 21000 41370
rect 21052 41318 24840 41370
rect 1104 41296 24840 41318
rect 3418 41256 3424 41268
rect 3379 41228 3424 41256
rect 3418 41216 3424 41228
rect 3476 41216 3482 41268
rect 4525 41259 4583 41265
rect 4525 41225 4537 41259
rect 4571 41256 4583 41259
rect 4614 41256 4620 41268
rect 4571 41228 4620 41256
rect 4571 41225 4583 41228
rect 4525 41219 4583 41225
rect 4614 41216 4620 41228
rect 4672 41216 4678 41268
rect 7374 41216 7380 41268
rect 7432 41256 7438 41268
rect 8389 41259 8447 41265
rect 8389 41256 8401 41259
rect 7432 41228 8401 41256
rect 7432 41216 7438 41228
rect 8389 41225 8401 41228
rect 8435 41225 8447 41259
rect 8389 41219 8447 41225
rect 9861 41259 9919 41265
rect 9861 41225 9873 41259
rect 9907 41256 9919 41259
rect 12710 41256 12716 41268
rect 9907 41228 12716 41256
rect 9907 41225 9919 41228
rect 9861 41219 9919 41225
rect 12710 41216 12716 41228
rect 12768 41216 12774 41268
rect 12897 41259 12955 41265
rect 12897 41225 12909 41259
rect 12943 41256 12955 41259
rect 17126 41256 17132 41268
rect 12943 41228 17132 41256
rect 12943 41225 12955 41228
rect 12897 41219 12955 41225
rect 17126 41216 17132 41228
rect 17184 41216 17190 41268
rect 16206 41148 16212 41200
rect 16264 41148 16270 41200
rect 4522 41080 4528 41132
rect 4580 41120 4586 41132
rect 5261 41123 5319 41129
rect 5261 41120 5273 41123
rect 4580 41092 5273 41120
rect 4580 41080 4586 41092
rect 5261 41089 5273 41092
rect 5307 41089 5319 41123
rect 5261 41083 5319 41089
rect 6822 41080 6828 41132
rect 6880 41120 6886 41132
rect 11149 41123 11207 41129
rect 6880 41092 9720 41120
rect 6880 41080 6886 41092
rect 2958 41052 2964 41064
rect 2919 41024 2964 41052
rect 2958 41012 2964 41024
rect 3016 41012 3022 41064
rect 3142 41052 3148 41064
rect 3103 41024 3148 41052
rect 3142 41012 3148 41024
rect 3200 41012 3206 41064
rect 3237 41055 3295 41061
rect 3237 41021 3249 41055
rect 3283 41052 3295 41055
rect 3694 41052 3700 41064
rect 3283 41024 3700 41052
rect 3283 41021 3295 41024
rect 3237 41015 3295 41021
rect 3694 41012 3700 41024
rect 3752 41012 3758 41064
rect 4798 41052 4804 41064
rect 4759 41024 4804 41052
rect 4798 41012 4804 41024
rect 4856 41012 4862 41064
rect 7006 41052 7012 41064
rect 6967 41024 7012 41052
rect 7006 41012 7012 41024
rect 7064 41012 7070 41064
rect 7282 41052 7288 41064
rect 7243 41024 7288 41052
rect 7282 41012 7288 41024
rect 7340 41012 7346 41064
rect 9692 41061 9720 41092
rect 11149 41089 11161 41123
rect 11195 41120 11207 41123
rect 12618 41120 12624 41132
rect 11195 41092 12624 41120
rect 11195 41089 11207 41092
rect 11149 41083 11207 41089
rect 12618 41080 12624 41092
rect 12676 41080 12682 41132
rect 14737 41123 14795 41129
rect 14737 41089 14749 41123
rect 14783 41120 14795 41123
rect 16224 41120 16252 41148
rect 14783 41092 16252 41120
rect 14783 41089 14795 41092
rect 14737 41083 14795 41089
rect 9677 41055 9735 41061
rect 9677 41021 9689 41055
rect 9723 41052 9735 41055
rect 9858 41052 9864 41064
rect 9723 41024 9864 41052
rect 9723 41021 9735 41024
rect 9677 41015 9735 41021
rect 9858 41012 9864 41024
rect 9916 41012 9922 41064
rect 10965 41055 11023 41061
rect 10965 41021 10977 41055
rect 11011 41052 11023 41055
rect 11054 41052 11060 41064
rect 11011 41024 11060 41052
rect 11011 41021 11023 41024
rect 10965 41015 11023 41021
rect 11054 41012 11060 41024
rect 11112 41012 11118 41064
rect 11330 41012 11336 41064
rect 11388 41052 11394 41064
rect 11514 41052 11520 41064
rect 11388 41024 11520 41052
rect 11388 41012 11394 41024
rect 11514 41012 11520 41024
rect 11572 41012 11578 41064
rect 13081 41055 13139 41061
rect 13081 41021 13093 41055
rect 13127 41052 13139 41055
rect 13262 41052 13268 41064
rect 13127 41024 13268 41052
rect 13127 41021 13139 41024
rect 13081 41015 13139 41021
rect 13262 41012 13268 41024
rect 13320 41012 13326 41064
rect 13541 41055 13599 41061
rect 13541 41021 13553 41055
rect 13587 41021 13599 41055
rect 14366 41052 14372 41064
rect 14327 41024 14372 41052
rect 13541 41015 13599 41021
rect 4062 40944 4068 40996
rect 4120 40984 4126 40996
rect 4709 40987 4767 40993
rect 4709 40984 4721 40987
rect 4120 40956 4721 40984
rect 4120 40944 4126 40956
rect 4709 40953 4721 40956
rect 4755 40953 4767 40987
rect 9876 40984 9904 41012
rect 11146 40984 11152 40996
rect 9876 40956 11152 40984
rect 4709 40947 4767 40953
rect 11146 40944 11152 40956
rect 11204 40944 11210 40996
rect 13556 40984 13584 41015
rect 14366 41012 14372 41024
rect 14424 41012 14430 41064
rect 14458 41012 14464 41064
rect 14516 41052 14522 41064
rect 14921 41055 14979 41061
rect 14921 41052 14933 41055
rect 14516 41024 14933 41052
rect 14516 41012 14522 41024
rect 14921 41021 14933 41024
rect 14967 41021 14979 41055
rect 16022 41052 16028 41064
rect 15983 41024 16028 41052
rect 14921 41015 14979 41021
rect 16022 41012 16028 41024
rect 16080 41012 16086 41064
rect 16206 41052 16212 41064
rect 16167 41024 16212 41052
rect 16206 41012 16212 41024
rect 16264 41012 16270 41064
rect 14476 40984 14504 41012
rect 16114 40984 16120 40996
rect 13556 40956 14504 40984
rect 16075 40956 16120 40984
rect 16114 40944 16120 40956
rect 16172 40944 16178 40996
rect 16666 40984 16672 40996
rect 16627 40956 16672 40984
rect 16666 40944 16672 40956
rect 16724 40944 16730 40996
rect 1104 40826 24840 40848
rect 1104 40774 8912 40826
rect 8964 40774 8976 40826
rect 9028 40774 9040 40826
rect 9092 40774 9104 40826
rect 9156 40774 16843 40826
rect 16895 40774 16907 40826
rect 16959 40774 16971 40826
rect 17023 40774 17035 40826
rect 17087 40774 24840 40826
rect 1104 40752 24840 40774
rect 3053 40715 3111 40721
rect 3053 40681 3065 40715
rect 3099 40712 3111 40715
rect 4154 40712 4160 40724
rect 3099 40684 4160 40712
rect 3099 40681 3111 40684
rect 3053 40675 3111 40681
rect 4154 40672 4160 40684
rect 4212 40672 4218 40724
rect 18141 40715 18199 40721
rect 18141 40712 18153 40715
rect 15580 40684 18153 40712
rect 5902 40604 5908 40656
rect 5960 40644 5966 40656
rect 6641 40647 6699 40653
rect 6641 40644 6653 40647
rect 5960 40616 6653 40644
rect 5960 40604 5966 40616
rect 6641 40613 6653 40616
rect 6687 40613 6699 40647
rect 6641 40607 6699 40613
rect 7193 40647 7251 40653
rect 7193 40613 7205 40647
rect 7239 40644 7251 40647
rect 7282 40644 7288 40656
rect 7239 40616 7288 40644
rect 7239 40613 7251 40616
rect 7193 40607 7251 40613
rect 7282 40604 7288 40616
rect 7340 40604 7346 40656
rect 15378 40644 15384 40656
rect 15339 40616 15384 40644
rect 15378 40604 15384 40616
rect 15436 40604 15442 40656
rect 1765 40579 1823 40585
rect 1765 40545 1777 40579
rect 1811 40576 1823 40579
rect 2869 40579 2927 40585
rect 2869 40576 2881 40579
rect 1811 40548 2881 40576
rect 1811 40545 1823 40548
rect 1765 40539 1823 40545
rect 2869 40545 2881 40548
rect 2915 40576 2927 40579
rect 3142 40576 3148 40588
rect 2915 40548 3148 40576
rect 2915 40545 2927 40548
rect 2869 40539 2927 40545
rect 3142 40536 3148 40548
rect 3200 40536 3206 40588
rect 4430 40576 4436 40588
rect 4391 40548 4436 40576
rect 4430 40536 4436 40548
rect 4488 40536 4494 40588
rect 4798 40576 4804 40588
rect 4759 40548 4804 40576
rect 4798 40536 4804 40548
rect 4856 40536 4862 40588
rect 5169 40579 5227 40585
rect 5169 40545 5181 40579
rect 5215 40576 5227 40579
rect 5350 40576 5356 40588
rect 5215 40548 5356 40576
rect 5215 40545 5227 40548
rect 5169 40539 5227 40545
rect 5350 40536 5356 40548
rect 5408 40536 5414 40588
rect 6730 40576 6736 40588
rect 6691 40548 6736 40576
rect 6730 40536 6736 40548
rect 6788 40536 6794 40588
rect 8202 40576 8208 40588
rect 8163 40548 8208 40576
rect 8202 40536 8208 40548
rect 8260 40536 8266 40588
rect 8754 40576 8760 40588
rect 8715 40548 8760 40576
rect 8754 40536 8760 40548
rect 8812 40536 8818 40588
rect 9858 40576 9864 40588
rect 9819 40548 9864 40576
rect 9858 40536 9864 40548
rect 9916 40536 9922 40588
rect 11146 40576 11152 40588
rect 11107 40548 11152 40576
rect 11146 40536 11152 40548
rect 11204 40536 11210 40588
rect 11514 40576 11520 40588
rect 11475 40548 11520 40576
rect 11514 40536 11520 40548
rect 11572 40536 11578 40588
rect 12434 40536 12440 40588
rect 12492 40576 12498 40588
rect 15580 40585 15608 40684
rect 18141 40681 18153 40684
rect 18187 40712 18199 40715
rect 18506 40712 18512 40724
rect 18187 40684 18512 40712
rect 18187 40681 18199 40684
rect 18141 40675 18199 40681
rect 18506 40672 18512 40684
rect 18564 40672 18570 40724
rect 15933 40647 15991 40653
rect 15933 40613 15945 40647
rect 15979 40644 15991 40647
rect 16114 40644 16120 40656
rect 15979 40616 16120 40644
rect 15979 40613 15991 40616
rect 15933 40607 15991 40613
rect 16114 40604 16120 40616
rect 16172 40604 16178 40656
rect 12529 40579 12587 40585
rect 12529 40576 12541 40579
rect 12492 40548 12541 40576
rect 12492 40536 12498 40548
rect 12529 40545 12541 40548
rect 12575 40545 12587 40579
rect 12529 40539 12587 40545
rect 15565 40579 15623 40585
rect 15565 40545 15577 40579
rect 15611 40545 15623 40579
rect 15565 40539 15623 40545
rect 16666 40536 16672 40588
rect 16724 40576 16730 40588
rect 17037 40579 17095 40585
rect 17037 40576 17049 40579
rect 16724 40548 17049 40576
rect 16724 40536 16730 40548
rect 17037 40545 17049 40548
rect 17083 40545 17095 40579
rect 17037 40539 17095 40545
rect 6457 40511 6515 40517
rect 6457 40477 6469 40511
rect 6503 40508 6515 40511
rect 7190 40508 7196 40520
rect 6503 40480 7196 40508
rect 6503 40477 6515 40480
rect 6457 40471 6515 40477
rect 7190 40468 7196 40480
rect 7248 40468 7254 40520
rect 8389 40511 8447 40517
rect 8389 40477 8401 40511
rect 8435 40508 8447 40511
rect 9674 40508 9680 40520
rect 8435 40480 9680 40508
rect 8435 40477 8447 40480
rect 8389 40471 8447 40477
rect 9674 40468 9680 40480
rect 9732 40468 9738 40520
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 12805 40511 12863 40517
rect 12805 40508 12817 40511
rect 12768 40480 12817 40508
rect 12768 40468 12774 40480
rect 12805 40477 12817 40480
rect 12851 40477 12863 40511
rect 12805 40471 12863 40477
rect 16574 40468 16580 40520
rect 16632 40508 16638 40520
rect 16761 40511 16819 40517
rect 16761 40508 16773 40511
rect 16632 40480 16773 40508
rect 16632 40468 16638 40480
rect 16761 40477 16773 40480
rect 16807 40477 16819 40511
rect 16761 40471 16819 40477
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 10042 40372 10048 40384
rect 10003 40344 10048 40372
rect 10042 40332 10048 40344
rect 10100 40332 10106 40384
rect 11057 40375 11115 40381
rect 11057 40341 11069 40375
rect 11103 40372 11115 40375
rect 13814 40372 13820 40384
rect 11103 40344 13820 40372
rect 11103 40341 11115 40344
rect 11057 40335 11115 40341
rect 13814 40332 13820 40344
rect 13872 40332 13878 40384
rect 13906 40332 13912 40384
rect 13964 40372 13970 40384
rect 13964 40344 14009 40372
rect 13964 40332 13970 40344
rect 14918 40332 14924 40384
rect 14976 40372 14982 40384
rect 17862 40372 17868 40384
rect 14976 40344 17868 40372
rect 14976 40332 14982 40344
rect 17862 40332 17868 40344
rect 17920 40332 17926 40384
rect 1104 40282 24840 40304
rect 1104 40230 4947 40282
rect 4999 40230 5011 40282
rect 5063 40230 5075 40282
rect 5127 40230 5139 40282
rect 5191 40230 12878 40282
rect 12930 40230 12942 40282
rect 12994 40230 13006 40282
rect 13058 40230 13070 40282
rect 13122 40230 20808 40282
rect 20860 40230 20872 40282
rect 20924 40230 20936 40282
rect 20988 40230 21000 40282
rect 21052 40230 24840 40282
rect 1104 40208 24840 40230
rect 4893 40171 4951 40177
rect 4893 40137 4905 40171
rect 4939 40168 4951 40171
rect 5258 40168 5264 40180
rect 4939 40140 5264 40168
rect 4939 40137 4951 40140
rect 4893 40131 4951 40137
rect 5258 40128 5264 40140
rect 5316 40128 5322 40180
rect 7745 40171 7803 40177
rect 7745 40137 7757 40171
rect 7791 40168 7803 40171
rect 9214 40168 9220 40180
rect 7791 40140 9220 40168
rect 7791 40137 7803 40140
rect 7745 40131 7803 40137
rect 9214 40128 9220 40140
rect 9272 40128 9278 40180
rect 9309 40171 9367 40177
rect 9309 40137 9321 40171
rect 9355 40168 9367 40171
rect 10410 40168 10416 40180
rect 9355 40140 10416 40168
rect 9355 40137 9367 40140
rect 9309 40131 9367 40137
rect 10410 40128 10416 40140
rect 10468 40128 10474 40180
rect 12710 40128 12716 40180
rect 12768 40168 12774 40180
rect 12897 40171 12955 40177
rect 12897 40168 12909 40171
rect 12768 40140 12909 40168
rect 12768 40128 12774 40140
rect 12897 40137 12909 40140
rect 12943 40137 12955 40171
rect 12897 40131 12955 40137
rect 15105 40171 15163 40177
rect 15105 40137 15117 40171
rect 15151 40168 15163 40171
rect 15378 40168 15384 40180
rect 15151 40140 15384 40168
rect 15151 40137 15163 40140
rect 15105 40131 15163 40137
rect 15378 40128 15384 40140
rect 15436 40128 15442 40180
rect 18325 40171 18383 40177
rect 18325 40168 18337 40171
rect 16592 40140 18337 40168
rect 11422 40100 11428 40112
rect 11164 40072 11428 40100
rect 3510 40032 3516 40044
rect 3471 40004 3516 40032
rect 3510 39992 3516 40004
rect 3568 39992 3574 40044
rect 6362 39992 6368 40044
rect 6420 40032 6426 40044
rect 11164 40041 11192 40072
rect 11422 40060 11428 40072
rect 11480 40060 11486 40112
rect 11149 40035 11207 40041
rect 6420 40004 10364 40032
rect 6420 39992 6426 40004
rect 2133 39967 2191 39973
rect 2133 39933 2145 39967
rect 2179 39933 2191 39967
rect 2133 39927 2191 39933
rect 2409 39967 2467 39973
rect 2409 39933 2421 39967
rect 2455 39964 2467 39967
rect 2498 39964 2504 39976
rect 2455 39936 2504 39964
rect 2455 39933 2467 39936
rect 2409 39927 2467 39933
rect 2148 39828 2176 39927
rect 2498 39924 2504 39936
rect 2556 39924 2562 39976
rect 4798 39964 4804 39976
rect 4759 39936 4804 39964
rect 4798 39924 4804 39936
rect 4856 39924 4862 39976
rect 5350 39964 5356 39976
rect 5311 39936 5356 39964
rect 5350 39924 5356 39936
rect 5408 39924 5414 39976
rect 6549 39967 6607 39973
rect 6549 39933 6561 39967
rect 6595 39933 6607 39967
rect 6549 39927 6607 39933
rect 7929 39967 7987 39973
rect 7929 39933 7941 39967
rect 7975 39933 7987 39967
rect 7929 39927 7987 39933
rect 8389 39967 8447 39973
rect 8389 39933 8401 39967
rect 8435 39964 8447 39967
rect 8754 39964 8760 39976
rect 8435 39936 8760 39964
rect 8435 39933 8447 39936
rect 8389 39927 8447 39933
rect 6564 39896 6592 39927
rect 7742 39896 7748 39908
rect 6564 39868 7748 39896
rect 7742 39856 7748 39868
rect 7800 39856 7806 39908
rect 7944 39896 7972 39927
rect 8754 39924 8760 39936
rect 8812 39924 8818 39976
rect 9214 39964 9220 39976
rect 9175 39936 9220 39964
rect 9214 39924 9220 39936
rect 9272 39924 9278 39976
rect 9858 39964 9864 39976
rect 9819 39936 9864 39964
rect 9858 39924 9864 39936
rect 9916 39924 9922 39976
rect 10226 39896 10232 39908
rect 7944 39868 10232 39896
rect 10226 39856 10232 39868
rect 10284 39856 10290 39908
rect 10336 39896 10364 40004
rect 11149 40001 11161 40035
rect 11195 40001 11207 40035
rect 11149 39995 11207 40001
rect 13909 40035 13967 40041
rect 13909 40001 13921 40035
rect 13955 40032 13967 40035
rect 15194 40032 15200 40044
rect 13955 40004 15200 40032
rect 13955 40001 13967 40004
rect 13909 39995 13967 40001
rect 15194 39992 15200 40004
rect 15252 39992 15258 40044
rect 16592 40032 16620 40140
rect 18325 40137 18337 40140
rect 18371 40137 18383 40171
rect 18325 40131 18383 40137
rect 16224 40004 16620 40032
rect 10962 39964 10968 39976
rect 10923 39936 10968 39964
rect 10962 39924 10968 39936
rect 11020 39924 11026 39976
rect 11422 39964 11428 39976
rect 11383 39936 11428 39964
rect 11422 39924 11428 39936
rect 11480 39924 11486 39976
rect 11606 39924 11612 39976
rect 11664 39964 11670 39976
rect 13449 39967 13507 39973
rect 13449 39964 13461 39967
rect 11664 39936 13461 39964
rect 11664 39924 11670 39936
rect 13449 39933 13461 39936
rect 13495 39933 13507 39967
rect 13449 39927 13507 39933
rect 13538 39924 13544 39976
rect 13596 39964 13602 39976
rect 13814 39964 13820 39976
rect 13596 39936 13641 39964
rect 13775 39936 13820 39964
rect 13596 39924 13602 39936
rect 13814 39924 13820 39936
rect 13872 39924 13878 39976
rect 14918 39964 14924 39976
rect 14879 39936 14924 39964
rect 14918 39924 14924 39936
rect 14976 39924 14982 39976
rect 16114 39964 16120 39976
rect 16075 39936 16120 39964
rect 16114 39924 16120 39936
rect 16172 39924 16178 39976
rect 16224 39973 16252 40004
rect 16209 39967 16267 39973
rect 16209 39933 16221 39967
rect 16255 39933 16267 39967
rect 16209 39927 16267 39933
rect 16298 39924 16304 39976
rect 16356 39964 16362 39976
rect 18049 39967 18107 39973
rect 18049 39964 18061 39967
rect 16356 39936 16401 39964
rect 16500 39936 18061 39964
rect 16356 39924 16362 39936
rect 14936 39896 14964 39924
rect 16500 39908 16528 39936
rect 18049 39933 18061 39936
rect 18095 39933 18107 39967
rect 18049 39927 18107 39933
rect 18233 39967 18291 39973
rect 18233 39933 18245 39967
rect 18279 39964 18291 39967
rect 18322 39964 18328 39976
rect 18279 39936 18328 39964
rect 18279 39933 18291 39936
rect 18233 39927 18291 39933
rect 18322 39924 18328 39936
rect 18380 39964 18386 39976
rect 22094 39964 22100 39976
rect 18380 39936 22100 39964
rect 18380 39924 18386 39936
rect 22094 39924 22100 39936
rect 22152 39924 22158 39976
rect 10336 39868 14964 39896
rect 15378 39856 15384 39908
rect 15436 39896 15442 39908
rect 16482 39896 16488 39908
rect 15436 39868 16488 39896
rect 15436 39856 15442 39868
rect 16482 39856 16488 39868
rect 16540 39856 16546 39908
rect 16666 39856 16672 39908
rect 16724 39896 16730 39908
rect 16761 39899 16819 39905
rect 16761 39896 16773 39899
rect 16724 39868 16773 39896
rect 16724 39856 16730 39868
rect 16761 39865 16773 39868
rect 16807 39865 16819 39899
rect 16761 39859 16819 39865
rect 4246 39828 4252 39840
rect 2148 39800 4252 39828
rect 4246 39788 4252 39800
rect 4304 39828 4310 39840
rect 5258 39828 5264 39840
rect 4304 39800 5264 39828
rect 4304 39788 4310 39800
rect 5258 39788 5264 39800
rect 5316 39828 5322 39840
rect 6365 39831 6423 39837
rect 6365 39828 6377 39831
rect 5316 39800 6377 39828
rect 5316 39788 5322 39800
rect 6365 39797 6377 39800
rect 6411 39797 6423 39831
rect 6365 39791 6423 39797
rect 1104 39738 24840 39760
rect 1104 39686 8912 39738
rect 8964 39686 8976 39738
rect 9028 39686 9040 39738
rect 9092 39686 9104 39738
rect 9156 39686 16843 39738
rect 16895 39686 16907 39738
rect 16959 39686 16971 39738
rect 17023 39686 17035 39738
rect 17087 39686 24840 39738
rect 1104 39664 24840 39686
rect 12069 39627 12127 39633
rect 12069 39593 12081 39627
rect 12115 39624 12127 39627
rect 13814 39624 13820 39636
rect 12115 39596 13820 39624
rect 12115 39593 12127 39596
rect 12069 39587 12127 39593
rect 13814 39584 13820 39596
rect 13872 39624 13878 39636
rect 18322 39624 18328 39636
rect 13872 39596 15424 39624
rect 18283 39596 18328 39624
rect 13872 39584 13878 39596
rect 2682 39516 2688 39568
rect 2740 39556 2746 39568
rect 6733 39559 6791 39565
rect 2740 39528 6500 39556
rect 2740 39516 2746 39528
rect 2869 39491 2927 39497
rect 2869 39457 2881 39491
rect 2915 39457 2927 39491
rect 4614 39488 4620 39500
rect 4575 39460 4620 39488
rect 2869 39451 2927 39457
rect 2884 39352 2912 39451
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 4706 39448 4712 39500
rect 4764 39488 4770 39500
rect 4801 39491 4859 39497
rect 4801 39488 4813 39491
rect 4764 39460 4813 39488
rect 4764 39448 4770 39460
rect 4801 39457 4813 39460
rect 4847 39457 4859 39491
rect 4801 39451 4859 39457
rect 5169 39491 5227 39497
rect 5169 39457 5181 39491
rect 5215 39488 5227 39491
rect 5350 39488 5356 39500
rect 5215 39460 5356 39488
rect 5215 39457 5227 39460
rect 5169 39451 5227 39457
rect 5350 39448 5356 39460
rect 5408 39448 5414 39500
rect 6472 39497 6500 39528
rect 6733 39525 6745 39559
rect 6779 39556 6791 39559
rect 6822 39556 6828 39568
rect 6779 39528 6828 39556
rect 6779 39525 6791 39528
rect 6733 39519 6791 39525
rect 6822 39516 6828 39528
rect 6880 39516 6886 39568
rect 15396 39500 15424 39596
rect 18322 39584 18328 39596
rect 18380 39584 18386 39636
rect 6273 39491 6331 39497
rect 6273 39457 6285 39491
rect 6319 39457 6331 39491
rect 6273 39451 6331 39457
rect 6457 39491 6515 39497
rect 6457 39457 6469 39491
rect 6503 39457 6515 39491
rect 7742 39488 7748 39500
rect 7703 39460 7748 39488
rect 6457 39451 6515 39457
rect 6288 39420 6316 39451
rect 7742 39448 7748 39460
rect 7800 39448 7806 39500
rect 8205 39491 8263 39497
rect 8205 39457 8217 39491
rect 8251 39457 8263 39491
rect 8386 39488 8392 39500
rect 8347 39460 8392 39488
rect 8205 39451 8263 39457
rect 6546 39420 6552 39432
rect 6288 39392 6552 39420
rect 6546 39380 6552 39392
rect 6604 39380 6610 39432
rect 6362 39352 6368 39364
rect 2884 39324 6368 39352
rect 6362 39312 6368 39324
rect 6420 39312 6426 39364
rect 8220 39352 8248 39451
rect 8386 39448 8392 39460
rect 8444 39448 8450 39500
rect 8754 39488 8760 39500
rect 8667 39460 8760 39488
rect 8754 39448 8760 39460
rect 8812 39488 8818 39500
rect 9858 39488 9864 39500
rect 8812 39460 9864 39488
rect 8812 39448 8818 39460
rect 9858 39448 9864 39460
rect 9916 39448 9922 39500
rect 10505 39491 10563 39497
rect 10505 39457 10517 39491
rect 10551 39488 10563 39491
rect 10870 39488 10876 39500
rect 10551 39460 10876 39488
rect 10551 39457 10563 39460
rect 10505 39451 10563 39457
rect 10870 39448 10876 39460
rect 10928 39488 10934 39500
rect 12434 39488 12440 39500
rect 10928 39460 12440 39488
rect 10928 39448 10934 39460
rect 12434 39448 12440 39460
rect 12492 39448 12498 39500
rect 13170 39488 13176 39500
rect 13131 39460 13176 39488
rect 13170 39448 13176 39460
rect 13228 39448 13234 39500
rect 13909 39491 13967 39497
rect 13909 39457 13921 39491
rect 13955 39457 13967 39491
rect 13909 39451 13967 39457
rect 14369 39491 14427 39497
rect 14369 39457 14381 39491
rect 14415 39488 14427 39491
rect 14458 39488 14464 39500
rect 14415 39460 14464 39488
rect 14415 39457 14427 39460
rect 14369 39451 14427 39457
rect 10778 39420 10784 39432
rect 10739 39392 10784 39420
rect 10778 39380 10784 39392
rect 10836 39380 10842 39432
rect 8386 39352 8392 39364
rect 8220 39324 8392 39352
rect 8386 39312 8392 39324
rect 8444 39312 8450 39364
rect 12452 39352 12480 39448
rect 12618 39352 12624 39364
rect 12452 39324 12624 39352
rect 12618 39312 12624 39324
rect 12676 39352 12682 39364
rect 12989 39355 13047 39361
rect 12989 39352 13001 39355
rect 12676 39324 13001 39352
rect 12676 39312 12682 39324
rect 12989 39321 13001 39324
rect 13035 39321 13047 39355
rect 13924 39352 13952 39451
rect 14458 39448 14464 39460
rect 14516 39448 14522 39500
rect 15194 39448 15200 39500
rect 15252 39488 15258 39500
rect 15289 39491 15347 39497
rect 15289 39488 15301 39491
rect 15252 39460 15301 39488
rect 15252 39448 15258 39460
rect 15289 39457 15301 39460
rect 15335 39457 15347 39491
rect 15289 39451 15347 39457
rect 15378 39448 15384 39500
rect 15436 39488 15442 39500
rect 15473 39491 15531 39497
rect 15473 39488 15485 39491
rect 15436 39460 15485 39488
rect 15436 39448 15442 39460
rect 15473 39457 15485 39460
rect 15519 39457 15531 39491
rect 15473 39451 15531 39457
rect 16666 39448 16672 39500
rect 16724 39488 16730 39500
rect 17037 39491 17095 39497
rect 17037 39488 17049 39491
rect 16724 39460 17049 39488
rect 16724 39448 16730 39460
rect 17037 39457 17049 39460
rect 17083 39457 17095 39491
rect 17037 39451 17095 39457
rect 14001 39423 14059 39429
rect 14001 39389 14013 39423
rect 14047 39420 14059 39423
rect 15654 39420 15660 39432
rect 14047 39392 15660 39420
rect 14047 39389 14059 39392
rect 14001 39383 14059 39389
rect 15654 39380 15660 39392
rect 15712 39380 15718 39432
rect 16574 39380 16580 39432
rect 16632 39420 16638 39432
rect 16761 39423 16819 39429
rect 16761 39420 16773 39423
rect 16632 39392 16773 39420
rect 16632 39380 16638 39392
rect 16761 39389 16773 39392
rect 16807 39389 16819 39423
rect 16761 39383 16819 39389
rect 14826 39352 14832 39364
rect 13924 39324 14832 39352
rect 12989 39315 13047 39321
rect 14826 39312 14832 39324
rect 14884 39312 14890 39364
rect 3053 39287 3111 39293
rect 3053 39253 3065 39287
rect 3099 39284 3111 39287
rect 4522 39284 4528 39296
rect 3099 39256 4528 39284
rect 3099 39253 3111 39256
rect 3053 39247 3111 39253
rect 4522 39244 4528 39256
rect 4580 39244 4586 39296
rect 7006 39244 7012 39296
rect 7064 39284 7070 39296
rect 7561 39287 7619 39293
rect 7561 39284 7573 39287
rect 7064 39256 7573 39284
rect 7064 39244 7070 39256
rect 7561 39253 7573 39256
rect 7607 39284 7619 39287
rect 7834 39284 7840 39296
rect 7607 39256 7840 39284
rect 7607 39253 7619 39256
rect 7561 39247 7619 39253
rect 7834 39244 7840 39256
rect 7892 39244 7898 39296
rect 14090 39244 14096 39296
rect 14148 39284 14154 39296
rect 15565 39287 15623 39293
rect 15565 39284 15577 39287
rect 14148 39256 15577 39284
rect 14148 39244 14154 39256
rect 15565 39253 15577 39256
rect 15611 39253 15623 39287
rect 15565 39247 15623 39253
rect 1104 39194 24840 39216
rect 1104 39142 4947 39194
rect 4999 39142 5011 39194
rect 5063 39142 5075 39194
rect 5127 39142 5139 39194
rect 5191 39142 12878 39194
rect 12930 39142 12942 39194
rect 12994 39142 13006 39194
rect 13058 39142 13070 39194
rect 13122 39142 20808 39194
rect 20860 39142 20872 39194
rect 20924 39142 20936 39194
rect 20988 39142 21000 39194
rect 21052 39142 24840 39194
rect 1104 39120 24840 39142
rect 2498 39080 2504 39092
rect 2459 39052 2504 39080
rect 2498 39040 2504 39052
rect 2556 39040 2562 39092
rect 3694 39080 3700 39092
rect 3655 39052 3700 39080
rect 3694 39040 3700 39052
rect 3752 39040 3758 39092
rect 11425 39083 11483 39089
rect 11425 39049 11437 39083
rect 11471 39080 11483 39083
rect 11606 39080 11612 39092
rect 11471 39052 11612 39080
rect 11471 39049 11483 39052
rect 11425 39043 11483 39049
rect 11606 39040 11612 39052
rect 11664 39040 11670 39092
rect 9582 38972 9588 39024
rect 9640 39012 9646 39024
rect 10042 39012 10048 39024
rect 9640 38984 10048 39012
rect 9640 38972 9646 38984
rect 10042 38972 10048 38984
rect 10100 39012 10106 39024
rect 12066 39012 12072 39024
rect 10100 38984 12072 39012
rect 10100 38972 10106 38984
rect 12066 38972 12072 38984
rect 12124 38972 12130 39024
rect 2041 38947 2099 38953
rect 2041 38913 2053 38947
rect 2087 38944 2099 38947
rect 2406 38944 2412 38956
rect 2087 38916 2412 38944
rect 2087 38913 2099 38916
rect 2041 38907 2099 38913
rect 2406 38904 2412 38916
rect 2464 38904 2470 38956
rect 4522 38944 4528 38956
rect 4356 38916 4528 38944
rect 2317 38879 2375 38885
rect 2317 38845 2329 38879
rect 2363 38876 2375 38879
rect 3418 38876 3424 38888
rect 2363 38848 3424 38876
rect 2363 38845 2375 38848
rect 2317 38839 2375 38845
rect 3418 38836 3424 38848
rect 3476 38836 3482 38888
rect 3694 38876 3700 38888
rect 3655 38848 3700 38876
rect 3694 38836 3700 38848
rect 3752 38836 3758 38888
rect 4356 38885 4384 38916
rect 4522 38904 4528 38916
rect 4580 38944 4586 38956
rect 5350 38944 5356 38956
rect 4580 38916 5356 38944
rect 4580 38904 4586 38916
rect 5350 38904 5356 38916
rect 5408 38904 5414 38956
rect 5534 38944 5540 38956
rect 5495 38916 5540 38944
rect 5534 38904 5540 38916
rect 5592 38904 5598 38956
rect 7466 38944 7472 38956
rect 7427 38916 7472 38944
rect 7466 38904 7472 38916
rect 7524 38904 7530 38956
rect 10137 38947 10195 38953
rect 10137 38913 10149 38947
rect 10183 38944 10195 38947
rect 10594 38944 10600 38956
rect 10183 38916 10600 38944
rect 10183 38913 10195 38916
rect 10137 38907 10195 38913
rect 10594 38904 10600 38916
rect 10652 38904 10658 38956
rect 12618 38944 12624 38956
rect 12579 38916 12624 38944
rect 12618 38904 12624 38916
rect 12676 38904 12682 38956
rect 15473 38947 15531 38953
rect 15473 38913 15485 38947
rect 15519 38944 15531 38947
rect 16206 38944 16212 38956
rect 15519 38916 16212 38944
rect 15519 38913 15531 38916
rect 15473 38907 15531 38913
rect 16206 38904 16212 38916
rect 16264 38904 16270 38956
rect 4341 38879 4399 38885
rect 4341 38845 4353 38879
rect 4387 38845 4399 38879
rect 4341 38839 4399 38845
rect 5445 38879 5503 38885
rect 5445 38845 5457 38879
rect 5491 38845 5503 38879
rect 5902 38876 5908 38888
rect 5863 38848 5908 38876
rect 5445 38839 5503 38845
rect 2225 38811 2283 38817
rect 2225 38777 2237 38811
rect 2271 38808 2283 38811
rect 3510 38808 3516 38820
rect 2271 38780 3516 38808
rect 2271 38777 2283 38780
rect 2225 38771 2283 38777
rect 3510 38768 3516 38780
rect 3568 38768 3574 38820
rect 5460 38808 5488 38839
rect 5902 38836 5908 38848
rect 5960 38836 5966 38888
rect 6822 38836 6828 38888
rect 6880 38876 6886 38888
rect 7101 38879 7159 38885
rect 7101 38876 7113 38879
rect 6880 38848 7113 38876
rect 6880 38836 6886 38848
rect 7101 38845 7113 38848
rect 7147 38845 7159 38879
rect 7650 38876 7656 38888
rect 7611 38848 7656 38876
rect 7101 38839 7159 38845
rect 7650 38836 7656 38848
rect 7708 38836 7714 38888
rect 8665 38879 8723 38885
rect 8665 38845 8677 38879
rect 8711 38845 8723 38879
rect 8665 38839 8723 38845
rect 9769 38879 9827 38885
rect 9769 38845 9781 38879
rect 9815 38845 9827 38879
rect 9769 38839 9827 38845
rect 5810 38808 5816 38820
rect 5460 38780 5816 38808
rect 5810 38768 5816 38780
rect 5868 38768 5874 38820
rect 5534 38700 5540 38752
rect 5592 38740 5598 38752
rect 8680 38740 8708 38839
rect 9784 38808 9812 38839
rect 9858 38836 9864 38888
rect 9916 38876 9922 38888
rect 11330 38885 11336 38888
rect 10321 38879 10379 38885
rect 10321 38876 10333 38879
rect 9916 38848 10333 38876
rect 9916 38836 9922 38848
rect 10321 38845 10333 38848
rect 10367 38845 10379 38879
rect 11325 38876 11336 38885
rect 11291 38848 11336 38876
rect 10321 38839 10379 38845
rect 11325 38839 11336 38848
rect 11330 38836 11336 38839
rect 11388 38836 11394 38888
rect 12710 38836 12716 38888
rect 12768 38876 12774 38888
rect 12897 38879 12955 38885
rect 12897 38876 12909 38879
rect 12768 38848 12909 38876
rect 12768 38836 12774 38848
rect 12897 38845 12909 38848
rect 12943 38845 12955 38879
rect 12897 38839 12955 38845
rect 15381 38879 15439 38885
rect 15381 38845 15393 38879
rect 15427 38845 15439 38879
rect 15838 38876 15844 38888
rect 15799 38848 15844 38876
rect 15381 38839 15439 38845
rect 10594 38808 10600 38820
rect 9784 38780 10600 38808
rect 10594 38768 10600 38780
rect 10652 38768 10658 38820
rect 15396 38808 15424 38839
rect 15838 38836 15844 38848
rect 15896 38836 15902 38888
rect 16666 38876 16672 38888
rect 16627 38848 16672 38876
rect 16666 38836 16672 38848
rect 16724 38836 16730 38888
rect 16390 38808 16396 38820
rect 15396 38780 16396 38808
rect 16390 38768 16396 38780
rect 16448 38768 16454 38820
rect 5592 38712 8708 38740
rect 5592 38700 5598 38712
rect 8754 38700 8760 38752
rect 8812 38740 8818 38752
rect 8849 38743 8907 38749
rect 8849 38740 8861 38743
rect 8812 38712 8861 38740
rect 8812 38700 8818 38712
rect 8849 38709 8861 38712
rect 8895 38709 8907 38743
rect 8849 38703 8907 38709
rect 13814 38700 13820 38752
rect 13872 38740 13878 38752
rect 14001 38743 14059 38749
rect 14001 38740 14013 38743
rect 13872 38712 14013 38740
rect 13872 38700 13878 38712
rect 14001 38709 14013 38712
rect 14047 38709 14059 38743
rect 14001 38703 14059 38709
rect 16114 38700 16120 38752
rect 16172 38740 16178 38752
rect 16853 38743 16911 38749
rect 16853 38740 16865 38743
rect 16172 38712 16865 38740
rect 16172 38700 16178 38712
rect 16853 38709 16865 38712
rect 16899 38709 16911 38743
rect 16853 38703 16911 38709
rect 1104 38650 24840 38672
rect 1104 38598 8912 38650
rect 8964 38598 8976 38650
rect 9028 38598 9040 38650
rect 9092 38598 9104 38650
rect 9156 38598 16843 38650
rect 16895 38598 16907 38650
rect 16959 38598 16971 38650
rect 17023 38598 17035 38650
rect 17087 38598 24840 38650
rect 1104 38576 24840 38598
rect 3510 38496 3516 38548
rect 3568 38536 3574 38548
rect 4341 38539 4399 38545
rect 4341 38536 4353 38539
rect 3568 38508 4353 38536
rect 3568 38496 3574 38508
rect 4341 38505 4353 38508
rect 4387 38505 4399 38539
rect 4341 38499 4399 38505
rect 7742 38496 7748 38548
rect 7800 38536 7806 38548
rect 8665 38539 8723 38545
rect 8665 38536 8677 38539
rect 7800 38508 8677 38536
rect 7800 38496 7806 38508
rect 8665 38505 8677 38508
rect 8711 38505 8723 38539
rect 9858 38536 9864 38548
rect 9819 38508 9864 38536
rect 8665 38499 8723 38505
rect 9858 38496 9864 38508
rect 9916 38496 9922 38548
rect 1946 38428 1952 38480
rect 2004 38468 2010 38480
rect 2004 38440 3556 38468
rect 2004 38428 2010 38440
rect 2869 38403 2927 38409
rect 2869 38369 2881 38403
rect 2915 38369 2927 38403
rect 3528 38400 3556 38440
rect 3602 38428 3608 38480
rect 3660 38468 3666 38480
rect 3660 38440 4292 38468
rect 3660 38428 3666 38440
rect 4062 38400 4068 38412
rect 3528 38372 4068 38400
rect 2869 38363 2927 38369
rect 2884 38196 2912 38363
rect 4062 38360 4068 38372
rect 4120 38360 4126 38412
rect 4264 38409 4292 38440
rect 8754 38428 8760 38480
rect 8812 38468 8818 38480
rect 12621 38471 12679 38477
rect 8812 38440 11100 38468
rect 8812 38428 8818 38440
rect 4249 38403 4307 38409
rect 4249 38369 4261 38403
rect 4295 38369 4307 38403
rect 4249 38363 4307 38369
rect 5813 38403 5871 38409
rect 5813 38369 5825 38403
rect 5859 38400 5871 38403
rect 5994 38400 6000 38412
rect 5859 38372 6000 38400
rect 5859 38369 5871 38372
rect 5813 38363 5871 38369
rect 5994 38360 6000 38372
rect 6052 38360 6058 38412
rect 6089 38403 6147 38409
rect 6089 38369 6101 38403
rect 6135 38369 6147 38403
rect 6089 38363 6147 38369
rect 5902 38332 5908 38344
rect 3068 38304 5908 38332
rect 3068 38273 3096 38304
rect 5902 38292 5908 38304
rect 5960 38332 5966 38344
rect 6104 38332 6132 38363
rect 6638 38360 6644 38412
rect 6696 38400 6702 38412
rect 7101 38403 7159 38409
rect 7101 38400 7113 38403
rect 6696 38372 7113 38400
rect 6696 38360 6702 38372
rect 7101 38369 7113 38372
rect 7147 38369 7159 38403
rect 7101 38363 7159 38369
rect 7469 38403 7527 38409
rect 7469 38369 7481 38403
rect 7515 38400 7527 38403
rect 7558 38400 7564 38412
rect 7515 38372 7564 38400
rect 7515 38369 7527 38372
rect 7469 38363 7527 38369
rect 7558 38360 7564 38372
rect 7616 38360 7622 38412
rect 7650 38360 7656 38412
rect 7708 38400 7714 38412
rect 7708 38372 7801 38400
rect 7708 38360 7714 38372
rect 8662 38360 8668 38412
rect 8720 38400 8726 38412
rect 9692 38409 9720 38440
rect 8849 38403 8907 38409
rect 8849 38400 8861 38403
rect 8720 38372 8861 38400
rect 8720 38360 8726 38372
rect 8849 38369 8861 38372
rect 8895 38369 8907 38403
rect 8849 38363 8907 38369
rect 9677 38403 9735 38409
rect 9677 38369 9689 38403
rect 9723 38369 9735 38403
rect 9677 38363 9735 38369
rect 10870 38360 10876 38412
rect 10928 38400 10934 38412
rect 10965 38403 11023 38409
rect 10965 38400 10977 38403
rect 10928 38372 10977 38400
rect 10928 38360 10934 38372
rect 10965 38369 10977 38372
rect 11011 38369 11023 38403
rect 11072 38400 11100 38440
rect 12621 38437 12633 38471
rect 12667 38468 12679 38471
rect 13814 38468 13820 38480
rect 12667 38440 13820 38468
rect 12667 38437 12679 38440
rect 12621 38431 12679 38437
rect 13814 38428 13820 38440
rect 13872 38428 13878 38480
rect 15746 38468 15752 38480
rect 14016 38440 15752 38468
rect 11330 38400 11336 38412
rect 11072 38372 11336 38400
rect 10965 38363 11023 38369
rect 11330 38360 11336 38372
rect 11388 38360 11394 38412
rect 14016 38409 14044 38440
rect 15746 38428 15752 38440
rect 15804 38428 15810 38480
rect 16482 38428 16488 38480
rect 16540 38468 16546 38480
rect 16853 38471 16911 38477
rect 16853 38468 16865 38471
rect 16540 38440 16865 38468
rect 16540 38428 16546 38440
rect 16853 38437 16865 38440
rect 16899 38437 16911 38471
rect 16853 38431 16911 38437
rect 13909 38403 13967 38409
rect 13909 38369 13921 38403
rect 13955 38369 13967 38403
rect 13909 38363 13967 38369
rect 14001 38403 14059 38409
rect 14001 38369 14013 38403
rect 14047 38369 14059 38403
rect 14001 38363 14059 38369
rect 14369 38403 14427 38409
rect 14369 38369 14381 38403
rect 14415 38400 14427 38403
rect 14458 38400 14464 38412
rect 14415 38372 14464 38400
rect 14415 38369 14427 38372
rect 14369 38363 14427 38369
rect 7668 38332 7696 38360
rect 11238 38332 11244 38344
rect 5960 38304 7696 38332
rect 11199 38304 11244 38332
rect 5960 38292 5966 38304
rect 11238 38292 11244 38304
rect 11296 38292 11302 38344
rect 13924 38332 13952 38363
rect 14458 38360 14464 38372
rect 14516 38360 14522 38412
rect 15562 38400 15568 38412
rect 15523 38372 15568 38400
rect 15562 38360 15568 38372
rect 15620 38360 15626 38412
rect 15838 38400 15844 38412
rect 15799 38372 15844 38400
rect 15838 38360 15844 38372
rect 15896 38360 15902 38412
rect 17037 38403 17095 38409
rect 17037 38369 17049 38403
rect 17083 38400 17095 38403
rect 19978 38400 19984 38412
rect 17083 38372 19984 38400
rect 17083 38369 17095 38372
rect 17037 38363 17095 38369
rect 19978 38360 19984 38372
rect 20036 38360 20042 38412
rect 14550 38332 14556 38344
rect 13924 38304 14556 38332
rect 14550 38292 14556 38304
rect 14608 38292 14614 38344
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38332 15715 38335
rect 16298 38332 16304 38344
rect 15703 38304 16304 38332
rect 15703 38301 15715 38304
rect 15657 38295 15715 38301
rect 16298 38292 16304 38304
rect 16356 38292 16362 38344
rect 3053 38267 3111 38273
rect 3053 38233 3065 38267
rect 3099 38233 3111 38267
rect 3053 38227 3111 38233
rect 5442 38224 5448 38276
rect 5500 38264 5506 38276
rect 5629 38267 5687 38273
rect 5629 38264 5641 38267
rect 5500 38236 5641 38264
rect 5500 38224 5506 38236
rect 5629 38233 5641 38236
rect 5675 38233 5687 38267
rect 5629 38227 5687 38233
rect 8754 38196 8760 38208
rect 2884 38168 8760 38196
rect 8754 38156 8760 38168
rect 8812 38156 8818 38208
rect 10962 38156 10968 38208
rect 11020 38196 11026 38208
rect 13170 38196 13176 38208
rect 11020 38168 13176 38196
rect 11020 38156 11026 38168
rect 13170 38156 13176 38168
rect 13228 38156 13234 38208
rect 16206 38156 16212 38208
rect 16264 38196 16270 38208
rect 17129 38199 17187 38205
rect 17129 38196 17141 38199
rect 16264 38168 17141 38196
rect 16264 38156 16270 38168
rect 17129 38165 17141 38168
rect 17175 38165 17187 38199
rect 17129 38159 17187 38165
rect 1104 38106 24840 38128
rect 1104 38054 4947 38106
rect 4999 38054 5011 38106
rect 5063 38054 5075 38106
rect 5127 38054 5139 38106
rect 5191 38054 12878 38106
rect 12930 38054 12942 38106
rect 12994 38054 13006 38106
rect 13058 38054 13070 38106
rect 13122 38054 20808 38106
rect 20860 38054 20872 38106
rect 20924 38054 20936 38106
rect 20988 38054 21000 38106
rect 21052 38054 24840 38106
rect 1104 38032 24840 38054
rect 3418 37952 3424 38004
rect 3476 37992 3482 38004
rect 3973 37995 4031 38001
rect 3973 37992 3985 37995
rect 3476 37964 3985 37992
rect 3476 37952 3482 37964
rect 3973 37961 3985 37964
rect 4019 37961 4031 37995
rect 3973 37955 4031 37961
rect 5813 37995 5871 38001
rect 5813 37961 5825 37995
rect 5859 37992 5871 37995
rect 6362 37992 6368 38004
rect 5859 37964 6368 37992
rect 5859 37961 5871 37964
rect 5813 37955 5871 37961
rect 6362 37952 6368 37964
rect 6420 37952 6426 38004
rect 6730 37952 6736 38004
rect 6788 37992 6794 38004
rect 6917 37995 6975 38001
rect 6917 37992 6929 37995
rect 6788 37964 6929 37992
rect 6788 37952 6794 37964
rect 6917 37961 6929 37964
rect 6963 37961 6975 37995
rect 10962 37992 10968 38004
rect 6917 37955 6975 37961
rect 7024 37964 9444 37992
rect 10923 37964 10968 37992
rect 6270 37884 6276 37936
rect 6328 37924 6334 37936
rect 7024 37924 7052 37964
rect 6328 37896 7052 37924
rect 9416 37924 9444 37964
rect 10962 37952 10968 37964
rect 11020 37952 11026 38004
rect 11422 37992 11428 38004
rect 11383 37964 11428 37992
rect 11422 37952 11428 37964
rect 11480 37952 11486 38004
rect 12710 37952 12716 38004
rect 12768 37992 12774 38004
rect 12989 37995 13047 38001
rect 12989 37992 13001 37995
rect 12768 37964 13001 37992
rect 12768 37952 12774 37964
rect 12989 37961 13001 37964
rect 13035 37961 13047 37995
rect 12989 37955 13047 37961
rect 12250 37924 12256 37936
rect 9416 37896 12256 37924
rect 6328 37884 6334 37896
rect 12250 37884 12256 37896
rect 12308 37884 12314 37936
rect 7834 37816 7840 37868
rect 7892 37856 7898 37868
rect 8481 37859 8539 37865
rect 8481 37856 8493 37859
rect 7892 37828 8493 37856
rect 7892 37816 7898 37828
rect 8481 37825 8493 37828
rect 8527 37825 8539 37859
rect 8481 37819 8539 37825
rect 10870 37816 10876 37868
rect 10928 37856 10934 37868
rect 12066 37856 12072 37868
rect 10928 37828 12072 37856
rect 10928 37816 10934 37828
rect 12066 37816 12072 37828
rect 12124 37816 12130 37868
rect 13446 37856 13452 37868
rect 13407 37828 13452 37856
rect 13446 37816 13452 37828
rect 13504 37816 13510 37868
rect 18141 37859 18199 37865
rect 18141 37856 18153 37859
rect 13556 37828 18153 37856
rect 2869 37791 2927 37797
rect 2869 37757 2881 37791
rect 2915 37757 2927 37791
rect 3878 37788 3884 37800
rect 3839 37760 3884 37788
rect 2869 37751 2927 37757
rect 2884 37652 2912 37751
rect 3878 37748 3884 37760
rect 3936 37748 3942 37800
rect 4522 37788 4528 37800
rect 4483 37760 4528 37788
rect 4522 37748 4528 37760
rect 4580 37748 4586 37800
rect 5534 37748 5540 37800
rect 5592 37788 5598 37800
rect 5629 37791 5687 37797
rect 5629 37788 5641 37791
rect 5592 37760 5641 37788
rect 5592 37748 5598 37760
rect 5629 37757 5641 37760
rect 5675 37757 5687 37791
rect 5629 37751 5687 37757
rect 6362 37748 6368 37800
rect 6420 37788 6426 37800
rect 6825 37791 6883 37797
rect 6825 37788 6837 37791
rect 6420 37760 6837 37788
rect 6420 37748 6426 37760
rect 6825 37757 6837 37760
rect 6871 37757 6883 37791
rect 6825 37751 6883 37757
rect 7561 37791 7619 37797
rect 7561 37757 7573 37791
rect 7607 37788 7619 37791
rect 7650 37788 7656 37800
rect 7607 37760 7656 37788
rect 7607 37757 7619 37760
rect 7561 37751 7619 37757
rect 7650 37748 7656 37760
rect 7708 37748 7714 37800
rect 8754 37788 8760 37800
rect 8715 37760 8760 37788
rect 8754 37748 8760 37760
rect 8812 37748 8818 37800
rect 11149 37791 11207 37797
rect 11149 37757 11161 37791
rect 11195 37757 11207 37791
rect 11149 37751 11207 37757
rect 11241 37791 11299 37797
rect 11241 37757 11253 37791
rect 11287 37788 11299 37791
rect 11330 37788 11336 37800
rect 11287 37760 11336 37788
rect 11287 37757 11299 37760
rect 11241 37751 11299 37757
rect 2961 37723 3019 37729
rect 2961 37689 2973 37723
rect 3007 37720 3019 37723
rect 8018 37720 8024 37732
rect 3007 37692 8024 37720
rect 3007 37689 3019 37692
rect 2961 37683 3019 37689
rect 8018 37680 8024 37692
rect 8076 37680 8082 37732
rect 11164 37720 11192 37751
rect 11330 37748 11336 37760
rect 11388 37788 11394 37800
rect 13556 37797 13584 37828
rect 18141 37825 18153 37828
rect 18187 37825 18199 37859
rect 18141 37819 18199 37825
rect 13541 37791 13599 37797
rect 11388 37760 13492 37788
rect 11388 37748 11394 37760
rect 11606 37720 11612 37732
rect 11164 37692 11612 37720
rect 11606 37680 11612 37692
rect 11664 37680 11670 37732
rect 13464 37720 13492 37760
rect 13541 37757 13553 37791
rect 13587 37757 13599 37791
rect 13541 37751 13599 37757
rect 13814 37748 13820 37800
rect 13872 37788 13878 37800
rect 13909 37791 13967 37797
rect 13909 37788 13921 37791
rect 13872 37760 13921 37788
rect 13872 37748 13878 37760
rect 13909 37757 13921 37760
rect 13955 37757 13967 37791
rect 14090 37788 14096 37800
rect 14051 37760 14096 37788
rect 13909 37751 13967 37757
rect 14090 37748 14096 37760
rect 14148 37748 14154 37800
rect 14921 37791 14979 37797
rect 14921 37757 14933 37791
rect 14967 37757 14979 37791
rect 14921 37751 14979 37757
rect 14936 37720 14964 37751
rect 15102 37748 15108 37800
rect 15160 37788 15166 37800
rect 16022 37788 16028 37800
rect 15160 37760 15884 37788
rect 15983 37760 16028 37788
rect 15160 37748 15166 37760
rect 15286 37720 15292 37732
rect 13464 37692 15292 37720
rect 15286 37680 15292 37692
rect 15344 37680 15350 37732
rect 10042 37652 10048 37664
rect 2884 37624 10048 37652
rect 10042 37612 10048 37624
rect 10100 37612 10106 37664
rect 11514 37612 11520 37664
rect 11572 37652 11578 37664
rect 13170 37652 13176 37664
rect 11572 37624 13176 37652
rect 11572 37612 11578 37624
rect 13170 37612 13176 37624
rect 13228 37612 13234 37664
rect 15105 37655 15163 37661
rect 15105 37621 15117 37655
rect 15151 37652 15163 37655
rect 15746 37652 15752 37664
rect 15151 37624 15752 37652
rect 15151 37621 15163 37624
rect 15105 37615 15163 37621
rect 15746 37612 15752 37624
rect 15804 37612 15810 37664
rect 15856 37652 15884 37760
rect 16022 37748 16028 37760
rect 16080 37748 16086 37800
rect 16298 37788 16304 37800
rect 16259 37760 16304 37788
rect 16298 37748 16304 37760
rect 16356 37748 16362 37800
rect 18049 37791 18107 37797
rect 18049 37757 18061 37791
rect 18095 37757 18107 37791
rect 18049 37751 18107 37757
rect 16206 37720 16212 37732
rect 16167 37692 16212 37720
rect 16206 37680 16212 37692
rect 16264 37680 16270 37732
rect 16666 37680 16672 37732
rect 16724 37720 16730 37732
rect 16761 37723 16819 37729
rect 16761 37720 16773 37723
rect 16724 37692 16773 37720
rect 16724 37680 16730 37692
rect 16761 37689 16773 37692
rect 16807 37689 16819 37723
rect 16761 37683 16819 37689
rect 18064 37652 18092 37751
rect 15856 37624 18092 37652
rect 1104 37562 24840 37584
rect 1104 37510 8912 37562
rect 8964 37510 8976 37562
rect 9028 37510 9040 37562
rect 9092 37510 9104 37562
rect 9156 37510 16843 37562
rect 16895 37510 16907 37562
rect 16959 37510 16971 37562
rect 17023 37510 17035 37562
rect 17087 37510 24840 37562
rect 1104 37488 24840 37510
rect 5626 37448 5632 37460
rect 2608 37420 5632 37448
rect 2608 37389 2636 37420
rect 5626 37408 5632 37420
rect 5684 37408 5690 37460
rect 5718 37408 5724 37460
rect 5776 37448 5782 37460
rect 6089 37451 6147 37457
rect 6089 37448 6101 37451
rect 5776 37420 6101 37448
rect 5776 37408 5782 37420
rect 6089 37417 6101 37420
rect 6135 37417 6147 37451
rect 6089 37411 6147 37417
rect 8018 37408 8024 37460
rect 8076 37448 8082 37460
rect 12066 37448 12072 37460
rect 8076 37420 11652 37448
rect 12027 37420 12072 37448
rect 8076 37408 8082 37420
rect 2593 37383 2651 37389
rect 2593 37349 2605 37383
rect 2639 37349 2651 37383
rect 8665 37383 8723 37389
rect 2593 37343 2651 37349
rect 7576 37352 8156 37380
rect 7576 37324 7604 37352
rect 2406 37312 2412 37324
rect 2367 37284 2412 37312
rect 2406 37272 2412 37284
rect 2464 37272 2470 37324
rect 2685 37315 2743 37321
rect 2685 37281 2697 37315
rect 2731 37312 2743 37315
rect 4154 37312 4160 37324
rect 2731 37284 4160 37312
rect 2731 37281 2743 37284
rect 2685 37275 2743 37281
rect 4154 37272 4160 37284
rect 4212 37272 4218 37324
rect 4709 37315 4767 37321
rect 4709 37281 4721 37315
rect 4755 37281 4767 37315
rect 4709 37275 4767 37281
rect 4985 37315 5043 37321
rect 4985 37281 4997 37315
rect 5031 37312 5043 37315
rect 7098 37312 7104 37324
rect 5031 37284 7104 37312
rect 5031 37281 5043 37284
rect 4985 37275 5043 37281
rect 4246 37204 4252 37256
rect 4304 37244 4310 37256
rect 4724 37244 4752 37275
rect 7098 37272 7104 37284
rect 7156 37272 7162 37324
rect 7558 37312 7564 37324
rect 7519 37284 7564 37312
rect 7558 37272 7564 37284
rect 7616 37272 7622 37324
rect 7653 37315 7711 37321
rect 7653 37281 7665 37315
rect 7699 37312 7711 37315
rect 8018 37312 8024 37324
rect 7699 37284 7788 37312
rect 7979 37284 8024 37312
rect 7699 37281 7711 37284
rect 7653 37275 7711 37281
rect 5442 37244 5448 37256
rect 4304 37216 5448 37244
rect 4304 37204 4310 37216
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 7760 37176 7788 37284
rect 8018 37272 8024 37284
rect 8076 37272 8082 37324
rect 8128 37321 8156 37352
rect 8665 37349 8677 37383
rect 8711 37380 8723 37383
rect 8754 37380 8760 37392
rect 8711 37352 8760 37380
rect 8711 37349 8723 37352
rect 8665 37343 8723 37349
rect 8754 37340 8760 37352
rect 8812 37340 8818 37392
rect 10410 37380 10416 37392
rect 9784 37352 10416 37380
rect 9784 37321 9812 37352
rect 10410 37340 10416 37352
rect 10468 37340 10474 37392
rect 11057 37383 11115 37389
rect 11057 37349 11069 37383
rect 11103 37380 11115 37383
rect 11238 37380 11244 37392
rect 11103 37352 11244 37380
rect 11103 37349 11115 37352
rect 11057 37343 11115 37349
rect 11238 37340 11244 37352
rect 11296 37340 11302 37392
rect 8113 37315 8171 37321
rect 8113 37281 8125 37315
rect 8159 37281 8171 37315
rect 9769 37315 9827 37321
rect 9769 37312 9781 37315
rect 8113 37275 8171 37281
rect 8496 37284 9781 37312
rect 8496 37176 8524 37284
rect 9769 37281 9781 37284
rect 9815 37281 9827 37315
rect 9769 37275 9827 37281
rect 9953 37315 10011 37321
rect 9953 37281 9965 37315
rect 9999 37312 10011 37315
rect 10318 37312 10324 37324
rect 9999 37284 10324 37312
rect 9999 37281 10011 37284
rect 9953 37275 10011 37281
rect 10318 37272 10324 37284
rect 10376 37312 10382 37324
rect 10505 37315 10563 37321
rect 10505 37312 10517 37315
rect 10376 37284 10517 37312
rect 10376 37272 10382 37284
rect 10505 37281 10517 37284
rect 10551 37281 10563 37315
rect 10505 37275 10563 37281
rect 10689 37315 10747 37321
rect 10689 37281 10701 37315
rect 10735 37312 10747 37315
rect 11514 37312 11520 37324
rect 10735 37284 11520 37312
rect 10735 37281 10747 37284
rect 10689 37275 10747 37281
rect 11514 37272 11520 37284
rect 11572 37272 11578 37324
rect 11624 37312 11652 37420
rect 12066 37408 12072 37420
rect 12124 37408 12130 37460
rect 14458 37408 14464 37460
rect 14516 37448 14522 37460
rect 15473 37451 15531 37457
rect 15473 37448 15485 37451
rect 14516 37420 15485 37448
rect 14516 37408 14522 37420
rect 15473 37417 15485 37420
rect 15519 37417 15531 37451
rect 15473 37411 15531 37417
rect 11698 37340 11704 37392
rect 11756 37380 11762 37392
rect 14093 37383 14151 37389
rect 14093 37380 14105 37383
rect 11756 37352 13032 37380
rect 11756 37340 11762 37352
rect 13004 37321 13032 37352
rect 13188 37352 14105 37380
rect 13188 37324 13216 37352
rect 14093 37349 14105 37352
rect 14139 37349 14151 37383
rect 14093 37343 14151 37349
rect 14918 37340 14924 37392
rect 14976 37380 14982 37392
rect 18141 37383 18199 37389
rect 14976 37352 16528 37380
rect 14976 37340 14982 37352
rect 12437 37315 12495 37321
rect 12437 37312 12449 37315
rect 11624 37284 12449 37312
rect 12437 37281 12449 37284
rect 12483 37281 12495 37315
rect 12621 37315 12679 37321
rect 12621 37312 12633 37315
rect 12437 37275 12495 37281
rect 12544 37284 12633 37312
rect 11238 37204 11244 37256
rect 11296 37244 11302 37256
rect 12544 37244 12572 37284
rect 12621 37281 12633 37284
rect 12667 37281 12679 37315
rect 12621 37275 12679 37281
rect 12989 37315 13047 37321
rect 12989 37281 13001 37315
rect 13035 37281 13047 37315
rect 13170 37312 13176 37324
rect 13131 37284 13176 37312
rect 12989 37275 13047 37281
rect 13170 37272 13176 37284
rect 13228 37272 13234 37324
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 14001 37315 14059 37321
rect 14001 37312 14013 37315
rect 13872 37284 14013 37312
rect 13872 37272 13878 37284
rect 14001 37281 14013 37284
rect 14047 37281 14059 37315
rect 15286 37312 15292 37324
rect 15247 37284 15292 37312
rect 14001 37275 14059 37281
rect 15286 37272 15292 37284
rect 15344 37272 15350 37324
rect 16500 37321 16528 37352
rect 18141 37349 18153 37383
rect 18187 37380 18199 37383
rect 19978 37380 19984 37392
rect 18187 37352 19984 37380
rect 18187 37349 18199 37352
rect 18141 37343 18199 37349
rect 19978 37340 19984 37352
rect 20036 37340 20042 37392
rect 16485 37315 16543 37321
rect 16485 37281 16497 37315
rect 16531 37281 16543 37315
rect 16758 37312 16764 37324
rect 16719 37284 16764 37312
rect 16485 37275 16543 37281
rect 16758 37272 16764 37284
rect 16816 37272 16822 37324
rect 11296 37216 12572 37244
rect 11296 37204 11302 37216
rect 7760 37148 8524 37176
rect 2869 37111 2927 37117
rect 2869 37077 2881 37111
rect 2915 37108 2927 37111
rect 3050 37108 3056 37120
rect 2915 37080 3056 37108
rect 2915 37077 2927 37080
rect 2869 37071 2927 37077
rect 3050 37068 3056 37080
rect 3108 37068 3114 37120
rect 8110 37068 8116 37120
rect 8168 37108 8174 37120
rect 16022 37108 16028 37120
rect 8168 37080 16028 37108
rect 8168 37068 8174 37080
rect 16022 37068 16028 37080
rect 16080 37068 16086 37120
rect 1104 37018 24840 37040
rect 1104 36966 4947 37018
rect 4999 36966 5011 37018
rect 5063 36966 5075 37018
rect 5127 36966 5139 37018
rect 5191 36966 12878 37018
rect 12930 36966 12942 37018
rect 12994 36966 13006 37018
rect 13058 36966 13070 37018
rect 13122 36966 20808 37018
rect 20860 36966 20872 37018
rect 20924 36966 20936 37018
rect 20988 36966 21000 37018
rect 21052 36966 24840 37018
rect 1104 36944 24840 36966
rect 4338 36904 4344 36916
rect 4299 36876 4344 36904
rect 4338 36864 4344 36876
rect 4396 36864 4402 36916
rect 5537 36907 5595 36913
rect 5537 36873 5549 36907
rect 5583 36904 5595 36907
rect 5626 36904 5632 36916
rect 5583 36876 5632 36904
rect 5583 36873 5595 36876
rect 5537 36867 5595 36873
rect 5626 36864 5632 36876
rect 5684 36864 5690 36916
rect 7098 36904 7104 36916
rect 7059 36876 7104 36904
rect 7098 36864 7104 36876
rect 7156 36864 7162 36916
rect 8110 36864 8116 36916
rect 8168 36904 8174 36916
rect 8389 36907 8447 36913
rect 8389 36904 8401 36907
rect 8168 36876 8401 36904
rect 8168 36864 8174 36876
rect 8389 36873 8401 36876
rect 8435 36873 8447 36907
rect 10778 36904 10784 36916
rect 10739 36876 10784 36904
rect 8389 36867 8447 36873
rect 10778 36864 10784 36876
rect 10836 36864 10842 36916
rect 10962 36864 10968 36916
rect 11020 36904 11026 36916
rect 12897 36907 12955 36913
rect 12897 36904 12909 36907
rect 11020 36876 12909 36904
rect 11020 36864 11026 36876
rect 12897 36873 12909 36876
rect 12943 36904 12955 36907
rect 15194 36904 15200 36916
rect 12943 36876 15200 36904
rect 12943 36873 12955 36876
rect 12897 36867 12955 36873
rect 15194 36864 15200 36876
rect 15252 36904 15258 36916
rect 15930 36904 15936 36916
rect 15252 36876 15936 36904
rect 15252 36864 15258 36876
rect 15930 36864 15936 36876
rect 15988 36864 15994 36916
rect 16117 36907 16175 36913
rect 16117 36873 16129 36907
rect 16163 36904 16175 36907
rect 16298 36904 16304 36916
rect 16163 36876 16304 36904
rect 16163 36873 16175 36876
rect 16117 36867 16175 36873
rect 16298 36864 16304 36876
rect 16356 36864 16362 36916
rect 3050 36768 3056 36780
rect 3011 36740 3056 36768
rect 3050 36728 3056 36740
rect 3108 36728 3114 36780
rect 4246 36768 4252 36780
rect 3988 36740 4252 36768
rect 2777 36703 2835 36709
rect 2777 36669 2789 36703
rect 2823 36700 2835 36703
rect 3988 36700 4016 36740
rect 4246 36728 4252 36740
rect 4304 36728 4310 36780
rect 4356 36768 4384 36864
rect 6825 36771 6883 36777
rect 4356 36740 5488 36768
rect 2823 36672 4016 36700
rect 2823 36669 2835 36672
rect 2777 36663 2835 36669
rect 4062 36660 4068 36712
rect 4120 36700 4126 36712
rect 5261 36703 5319 36709
rect 5261 36700 5273 36703
rect 4120 36672 5273 36700
rect 4120 36660 4126 36672
rect 5261 36669 5273 36672
rect 5307 36700 5319 36703
rect 5350 36700 5356 36712
rect 5307 36672 5356 36700
rect 5307 36669 5319 36672
rect 5261 36663 5319 36669
rect 5350 36660 5356 36672
rect 5408 36660 5414 36712
rect 5460 36709 5488 36740
rect 6825 36737 6837 36771
rect 6871 36768 6883 36771
rect 8128 36768 8156 36864
rect 9674 36768 9680 36780
rect 6871 36740 8156 36768
rect 9635 36740 9680 36768
rect 6871 36737 6883 36740
rect 6825 36731 6883 36737
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 12434 36768 12440 36780
rect 11992 36740 12440 36768
rect 5445 36703 5503 36709
rect 5445 36669 5457 36703
rect 5491 36669 5503 36703
rect 5445 36663 5503 36669
rect 6914 36660 6920 36712
rect 6972 36700 6978 36712
rect 6972 36672 7017 36700
rect 6972 36660 6978 36672
rect 7926 36660 7932 36712
rect 7984 36700 7990 36712
rect 8205 36703 8263 36709
rect 8205 36700 8217 36703
rect 7984 36672 8217 36700
rect 7984 36660 7990 36672
rect 8205 36669 8217 36672
rect 8251 36669 8263 36703
rect 8205 36663 8263 36669
rect 9493 36703 9551 36709
rect 9493 36669 9505 36703
rect 9539 36669 9551 36703
rect 9766 36700 9772 36712
rect 9727 36672 9772 36700
rect 9493 36663 9551 36669
rect 9508 36632 9536 36663
rect 9766 36660 9772 36672
rect 9824 36660 9830 36712
rect 10318 36660 10324 36712
rect 10376 36700 10382 36712
rect 10505 36703 10563 36709
rect 10376 36672 10421 36700
rect 10376 36660 10382 36672
rect 10505 36669 10517 36703
rect 10551 36700 10563 36703
rect 11330 36700 11336 36712
rect 10551 36672 11336 36700
rect 10551 36669 10563 36672
rect 10505 36663 10563 36669
rect 11330 36660 11336 36672
rect 11388 36660 11394 36712
rect 11992 36709 12020 36740
rect 12434 36728 12440 36740
rect 12492 36728 12498 36780
rect 14458 36728 14464 36780
rect 14516 36768 14522 36780
rect 15102 36768 15108 36780
rect 14516 36740 15108 36768
rect 14516 36728 14522 36740
rect 15102 36728 15108 36740
rect 15160 36728 15166 36780
rect 11977 36703 12035 36709
rect 11977 36669 11989 36703
rect 12023 36669 12035 36703
rect 11977 36663 12035 36669
rect 12805 36703 12863 36709
rect 12805 36669 12817 36703
rect 12851 36700 12863 36703
rect 13354 36700 13360 36712
rect 12851 36672 13360 36700
rect 12851 36669 12863 36672
rect 12805 36663 12863 36669
rect 11992 36632 12020 36663
rect 13354 36660 13360 36672
rect 13412 36660 13418 36712
rect 14642 36700 14648 36712
rect 14603 36672 14648 36700
rect 14642 36660 14648 36672
rect 14700 36660 14706 36712
rect 14734 36660 14740 36712
rect 14792 36700 14798 36712
rect 15010 36700 15016 36712
rect 14792 36672 14837 36700
rect 14971 36672 15016 36700
rect 14792 36660 14798 36672
rect 15010 36660 15016 36672
rect 15068 36660 15074 36712
rect 15470 36660 15476 36712
rect 15528 36700 15534 36712
rect 16025 36703 16083 36709
rect 16025 36700 16037 36703
rect 15528 36672 16037 36700
rect 15528 36660 15534 36672
rect 16025 36669 16037 36672
rect 16071 36669 16083 36703
rect 16025 36663 16083 36669
rect 16577 36703 16635 36709
rect 16577 36669 16589 36703
rect 16623 36669 16635 36703
rect 16577 36663 16635 36669
rect 9508 36604 12020 36632
rect 12621 36635 12679 36641
rect 12621 36601 12633 36635
rect 12667 36632 12679 36635
rect 13630 36632 13636 36644
rect 12667 36604 13636 36632
rect 12667 36601 12679 36604
rect 12621 36595 12679 36601
rect 13630 36592 13636 36604
rect 13688 36592 13694 36644
rect 14001 36635 14059 36641
rect 14001 36601 14013 36635
rect 14047 36632 14059 36635
rect 15102 36632 15108 36644
rect 14047 36604 15108 36632
rect 14047 36601 14059 36604
rect 14001 36595 14059 36601
rect 15102 36592 15108 36604
rect 15160 36592 15166 36644
rect 15746 36592 15752 36644
rect 15804 36632 15810 36644
rect 16592 36632 16620 36663
rect 15804 36604 16620 36632
rect 15804 36592 15810 36604
rect 3142 36524 3148 36576
rect 3200 36564 3206 36576
rect 5534 36564 5540 36576
rect 3200 36536 5540 36564
rect 3200 36524 3206 36536
rect 5534 36524 5540 36536
rect 5592 36524 5598 36576
rect 8754 36524 8760 36576
rect 8812 36564 8818 36576
rect 9309 36567 9367 36573
rect 9309 36564 9321 36567
rect 8812 36536 9321 36564
rect 8812 36524 8818 36536
rect 9309 36533 9321 36536
rect 9355 36533 9367 36567
rect 9309 36527 9367 36533
rect 9766 36524 9772 36576
rect 9824 36564 9830 36576
rect 10318 36564 10324 36576
rect 9824 36536 10324 36564
rect 9824 36524 9830 36536
rect 10318 36524 10324 36536
rect 10376 36524 10382 36576
rect 11606 36524 11612 36576
rect 11664 36564 11670 36576
rect 11793 36567 11851 36573
rect 11793 36564 11805 36567
rect 11664 36536 11805 36564
rect 11664 36524 11670 36536
rect 11793 36533 11805 36536
rect 11839 36564 11851 36567
rect 13538 36564 13544 36576
rect 11839 36536 13544 36564
rect 11839 36533 11851 36536
rect 11793 36527 11851 36533
rect 13538 36524 13544 36536
rect 13596 36524 13602 36576
rect 1104 36474 24840 36496
rect 1104 36422 8912 36474
rect 8964 36422 8976 36474
rect 9028 36422 9040 36474
rect 9092 36422 9104 36474
rect 9156 36422 16843 36474
rect 16895 36422 16907 36474
rect 16959 36422 16971 36474
rect 17023 36422 17035 36474
rect 17087 36422 24840 36474
rect 1104 36400 24840 36422
rect 6454 36360 6460 36372
rect 2976 36332 6460 36360
rect 2976 36233 3004 36332
rect 6454 36320 6460 36332
rect 6512 36320 6518 36372
rect 10597 36363 10655 36369
rect 10597 36329 10609 36363
rect 10643 36360 10655 36363
rect 10686 36360 10692 36372
rect 10643 36332 10692 36360
rect 10643 36329 10655 36332
rect 10597 36323 10655 36329
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 15378 36320 15384 36372
rect 15436 36360 15442 36372
rect 15749 36363 15807 36369
rect 15749 36360 15761 36363
rect 15436 36332 15761 36360
rect 15436 36320 15442 36332
rect 15749 36329 15761 36332
rect 15795 36329 15807 36363
rect 15749 36323 15807 36329
rect 3053 36295 3111 36301
rect 3053 36261 3065 36295
rect 3099 36292 3111 36295
rect 3142 36292 3148 36304
rect 3099 36264 3148 36292
rect 3099 36261 3111 36264
rect 3053 36255 3111 36261
rect 3142 36252 3148 36264
rect 3200 36252 3206 36304
rect 4617 36295 4675 36301
rect 4617 36261 4629 36295
rect 4663 36292 4675 36295
rect 6914 36292 6920 36304
rect 4663 36264 6920 36292
rect 4663 36261 4675 36264
rect 4617 36255 4675 36261
rect 6914 36252 6920 36264
rect 6972 36252 6978 36304
rect 11238 36292 11244 36304
rect 10980 36264 11244 36292
rect 2961 36227 3019 36233
rect 2961 36193 2973 36227
rect 3007 36193 3019 36227
rect 5166 36224 5172 36236
rect 5127 36196 5172 36224
rect 2961 36187 3019 36193
rect 5166 36184 5172 36196
rect 5224 36184 5230 36236
rect 5261 36227 5319 36233
rect 5261 36193 5273 36227
rect 5307 36193 5319 36227
rect 5261 36187 5319 36193
rect 3234 35980 3240 36032
rect 3292 36020 3298 36032
rect 5276 36020 5304 36187
rect 5350 36184 5356 36236
rect 5408 36224 5414 36236
rect 5445 36227 5503 36233
rect 5445 36224 5457 36227
rect 5408 36196 5457 36224
rect 5408 36184 5414 36196
rect 5445 36193 5457 36196
rect 5491 36193 5503 36227
rect 5718 36224 5724 36236
rect 5679 36196 5724 36224
rect 5445 36187 5503 36193
rect 5718 36184 5724 36196
rect 5776 36184 5782 36236
rect 6089 36227 6147 36233
rect 6089 36193 6101 36227
rect 6135 36224 6147 36227
rect 6454 36224 6460 36236
rect 6135 36196 6460 36224
rect 6135 36193 6147 36196
rect 6089 36187 6147 36193
rect 6454 36184 6460 36196
rect 6512 36184 6518 36236
rect 10980 36233 11008 36264
rect 11238 36252 11244 36264
rect 11296 36252 11302 36304
rect 11514 36292 11520 36304
rect 11348 36264 11520 36292
rect 11348 36233 11376 36264
rect 11514 36252 11520 36264
rect 11572 36252 11578 36304
rect 13814 36252 13820 36304
rect 13872 36292 13878 36304
rect 15764 36292 15792 36323
rect 13872 36264 15608 36292
rect 15764 36264 17080 36292
rect 13872 36252 13878 36264
rect 10965 36227 11023 36233
rect 10965 36193 10977 36227
rect 11011 36193 11023 36227
rect 10965 36187 11023 36193
rect 11333 36227 11391 36233
rect 11333 36193 11345 36227
rect 11379 36193 11391 36227
rect 11333 36187 11391 36193
rect 11422 36184 11428 36236
rect 11480 36224 11486 36236
rect 12989 36227 13047 36233
rect 12989 36224 13001 36227
rect 11480 36196 13001 36224
rect 11480 36184 11486 36196
rect 12989 36193 13001 36196
rect 13035 36193 13047 36227
rect 13354 36224 13360 36236
rect 13315 36196 13360 36224
rect 12989 36187 13047 36193
rect 13354 36184 13360 36196
rect 13412 36184 13418 36236
rect 13541 36227 13599 36233
rect 13541 36193 13553 36227
rect 13587 36224 13599 36227
rect 13630 36224 13636 36236
rect 13587 36196 13636 36224
rect 13587 36193 13599 36196
rect 13541 36187 13599 36193
rect 13630 36184 13636 36196
rect 13688 36184 13694 36236
rect 14090 36184 14096 36236
rect 14148 36224 14154 36236
rect 15010 36224 15016 36236
rect 14148 36196 15016 36224
rect 14148 36184 14154 36196
rect 15010 36184 15016 36196
rect 15068 36224 15074 36236
rect 15580 36233 15608 36264
rect 15289 36227 15347 36233
rect 15289 36224 15301 36227
rect 15068 36196 15301 36224
rect 15068 36184 15074 36196
rect 15289 36193 15301 36196
rect 15335 36193 15347 36227
rect 15289 36187 15347 36193
rect 15565 36227 15623 36233
rect 15565 36193 15577 36227
rect 15611 36193 15623 36227
rect 15565 36187 15623 36193
rect 15930 36184 15936 36236
rect 15988 36224 15994 36236
rect 17052 36233 17080 36264
rect 16853 36227 16911 36233
rect 16853 36224 16865 36227
rect 15988 36196 16865 36224
rect 15988 36184 15994 36196
rect 16853 36193 16865 36196
rect 16899 36193 16911 36227
rect 16853 36187 16911 36193
rect 17037 36227 17095 36233
rect 17037 36193 17049 36227
rect 17083 36193 17095 36227
rect 17037 36187 17095 36193
rect 5534 36116 5540 36168
rect 5592 36156 5598 36168
rect 7101 36159 7159 36165
rect 7101 36156 7113 36159
rect 5592 36128 7113 36156
rect 5592 36116 5598 36128
rect 7101 36125 7113 36128
rect 7147 36125 7159 36159
rect 7374 36156 7380 36168
rect 7335 36128 7380 36156
rect 7101 36119 7159 36125
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 8662 36116 8668 36168
rect 8720 36156 8726 36168
rect 10781 36159 10839 36165
rect 10781 36156 10793 36159
rect 8720 36128 10793 36156
rect 8720 36116 8726 36128
rect 10781 36125 10793 36128
rect 10827 36125 10839 36159
rect 10781 36119 10839 36125
rect 11241 36159 11299 36165
rect 11241 36125 11253 36159
rect 11287 36156 11299 36159
rect 13081 36159 13139 36165
rect 11287 36128 11376 36156
rect 11287 36125 11299 36128
rect 11241 36119 11299 36125
rect 11348 36100 11376 36128
rect 13081 36125 13093 36159
rect 13127 36156 13139 36159
rect 13446 36156 13452 36168
rect 13127 36128 13452 36156
rect 13127 36125 13139 36128
rect 13081 36119 13139 36125
rect 13446 36116 13452 36128
rect 13504 36156 13510 36168
rect 14734 36156 14740 36168
rect 13504 36128 14740 36156
rect 13504 36116 13510 36128
rect 14734 36116 14740 36128
rect 14792 36116 14798 36168
rect 11330 36048 11336 36100
rect 11388 36048 11394 36100
rect 15286 36048 15292 36100
rect 15344 36088 15350 36100
rect 15381 36091 15439 36097
rect 15381 36088 15393 36091
rect 15344 36060 15393 36088
rect 15344 36048 15350 36060
rect 15381 36057 15393 36060
rect 15427 36057 15439 36091
rect 15381 36051 15439 36057
rect 3292 35992 5304 36020
rect 8665 36023 8723 36029
rect 3292 35980 3298 35992
rect 8665 35989 8677 36023
rect 8711 36020 8723 36023
rect 8846 36020 8852 36032
rect 8711 35992 8852 36020
rect 8711 35989 8723 35992
rect 8665 35983 8723 35989
rect 8846 35980 8852 35992
rect 8904 35980 8910 36032
rect 12437 36023 12495 36029
rect 12437 35989 12449 36023
rect 12483 36020 12495 36023
rect 12710 36020 12716 36032
rect 12483 35992 12716 36020
rect 12483 35989 12495 35992
rect 12437 35983 12495 35989
rect 12710 35980 12716 35992
rect 12768 35980 12774 36032
rect 17126 36020 17132 36032
rect 17087 35992 17132 36020
rect 17126 35980 17132 35992
rect 17184 35980 17190 36032
rect 1104 35930 24840 35952
rect 1104 35878 4947 35930
rect 4999 35878 5011 35930
rect 5063 35878 5075 35930
rect 5127 35878 5139 35930
rect 5191 35878 12878 35930
rect 12930 35878 12942 35930
rect 12994 35878 13006 35930
rect 13058 35878 13070 35930
rect 13122 35878 20808 35930
rect 20860 35878 20872 35930
rect 20924 35878 20936 35930
rect 20988 35878 21000 35930
rect 21052 35878 24840 35930
rect 1104 35856 24840 35878
rect 8846 35816 8852 35828
rect 3528 35788 8852 35816
rect 2038 35640 2044 35692
rect 2096 35680 2102 35692
rect 2682 35680 2688 35692
rect 2096 35652 2688 35680
rect 2096 35640 2102 35652
rect 2682 35640 2688 35652
rect 2740 35640 2746 35692
rect 3528 35621 3556 35788
rect 8846 35776 8852 35788
rect 8904 35776 8910 35828
rect 10413 35819 10471 35825
rect 10413 35785 10425 35819
rect 10459 35816 10471 35819
rect 11422 35816 11428 35828
rect 10459 35788 11428 35816
rect 10459 35785 10471 35788
rect 10413 35779 10471 35785
rect 11422 35776 11428 35788
rect 11480 35776 11486 35828
rect 11698 35776 11704 35828
rect 11756 35816 11762 35828
rect 11756 35788 14780 35816
rect 11756 35776 11762 35788
rect 3605 35751 3663 35757
rect 3605 35717 3617 35751
rect 3651 35748 3663 35751
rect 3651 35720 7328 35748
rect 3651 35717 3663 35720
rect 3605 35711 3663 35717
rect 7300 35680 7328 35720
rect 7374 35708 7380 35760
rect 7432 35748 7438 35760
rect 9125 35751 9183 35757
rect 9125 35748 9137 35751
rect 7432 35720 9137 35748
rect 7432 35708 7438 35720
rect 9125 35717 9137 35720
rect 9171 35717 9183 35751
rect 9125 35711 9183 35717
rect 12710 35680 12716 35692
rect 7300 35652 8432 35680
rect 12671 35652 12716 35680
rect 3513 35615 3571 35621
rect 3513 35581 3525 35615
rect 3559 35581 3571 35615
rect 3513 35575 3571 35581
rect 4430 35572 4436 35624
rect 4488 35612 4494 35624
rect 4525 35615 4583 35621
rect 4525 35612 4537 35615
rect 4488 35584 4537 35612
rect 4488 35572 4494 35584
rect 4525 35581 4537 35584
rect 4571 35581 4583 35615
rect 4706 35612 4712 35624
rect 4667 35584 4712 35612
rect 4525 35575 4583 35581
rect 4706 35572 4712 35584
rect 4764 35572 4770 35624
rect 5169 35615 5227 35621
rect 5169 35581 5181 35615
rect 5215 35581 5227 35615
rect 5169 35575 5227 35581
rect 5261 35615 5319 35621
rect 5261 35581 5273 35615
rect 5307 35581 5319 35615
rect 5261 35575 5319 35581
rect 2682 35504 2688 35556
rect 2740 35544 2746 35556
rect 5184 35544 5212 35575
rect 2740 35516 5212 35544
rect 2740 35504 2746 35516
rect 4706 35436 4712 35488
rect 4764 35476 4770 35488
rect 5276 35476 5304 35575
rect 5626 35572 5632 35624
rect 5684 35612 5690 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 5684 35584 6837 35612
rect 5684 35572 5690 35584
rect 6825 35581 6837 35584
rect 6871 35581 6883 35615
rect 6825 35575 6883 35581
rect 8021 35615 8079 35621
rect 8021 35581 8033 35615
rect 8067 35581 8079 35615
rect 8021 35575 8079 35581
rect 8205 35615 8263 35621
rect 8205 35581 8217 35615
rect 8251 35581 8263 35615
rect 8404 35612 8432 35652
rect 12710 35640 12716 35652
rect 12768 35640 12774 35692
rect 12802 35640 12808 35692
rect 12860 35680 12866 35692
rect 13817 35683 13875 35689
rect 13817 35680 13829 35683
rect 12860 35652 13829 35680
rect 12860 35640 12866 35652
rect 13817 35649 13829 35652
rect 13863 35649 13875 35683
rect 13817 35643 13875 35649
rect 8662 35612 8668 35624
rect 8404 35584 8668 35612
rect 8205 35575 8263 35581
rect 5813 35547 5871 35553
rect 5813 35513 5825 35547
rect 5859 35544 5871 35547
rect 6086 35544 6092 35556
rect 5859 35516 6092 35544
rect 5859 35513 5871 35516
rect 5813 35507 5871 35513
rect 6086 35504 6092 35516
rect 6144 35504 6150 35556
rect 7006 35476 7012 35488
rect 4764 35448 5304 35476
rect 6967 35448 7012 35476
rect 4764 35436 4770 35448
rect 7006 35436 7012 35448
rect 7064 35436 7070 35488
rect 8036 35476 8064 35575
rect 8220 35544 8248 35575
rect 8662 35572 8668 35584
rect 8720 35572 8726 35624
rect 8757 35615 8815 35621
rect 8757 35581 8769 35615
rect 8803 35581 8815 35615
rect 8757 35575 8815 35581
rect 10321 35615 10379 35621
rect 10321 35581 10333 35615
rect 10367 35612 10379 35615
rect 10962 35612 10968 35624
rect 10367 35584 10968 35612
rect 10367 35581 10379 35584
rect 10321 35575 10379 35581
rect 8478 35544 8484 35556
rect 8220 35516 8484 35544
rect 8478 35504 8484 35516
rect 8536 35544 8542 35556
rect 8772 35544 8800 35575
rect 10962 35572 10968 35584
rect 11020 35572 11026 35624
rect 11333 35615 11391 35621
rect 11333 35581 11345 35615
rect 11379 35612 11391 35615
rect 11882 35612 11888 35624
rect 11379 35584 11888 35612
rect 11379 35581 11391 35584
rect 11333 35575 11391 35581
rect 11882 35572 11888 35584
rect 11940 35572 11946 35624
rect 12437 35615 12495 35621
rect 12437 35581 12449 35615
rect 12483 35612 12495 35615
rect 12483 35584 13860 35612
rect 12483 35581 12495 35584
rect 12437 35575 12495 35581
rect 8536 35516 8800 35544
rect 8536 35504 8542 35516
rect 8846 35504 8852 35556
rect 8904 35544 8910 35556
rect 11606 35544 11612 35556
rect 8904 35516 11612 35544
rect 8904 35504 8910 35516
rect 11606 35504 11612 35516
rect 11664 35504 11670 35556
rect 9674 35476 9680 35488
rect 8036 35448 9680 35476
rect 9674 35436 9680 35448
rect 9732 35436 9738 35488
rect 11422 35476 11428 35488
rect 11383 35448 11428 35476
rect 11422 35436 11428 35448
rect 11480 35436 11486 35488
rect 13832 35476 13860 35584
rect 14752 35544 14780 35788
rect 15102 35776 15108 35828
rect 15160 35816 15166 35828
rect 16301 35819 16359 35825
rect 16301 35816 16313 35819
rect 15160 35788 16313 35816
rect 15160 35776 15166 35788
rect 16301 35785 16313 35788
rect 16347 35785 16359 35819
rect 16301 35779 16359 35785
rect 15194 35680 15200 35692
rect 15155 35652 15200 35680
rect 15194 35640 15200 35652
rect 15252 35640 15258 35692
rect 14918 35612 14924 35624
rect 14879 35584 14924 35612
rect 14918 35572 14924 35584
rect 14976 35572 14982 35624
rect 18049 35615 18107 35621
rect 18049 35612 18061 35615
rect 15028 35584 18061 35612
rect 15028 35544 15056 35584
rect 18049 35581 18061 35584
rect 18095 35581 18107 35615
rect 18049 35575 18107 35581
rect 18233 35615 18291 35621
rect 18233 35581 18245 35615
rect 18279 35612 18291 35615
rect 18414 35612 18420 35624
rect 18279 35584 18420 35612
rect 18279 35581 18291 35584
rect 18233 35575 18291 35581
rect 14752 35516 15056 35544
rect 18064 35544 18092 35575
rect 18414 35572 18420 35584
rect 18472 35572 18478 35624
rect 19610 35544 19616 35556
rect 18064 35516 19616 35544
rect 19610 35504 19616 35516
rect 19668 35504 19674 35556
rect 14918 35476 14924 35488
rect 13832 35448 14924 35476
rect 14918 35436 14924 35448
rect 14976 35436 14982 35488
rect 16574 35436 16580 35488
rect 16632 35476 16638 35488
rect 18325 35479 18383 35485
rect 18325 35476 18337 35479
rect 16632 35448 18337 35476
rect 16632 35436 16638 35448
rect 18325 35445 18337 35448
rect 18371 35445 18383 35479
rect 18325 35439 18383 35445
rect 1104 35386 24840 35408
rect 1104 35334 8912 35386
rect 8964 35334 8976 35386
rect 9028 35334 9040 35386
rect 9092 35334 9104 35386
rect 9156 35334 16843 35386
rect 16895 35334 16907 35386
rect 16959 35334 16971 35386
rect 17023 35334 17035 35386
rect 17087 35334 24840 35386
rect 1104 35312 24840 35334
rect 5350 35272 5356 35284
rect 4816 35244 5356 35272
rect 4246 35136 4252 35148
rect 4207 35108 4252 35136
rect 4246 35096 4252 35108
rect 4304 35096 4310 35148
rect 4816 35145 4844 35244
rect 5350 35232 5356 35244
rect 5408 35272 5414 35284
rect 7006 35272 7012 35284
rect 5408 35244 7012 35272
rect 5408 35232 5414 35244
rect 7006 35232 7012 35244
rect 7064 35272 7070 35284
rect 11698 35272 11704 35284
rect 7064 35244 11704 35272
rect 7064 35232 7070 35244
rect 11698 35232 11704 35244
rect 11756 35232 11762 35284
rect 11974 35232 11980 35284
rect 12032 35272 12038 35284
rect 12032 35244 12572 35272
rect 12032 35232 12038 35244
rect 8110 35164 8116 35216
rect 8168 35204 8174 35216
rect 8168 35176 8248 35204
rect 8168 35164 8174 35176
rect 4801 35139 4859 35145
rect 4801 35105 4813 35139
rect 4847 35105 4859 35139
rect 4801 35099 4859 35105
rect 5629 35139 5687 35145
rect 5629 35105 5641 35139
rect 5675 35136 5687 35139
rect 5718 35136 5724 35148
rect 5675 35108 5724 35136
rect 5675 35105 5687 35108
rect 5629 35099 5687 35105
rect 5718 35096 5724 35108
rect 5776 35096 5782 35148
rect 8220 35145 8248 35176
rect 12544 35148 12572 35244
rect 14642 35232 14648 35284
rect 14700 35272 14706 35284
rect 15381 35275 15439 35281
rect 15381 35272 15393 35275
rect 14700 35244 15393 35272
rect 14700 35232 14706 35244
rect 15381 35241 15393 35244
rect 15427 35241 15439 35275
rect 15381 35235 15439 35241
rect 14369 35207 14427 35213
rect 14369 35173 14381 35207
rect 14415 35204 14427 35207
rect 14458 35204 14464 35216
rect 14415 35176 14464 35204
rect 14415 35173 14427 35176
rect 14369 35167 14427 35173
rect 14458 35164 14464 35176
rect 14516 35164 14522 35216
rect 18233 35207 18291 35213
rect 18233 35173 18245 35207
rect 18279 35204 18291 35207
rect 21358 35204 21364 35216
rect 18279 35176 21364 35204
rect 18279 35173 18291 35176
rect 18233 35167 18291 35173
rect 21358 35164 21364 35176
rect 21416 35164 21422 35216
rect 8205 35139 8263 35145
rect 8205 35105 8217 35139
rect 8251 35105 8263 35139
rect 8205 35099 8263 35105
rect 9953 35139 10011 35145
rect 9953 35105 9965 35139
rect 9999 35136 10011 35139
rect 9999 35108 11652 35136
rect 9999 35105 10011 35108
rect 9953 35099 10011 35105
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 5905 35071 5963 35077
rect 2096 35040 4384 35068
rect 2096 35028 2102 35040
rect 4154 34932 4160 34944
rect 4115 34904 4160 34932
rect 4154 34892 4160 34904
rect 4212 34892 4218 34944
rect 4356 34932 4384 35040
rect 5905 35037 5917 35071
rect 5951 35068 5963 35071
rect 5951 35040 7052 35068
rect 5951 35037 5963 35040
rect 5905 35031 5963 35037
rect 7024 35000 7052 35040
rect 7282 35028 7288 35080
rect 7340 35068 7346 35080
rect 8113 35071 8171 35077
rect 8113 35068 8125 35071
rect 7340 35040 8125 35068
rect 7340 35028 7346 35040
rect 8113 35037 8125 35040
rect 8159 35037 8171 35071
rect 10226 35068 10232 35080
rect 10187 35040 10232 35068
rect 8113 35031 8171 35037
rect 10226 35028 10232 35040
rect 10284 35028 10290 35080
rect 11624 35068 11652 35108
rect 12526 35096 12532 35148
rect 12584 35145 12590 35148
rect 12584 35136 12593 35145
rect 13630 35136 13636 35148
rect 12584 35108 12629 35136
rect 13591 35108 13636 35136
rect 12584 35099 12593 35108
rect 12584 35096 12590 35099
rect 13630 35096 13636 35108
rect 13688 35096 13694 35148
rect 15289 35139 15347 35145
rect 15289 35105 15301 35139
rect 15335 35136 15347 35139
rect 16666 35136 16672 35148
rect 15335 35108 16672 35136
rect 15335 35105 15347 35108
rect 15289 35099 15347 35105
rect 16666 35096 16672 35108
rect 16724 35136 16730 35148
rect 17126 35136 17132 35148
rect 16724 35108 17132 35136
rect 16724 35096 16730 35108
rect 17126 35096 17132 35108
rect 17184 35096 17190 35148
rect 11624 35040 12572 35068
rect 12544 35012 12572 35040
rect 13814 35028 13820 35080
rect 13872 35068 13878 35080
rect 14001 35071 14059 35077
rect 14001 35068 14013 35071
rect 13872 35040 14013 35068
rect 13872 35028 13878 35040
rect 14001 35037 14013 35040
rect 14047 35037 14059 35071
rect 14001 35031 14059 35037
rect 14458 35028 14464 35080
rect 14516 35068 14522 35080
rect 14734 35068 14740 35080
rect 14516 35040 14740 35068
rect 14516 35028 14522 35040
rect 14734 35028 14740 35040
rect 14792 35028 14798 35080
rect 16577 35071 16635 35077
rect 16577 35037 16589 35071
rect 16623 35037 16635 35071
rect 16577 35031 16635 35037
rect 16853 35071 16911 35077
rect 16853 35037 16865 35071
rect 16899 35068 16911 35071
rect 18506 35068 18512 35080
rect 16899 35040 18512 35068
rect 16899 35037 16911 35040
rect 16853 35031 16911 35037
rect 7024 34972 8432 35000
rect 8404 34941 8432 34972
rect 11882 34960 11888 35012
rect 11940 35000 11946 35012
rect 11940 34972 12480 35000
rect 11940 34960 11946 34972
rect 7009 34935 7067 34941
rect 7009 34932 7021 34935
rect 4356 34904 7021 34932
rect 7009 34901 7021 34904
rect 7055 34901 7067 34935
rect 7009 34895 7067 34901
rect 8389 34935 8447 34941
rect 8389 34901 8401 34935
rect 8435 34901 8447 34935
rect 8389 34895 8447 34901
rect 11330 34892 11336 34944
rect 11388 34932 11394 34944
rect 11517 34935 11575 34941
rect 11517 34932 11529 34935
rect 11388 34904 11529 34932
rect 11388 34892 11394 34904
rect 11517 34901 11529 34904
rect 11563 34932 11575 34935
rect 11974 34932 11980 34944
rect 11563 34904 11980 34932
rect 11563 34901 11575 34904
rect 11517 34895 11575 34901
rect 11974 34892 11980 34904
rect 12032 34892 12038 34944
rect 12452 34932 12480 34972
rect 12526 34960 12532 35012
rect 12584 34960 12590 35012
rect 13909 35003 13967 35009
rect 13909 35000 13921 35003
rect 12636 34972 13921 35000
rect 12636 34932 12664 34972
rect 13909 34969 13921 34972
rect 13955 35000 13967 35003
rect 15286 35000 15292 35012
rect 13955 34972 15292 35000
rect 13955 34969 13967 34972
rect 13909 34963 13967 34969
rect 15286 34960 15292 34972
rect 15344 34960 15350 35012
rect 12452 34904 12664 34932
rect 12713 34935 12771 34941
rect 12713 34901 12725 34935
rect 12759 34932 12771 34935
rect 13354 34932 13360 34944
rect 12759 34904 13360 34932
rect 12759 34901 12771 34904
rect 12713 34895 12771 34901
rect 13354 34892 13360 34904
rect 13412 34932 13418 34944
rect 13814 34941 13820 34944
rect 13798 34935 13820 34941
rect 13798 34932 13810 34935
rect 13412 34904 13810 34932
rect 13412 34892 13418 34904
rect 13798 34901 13810 34904
rect 13798 34895 13820 34901
rect 13814 34892 13820 34895
rect 13872 34892 13878 34944
rect 16592 34932 16620 35031
rect 18506 35028 18512 35040
rect 18564 35028 18570 35080
rect 17218 34932 17224 34944
rect 16592 34904 17224 34932
rect 17218 34892 17224 34904
rect 17276 34892 17282 34944
rect 1104 34842 24840 34864
rect 1104 34790 4947 34842
rect 4999 34790 5011 34842
rect 5063 34790 5075 34842
rect 5127 34790 5139 34842
rect 5191 34790 12878 34842
rect 12930 34790 12942 34842
rect 12994 34790 13006 34842
rect 13058 34790 13070 34842
rect 13122 34790 20808 34842
rect 20860 34790 20872 34842
rect 20924 34790 20936 34842
rect 20988 34790 21000 34842
rect 21052 34790 24840 34842
rect 1104 34768 24840 34790
rect 2777 34731 2835 34737
rect 2777 34697 2789 34731
rect 2823 34728 2835 34731
rect 4338 34728 4344 34740
rect 2823 34700 4344 34728
rect 2823 34697 2835 34700
rect 2777 34691 2835 34697
rect 4338 34688 4344 34700
rect 4396 34688 4402 34740
rect 6454 34688 6460 34740
rect 6512 34728 6518 34740
rect 6822 34728 6828 34740
rect 6512 34700 6828 34728
rect 6512 34688 6518 34700
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 9306 34728 9312 34740
rect 6932 34700 9312 34728
rect 5626 34660 5632 34672
rect 2976 34632 5632 34660
rect 2590 34484 2596 34536
rect 2648 34524 2654 34536
rect 2976 34524 3004 34632
rect 5626 34620 5632 34632
rect 5684 34620 5690 34672
rect 3050 34552 3056 34604
rect 3108 34592 3114 34604
rect 3237 34595 3295 34601
rect 3237 34592 3249 34595
rect 3108 34564 3249 34592
rect 3108 34552 3114 34564
rect 3237 34561 3249 34564
rect 3283 34592 3295 34595
rect 5813 34595 5871 34601
rect 3283 34564 4936 34592
rect 3283 34561 3295 34564
rect 3237 34555 3295 34561
rect 3145 34527 3203 34533
rect 3145 34524 3157 34527
rect 2648 34496 3157 34524
rect 2648 34484 2654 34496
rect 3145 34493 3157 34496
rect 3191 34493 3203 34527
rect 3145 34487 3203 34493
rect 3513 34527 3571 34533
rect 3513 34493 3525 34527
rect 3559 34493 3571 34527
rect 3513 34487 3571 34493
rect 3697 34527 3755 34533
rect 3697 34493 3709 34527
rect 3743 34524 3755 34527
rect 4062 34524 4068 34536
rect 3743 34496 4068 34524
rect 3743 34493 3755 34496
rect 3697 34487 3755 34493
rect 2958 34348 2964 34400
rect 3016 34388 3022 34400
rect 3528 34388 3556 34487
rect 4062 34484 4068 34496
rect 4120 34484 4126 34536
rect 4522 34524 4528 34536
rect 4483 34496 4528 34524
rect 4522 34484 4528 34496
rect 4580 34484 4586 34536
rect 4706 34524 4712 34536
rect 4619 34496 4712 34524
rect 4706 34484 4712 34496
rect 4764 34484 4770 34536
rect 4908 34524 4936 34564
rect 5813 34561 5825 34595
rect 5859 34592 5871 34595
rect 6454 34592 6460 34604
rect 5859 34564 6460 34592
rect 5859 34561 5871 34564
rect 5813 34555 5871 34561
rect 6454 34552 6460 34564
rect 6512 34552 6518 34604
rect 6932 34601 6960 34700
rect 9306 34688 9312 34700
rect 9364 34688 9370 34740
rect 10226 34728 10232 34740
rect 10187 34700 10232 34728
rect 10226 34688 10232 34700
rect 10284 34688 10290 34740
rect 11422 34688 11428 34740
rect 11480 34728 11486 34740
rect 12575 34731 12633 34737
rect 12575 34728 12587 34731
rect 11480 34700 12587 34728
rect 11480 34688 11486 34700
rect 12575 34697 12587 34700
rect 12621 34697 12633 34731
rect 12575 34691 12633 34697
rect 12713 34731 12771 34737
rect 12713 34697 12725 34731
rect 12759 34728 12771 34731
rect 13170 34728 13176 34740
rect 12759 34700 13176 34728
rect 12759 34697 12771 34700
rect 12713 34691 12771 34697
rect 13170 34688 13176 34700
rect 13228 34688 13234 34740
rect 16022 34688 16028 34740
rect 16080 34728 16086 34740
rect 18049 34731 18107 34737
rect 18049 34728 18061 34731
rect 16080 34700 18061 34728
rect 16080 34688 16086 34700
rect 18049 34697 18061 34700
rect 18095 34697 18107 34731
rect 18506 34728 18512 34740
rect 18467 34700 18512 34728
rect 18049 34691 18107 34697
rect 18506 34688 18512 34700
rect 18564 34688 18570 34740
rect 8294 34660 8300 34672
rect 7024 34632 8300 34660
rect 6917 34595 6975 34601
rect 6917 34561 6929 34595
rect 6963 34561 6975 34595
rect 6917 34555 6975 34561
rect 5169 34527 5227 34533
rect 5169 34524 5181 34527
rect 4908 34496 5181 34524
rect 5169 34493 5181 34496
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 5258 34484 5264 34536
rect 5316 34524 5322 34536
rect 7024 34533 7052 34632
rect 8294 34620 8300 34632
rect 8352 34620 8358 34672
rect 9858 34660 9864 34672
rect 9232 34632 9864 34660
rect 7009 34527 7067 34533
rect 5316 34496 5361 34524
rect 5316 34484 5322 34496
rect 7009 34493 7021 34527
rect 7055 34493 7067 34527
rect 7466 34524 7472 34536
rect 7427 34496 7472 34524
rect 7009 34487 7067 34493
rect 7466 34484 7472 34496
rect 7524 34484 7530 34536
rect 7558 34484 7564 34536
rect 7616 34524 7622 34536
rect 8478 34524 8484 34536
rect 7616 34496 8484 34524
rect 7616 34484 7622 34496
rect 8478 34484 8484 34496
rect 8536 34484 8542 34536
rect 9232 34533 9260 34632
rect 9858 34620 9864 34632
rect 9916 34620 9922 34672
rect 14093 34663 14151 34669
rect 14093 34660 14105 34663
rect 12820 34632 14105 34660
rect 12820 34604 12848 34632
rect 14093 34629 14105 34632
rect 14139 34629 14151 34663
rect 14093 34623 14151 34629
rect 12802 34592 12808 34604
rect 12715 34564 12808 34592
rect 12802 34552 12808 34564
rect 12860 34552 12866 34604
rect 12897 34595 12955 34601
rect 12897 34561 12909 34595
rect 12943 34561 12955 34595
rect 12897 34555 12955 34561
rect 15565 34595 15623 34601
rect 15565 34561 15577 34595
rect 15611 34592 15623 34595
rect 16298 34592 16304 34604
rect 15611 34564 16304 34592
rect 15611 34561 15623 34564
rect 15565 34555 15623 34561
rect 9217 34527 9275 34533
rect 9217 34493 9229 34527
rect 9263 34493 9275 34527
rect 9217 34487 9275 34493
rect 9306 34484 9312 34536
rect 9364 34524 9370 34536
rect 9677 34527 9735 34533
rect 9364 34496 9409 34524
rect 9364 34484 9370 34496
rect 9677 34493 9689 34527
rect 9723 34493 9735 34527
rect 9677 34487 9735 34493
rect 4724 34456 4752 34484
rect 5276 34456 5304 34484
rect 4724 34428 5304 34456
rect 9692 34456 9720 34487
rect 9766 34484 9772 34536
rect 9824 34524 9830 34536
rect 9950 34524 9956 34536
rect 9824 34496 9956 34524
rect 9824 34484 9830 34496
rect 9950 34484 9956 34496
rect 10008 34484 10014 34536
rect 11330 34524 11336 34536
rect 11291 34496 11336 34524
rect 11330 34484 11336 34496
rect 11388 34484 11394 34536
rect 11425 34527 11483 34533
rect 11425 34493 11437 34527
rect 11471 34493 11483 34527
rect 11425 34487 11483 34493
rect 10134 34456 10140 34468
rect 9692 34428 10140 34456
rect 10134 34416 10140 34428
rect 10192 34456 10198 34468
rect 11440 34456 11468 34487
rect 12618 34484 12624 34536
rect 12676 34524 12682 34536
rect 12912 34524 12940 34555
rect 16298 34552 16304 34564
rect 16356 34552 16362 34604
rect 16390 34552 16396 34604
rect 16448 34592 16454 34604
rect 16448 34564 18368 34592
rect 16448 34552 16454 34564
rect 13998 34524 14004 34536
rect 12676 34496 12940 34524
rect 13959 34496 14004 34524
rect 12676 34484 12682 34496
rect 13998 34484 14004 34496
rect 14056 34484 14062 34536
rect 15473 34527 15531 34533
rect 15473 34493 15485 34527
rect 15519 34524 15531 34527
rect 15654 34524 15660 34536
rect 15519 34496 15660 34524
rect 15519 34493 15531 34496
rect 15473 34487 15531 34493
rect 15654 34484 15660 34496
rect 15712 34484 15718 34536
rect 15746 34484 15752 34536
rect 15804 34524 15810 34536
rect 18340 34533 18368 34564
rect 18325 34527 18383 34533
rect 15804 34496 15849 34524
rect 15804 34484 15810 34496
rect 18325 34493 18337 34527
rect 18371 34493 18383 34527
rect 18325 34487 18383 34493
rect 19797 34527 19855 34533
rect 19797 34493 19809 34527
rect 19843 34524 19855 34527
rect 21358 34524 21364 34536
rect 19843 34496 21364 34524
rect 19843 34493 19855 34496
rect 19797 34487 19855 34493
rect 21358 34484 21364 34496
rect 21416 34484 21422 34536
rect 12437 34459 12495 34465
rect 12437 34456 12449 34459
rect 10192 34428 12449 34456
rect 10192 34416 10198 34428
rect 12437 34425 12449 34428
rect 12483 34425 12495 34459
rect 12437 34419 12495 34425
rect 18233 34459 18291 34465
rect 18233 34425 18245 34459
rect 18279 34425 18291 34459
rect 19610 34456 19616 34468
rect 19571 34428 19616 34456
rect 18233 34419 18291 34425
rect 5534 34388 5540 34400
rect 3016 34360 5540 34388
rect 3016 34348 3022 34360
rect 5534 34348 5540 34360
rect 5592 34348 5598 34400
rect 7742 34348 7748 34400
rect 7800 34388 7806 34400
rect 8021 34391 8079 34397
rect 8021 34388 8033 34391
rect 7800 34360 8033 34388
rect 7800 34348 7806 34360
rect 8021 34357 8033 34360
rect 8067 34357 8079 34391
rect 18248 34388 18276 34419
rect 19610 34416 19616 34428
rect 19668 34416 19674 34468
rect 19889 34391 19947 34397
rect 19889 34388 19901 34391
rect 18248 34360 19901 34388
rect 8021 34351 8079 34357
rect 19889 34357 19901 34360
rect 19935 34357 19947 34391
rect 19889 34351 19947 34357
rect 1104 34298 24840 34320
rect 1104 34246 8912 34298
rect 8964 34246 8976 34298
rect 9028 34246 9040 34298
rect 9092 34246 9104 34298
rect 9156 34246 16843 34298
rect 16895 34246 16907 34298
rect 16959 34246 16971 34298
rect 17023 34246 17035 34298
rect 17087 34246 24840 34298
rect 1104 34224 24840 34246
rect 2225 34187 2283 34193
rect 2225 34153 2237 34187
rect 2271 34184 2283 34187
rect 3694 34184 3700 34196
rect 2271 34156 3700 34184
rect 2271 34153 2283 34156
rect 2225 34147 2283 34153
rect 3694 34144 3700 34156
rect 3752 34144 3758 34196
rect 4893 34187 4951 34193
rect 4893 34153 4905 34187
rect 4939 34184 4951 34187
rect 7466 34184 7472 34196
rect 4939 34156 7472 34184
rect 4939 34153 4951 34156
rect 4893 34147 4951 34153
rect 7466 34144 7472 34156
rect 7524 34144 7530 34196
rect 8478 34184 8484 34196
rect 8439 34156 8484 34184
rect 8478 34144 8484 34156
rect 8536 34144 8542 34196
rect 9950 34184 9956 34196
rect 9911 34156 9956 34184
rect 9950 34144 9956 34156
rect 10008 34144 10014 34196
rect 11054 34184 11060 34196
rect 11015 34156 11060 34184
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 12989 34187 13047 34193
rect 12989 34184 13001 34187
rect 12492 34156 13001 34184
rect 12492 34144 12498 34156
rect 12989 34153 13001 34156
rect 13035 34153 13047 34187
rect 12989 34147 13047 34153
rect 11422 34076 11428 34128
rect 11480 34116 11486 34128
rect 18233 34119 18291 34125
rect 11480 34088 12020 34116
rect 11480 34076 11486 34088
rect 2590 34048 2596 34060
rect 2551 34020 2596 34048
rect 2590 34008 2596 34020
rect 2648 34008 2654 34060
rect 2958 34048 2964 34060
rect 2919 34020 2964 34048
rect 2958 34008 2964 34020
rect 3016 34008 3022 34060
rect 3142 34048 3148 34060
rect 3103 34020 3148 34048
rect 3142 34008 3148 34020
rect 3200 34008 3206 34060
rect 4801 34051 4859 34057
rect 4801 34017 4813 34051
rect 4847 34048 4859 34051
rect 5902 34048 5908 34060
rect 4847 34020 5908 34048
rect 4847 34017 4859 34020
rect 4801 34011 4859 34017
rect 5902 34008 5908 34020
rect 5960 34008 5966 34060
rect 6086 34048 6092 34060
rect 6047 34020 6092 34048
rect 6086 34008 6092 34020
rect 6144 34008 6150 34060
rect 8294 34048 8300 34060
rect 8255 34020 8300 34048
rect 8294 34008 8300 34020
rect 8352 34008 8358 34060
rect 9769 34051 9827 34057
rect 9769 34017 9781 34051
rect 9815 34048 9827 34051
rect 9858 34048 9864 34060
rect 9815 34020 9864 34048
rect 9815 34017 9827 34020
rect 9769 34011 9827 34017
rect 9858 34008 9864 34020
rect 9916 34048 9922 34060
rect 10410 34048 10416 34060
rect 9916 34020 10416 34048
rect 9916 34008 9922 34020
rect 10410 34008 10416 34020
rect 10468 34008 10474 34060
rect 11238 34008 11244 34060
rect 11296 34048 11302 34060
rect 11992 34057 12020 34088
rect 18233 34085 18245 34119
rect 18279 34116 18291 34119
rect 18414 34116 18420 34128
rect 18279 34088 18420 34116
rect 18279 34085 18291 34088
rect 18233 34079 18291 34085
rect 18414 34076 18420 34088
rect 18472 34076 18478 34128
rect 11609 34051 11667 34057
rect 11609 34048 11621 34051
rect 11296 34020 11621 34048
rect 11296 34008 11302 34020
rect 11609 34017 11621 34020
rect 11655 34017 11667 34051
rect 11609 34011 11667 34017
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34017 12035 34051
rect 11977 34011 12035 34017
rect 12161 34051 12219 34057
rect 12161 34017 12173 34051
rect 12207 34048 12219 34051
rect 12434 34048 12440 34060
rect 12207 34020 12440 34048
rect 12207 34017 12219 34020
rect 12161 34011 12219 34017
rect 2682 33980 2688 33992
rect 2643 33952 2688 33980
rect 2682 33940 2688 33952
rect 2740 33940 2746 33992
rect 5718 33940 5724 33992
rect 5776 33980 5782 33992
rect 5813 33983 5871 33989
rect 5813 33980 5825 33983
rect 5776 33952 5825 33980
rect 5776 33940 5782 33952
rect 5813 33949 5825 33952
rect 5859 33949 5871 33983
rect 5813 33943 5871 33949
rect 10594 33940 10600 33992
rect 10652 33980 10658 33992
rect 11425 33983 11483 33989
rect 11425 33980 11437 33983
rect 10652 33952 11437 33980
rect 10652 33940 10658 33952
rect 11425 33949 11437 33952
rect 11471 33949 11483 33983
rect 11425 33943 11483 33949
rect 10042 33872 10048 33924
rect 10100 33912 10106 33924
rect 11054 33912 11060 33924
rect 10100 33884 11060 33912
rect 10100 33872 10106 33884
rect 11054 33872 11060 33884
rect 11112 33872 11118 33924
rect 11624 33912 11652 34011
rect 12434 34008 12440 34020
rect 12492 34048 12498 34060
rect 12802 34048 12808 34060
rect 12492 34020 12808 34048
rect 12492 34008 12498 34020
rect 12802 34008 12808 34020
rect 12860 34008 12866 34060
rect 13173 34051 13231 34057
rect 13173 34017 13185 34051
rect 13219 34017 13231 34051
rect 13173 34011 13231 34017
rect 13909 34051 13967 34057
rect 13909 34017 13921 34051
rect 13955 34017 13967 34051
rect 13909 34011 13967 34017
rect 14369 34051 14427 34057
rect 14369 34017 14381 34051
rect 14415 34048 14427 34051
rect 15746 34048 15752 34060
rect 14415 34020 15752 34048
rect 14415 34017 14427 34020
rect 14369 34011 14427 34017
rect 11882 33940 11888 33992
rect 11940 33980 11946 33992
rect 13188 33980 13216 34011
rect 11940 33952 13216 33980
rect 11940 33940 11946 33952
rect 12158 33912 12164 33924
rect 11624 33884 12164 33912
rect 12158 33872 12164 33884
rect 12216 33872 12222 33924
rect 13924 33912 13952 34011
rect 15746 34008 15752 34020
rect 15804 34008 15810 34060
rect 16577 34051 16635 34057
rect 16577 34017 16589 34051
rect 16623 34048 16635 34051
rect 17218 34048 17224 34060
rect 16623 34020 17224 34048
rect 16623 34017 16635 34020
rect 16577 34011 16635 34017
rect 14001 33983 14059 33989
rect 14001 33949 14013 33983
rect 14047 33980 14059 33983
rect 16390 33980 16396 33992
rect 14047 33952 16396 33980
rect 14047 33949 14059 33952
rect 14001 33943 14059 33949
rect 16390 33940 16396 33952
rect 16448 33940 16454 33992
rect 14734 33912 14740 33924
rect 13924 33884 14740 33912
rect 14734 33872 14740 33884
rect 14792 33872 14798 33924
rect 15286 33872 15292 33924
rect 15344 33912 15350 33924
rect 16592 33912 16620 34011
rect 17218 34008 17224 34020
rect 17276 34008 17282 34060
rect 16758 33940 16764 33992
rect 16816 33980 16822 33992
rect 16853 33983 16911 33989
rect 16853 33980 16865 33983
rect 16816 33952 16865 33980
rect 16816 33940 16822 33952
rect 16853 33949 16865 33952
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 15344 33884 16620 33912
rect 15344 33872 15350 33884
rect 1946 33804 1952 33856
rect 2004 33844 2010 33856
rect 7190 33844 7196 33856
rect 2004 33816 7196 33844
rect 2004 33804 2010 33816
rect 7190 33804 7196 33816
rect 7248 33804 7254 33856
rect 1104 33754 24840 33776
rect 1104 33702 4947 33754
rect 4999 33702 5011 33754
rect 5063 33702 5075 33754
rect 5127 33702 5139 33754
rect 5191 33702 12878 33754
rect 12930 33702 12942 33754
rect 12994 33702 13006 33754
rect 13058 33702 13070 33754
rect 13122 33702 20808 33754
rect 20860 33702 20872 33754
rect 20924 33702 20936 33754
rect 20988 33702 21000 33754
rect 21052 33702 24840 33754
rect 1104 33680 24840 33702
rect 5902 33600 5908 33652
rect 5960 33640 5966 33652
rect 8849 33643 8907 33649
rect 8849 33640 8861 33643
rect 5960 33612 8861 33640
rect 5960 33600 5966 33612
rect 8849 33609 8861 33612
rect 8895 33609 8907 33643
rect 13998 33640 14004 33652
rect 13959 33612 14004 33640
rect 8849 33603 8907 33609
rect 5718 33572 5724 33584
rect 4540 33544 5724 33572
rect 1486 33464 1492 33516
rect 1544 33504 1550 33516
rect 2225 33507 2283 33513
rect 2225 33504 2237 33507
rect 1544 33476 2237 33504
rect 1544 33464 1550 33476
rect 2225 33473 2237 33476
rect 2271 33504 2283 33507
rect 4540 33504 4568 33544
rect 5718 33532 5724 33544
rect 5776 33532 5782 33584
rect 8864 33572 8892 33603
rect 13998 33600 14004 33612
rect 14056 33600 14062 33652
rect 16022 33640 16028 33652
rect 15983 33612 16028 33640
rect 16022 33600 16028 33612
rect 16080 33600 16086 33652
rect 11514 33572 11520 33584
rect 8864 33544 11520 33572
rect 11514 33532 11520 33544
rect 11572 33532 11578 33584
rect 2271 33476 4568 33504
rect 2271 33473 2283 33476
rect 2225 33467 2283 33473
rect 4614 33464 4620 33516
rect 4672 33504 4678 33516
rect 4709 33507 4767 33513
rect 4709 33504 4721 33507
rect 4672 33476 4721 33504
rect 4672 33464 4678 33476
rect 4709 33473 4721 33476
rect 4755 33473 4767 33507
rect 5629 33507 5687 33513
rect 5629 33504 5641 33507
rect 4709 33467 4767 33473
rect 4816 33476 5641 33504
rect 2501 33439 2559 33445
rect 2501 33405 2513 33439
rect 2547 33436 2559 33439
rect 3970 33436 3976 33448
rect 2547 33408 3976 33436
rect 2547 33405 2559 33408
rect 2501 33399 2559 33405
rect 3970 33396 3976 33408
rect 4028 33396 4034 33448
rect 4154 33396 4160 33448
rect 4212 33436 4218 33448
rect 4816 33436 4844 33476
rect 5629 33473 5641 33476
rect 5675 33473 5687 33507
rect 7742 33504 7748 33516
rect 7703 33476 7748 33504
rect 5629 33467 5687 33473
rect 7742 33464 7748 33476
rect 7800 33464 7806 33516
rect 16758 33504 16764 33516
rect 16719 33476 16764 33504
rect 16758 33464 16764 33476
rect 16816 33464 16822 33516
rect 4212 33408 4844 33436
rect 5169 33439 5227 33445
rect 4212 33396 4218 33408
rect 5169 33405 5181 33439
rect 5215 33405 5227 33439
rect 5169 33399 5227 33405
rect 5353 33439 5411 33445
rect 5353 33405 5365 33439
rect 5399 33436 5411 33439
rect 5399 33408 5488 33436
rect 5399 33405 5411 33408
rect 5353 33399 5411 33405
rect 5184 33368 5212 33399
rect 5460 33368 5488 33408
rect 5534 33396 5540 33448
rect 5592 33436 5598 33448
rect 5721 33439 5779 33445
rect 5721 33436 5733 33439
rect 5592 33408 5733 33436
rect 5592 33396 5598 33408
rect 5721 33405 5733 33408
rect 5767 33405 5779 33439
rect 5721 33399 5779 33405
rect 5626 33368 5632 33380
rect 5184 33340 5396 33368
rect 5460 33340 5632 33368
rect 5368 33312 5396 33340
rect 5626 33328 5632 33340
rect 5684 33328 5690 33380
rect 3694 33260 3700 33312
rect 3752 33300 3758 33312
rect 3789 33303 3847 33309
rect 3789 33300 3801 33303
rect 3752 33272 3801 33300
rect 3752 33260 3758 33272
rect 3789 33269 3801 33272
rect 3835 33269 3847 33303
rect 3789 33263 3847 33269
rect 5350 33260 5356 33312
rect 5408 33260 5414 33312
rect 5534 33260 5540 33312
rect 5592 33300 5598 33312
rect 5736 33300 5764 33399
rect 6178 33396 6184 33448
rect 6236 33436 6242 33448
rect 7469 33439 7527 33445
rect 7469 33436 7481 33439
rect 6236 33408 7481 33436
rect 6236 33396 6242 33408
rect 7469 33405 7481 33408
rect 7515 33405 7527 33439
rect 7469 33399 7527 33405
rect 10042 33396 10048 33448
rect 10100 33436 10106 33448
rect 10137 33439 10195 33445
rect 10137 33436 10149 33439
rect 10100 33408 10149 33436
rect 10100 33396 10106 33408
rect 10137 33405 10149 33408
rect 10183 33405 10195 33439
rect 10137 33399 10195 33405
rect 10152 33368 10180 33399
rect 10226 33396 10232 33448
rect 10284 33436 10290 33448
rect 10594 33436 10600 33448
rect 10284 33408 10329 33436
rect 10555 33408 10600 33436
rect 10284 33396 10290 33408
rect 10594 33396 10600 33408
rect 10652 33396 10658 33448
rect 10689 33439 10747 33445
rect 10689 33405 10701 33439
rect 10735 33405 10747 33439
rect 10689 33399 10747 33405
rect 12437 33439 12495 33445
rect 12437 33405 12449 33439
rect 12483 33436 12495 33439
rect 12526 33436 12532 33448
rect 12483 33408 12532 33436
rect 12483 33405 12495 33408
rect 12437 33399 12495 33405
rect 10704 33368 10732 33399
rect 12526 33396 12532 33408
rect 12584 33396 12590 33448
rect 12710 33436 12716 33448
rect 12671 33408 12716 33436
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 14918 33436 14924 33448
rect 14879 33408 14924 33436
rect 14918 33396 14924 33408
rect 14976 33396 14982 33448
rect 16298 33436 16304 33448
rect 16259 33408 16304 33436
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 10152 33340 10732 33368
rect 16209 33371 16267 33377
rect 16209 33337 16221 33371
rect 16255 33368 16267 33371
rect 16574 33368 16580 33380
rect 16255 33340 16580 33368
rect 16255 33337 16267 33340
rect 16209 33331 16267 33337
rect 16574 33328 16580 33340
rect 16632 33328 16638 33380
rect 5592 33272 5764 33300
rect 5592 33260 5598 33272
rect 5902 33260 5908 33312
rect 5960 33300 5966 33312
rect 8754 33300 8760 33312
rect 5960 33272 8760 33300
rect 5960 33260 5966 33272
rect 8754 33260 8760 33272
rect 8812 33260 8818 33312
rect 9674 33260 9680 33312
rect 9732 33300 9738 33312
rect 11149 33303 11207 33309
rect 11149 33300 11161 33303
rect 9732 33272 11161 33300
rect 9732 33260 9738 33272
rect 11149 33269 11161 33272
rect 11195 33269 11207 33303
rect 15010 33300 15016 33312
rect 14971 33272 15016 33300
rect 11149 33263 11207 33269
rect 15010 33260 15016 33272
rect 15068 33260 15074 33312
rect 1104 33210 24840 33232
rect 1104 33158 8912 33210
rect 8964 33158 8976 33210
rect 9028 33158 9040 33210
rect 9092 33158 9104 33210
rect 9156 33158 16843 33210
rect 16895 33158 16907 33210
rect 16959 33158 16971 33210
rect 17023 33158 17035 33210
rect 17087 33158 24840 33210
rect 1104 33136 24840 33158
rect 2041 33099 2099 33105
rect 2041 33065 2053 33099
rect 2087 33096 2099 33099
rect 2682 33096 2688 33108
rect 2087 33068 2688 33096
rect 2087 33065 2099 33068
rect 2041 33059 2099 33065
rect 2682 33056 2688 33068
rect 2740 33056 2746 33108
rect 3050 33096 3056 33108
rect 3011 33068 3056 33096
rect 3050 33056 3056 33068
rect 3108 33056 3114 33108
rect 4062 33056 4068 33108
rect 4120 33096 4126 33108
rect 4157 33099 4215 33105
rect 4157 33096 4169 33099
rect 4120 33068 4169 33096
rect 4120 33056 4126 33068
rect 4157 33065 4169 33068
rect 4203 33065 4215 33099
rect 7374 33096 7380 33108
rect 4157 33059 4215 33065
rect 6104 33068 7380 33096
rect 6104 33028 6132 33068
rect 7374 33056 7380 33068
rect 7432 33056 7438 33108
rect 8665 33099 8723 33105
rect 8665 33065 8677 33099
rect 8711 33096 8723 33099
rect 10594 33096 10600 33108
rect 8711 33068 10600 33096
rect 8711 33065 8723 33068
rect 8665 33059 8723 33065
rect 10594 33056 10600 33068
rect 10652 33056 10658 33108
rect 12345 33099 12403 33105
rect 12345 33065 12357 33099
rect 12391 33096 12403 33099
rect 12710 33096 12716 33108
rect 12391 33068 12716 33096
rect 12391 33065 12403 33068
rect 12345 33059 12403 33065
rect 12710 33056 12716 33068
rect 12768 33056 12774 33108
rect 2976 33000 6132 33028
rect 13633 33031 13691 33037
rect 1946 32960 1952 32972
rect 1907 32932 1952 32960
rect 1946 32920 1952 32932
rect 2004 32920 2010 32972
rect 2976 32969 3004 33000
rect 13633 32997 13645 33031
rect 13679 33028 13691 33031
rect 15194 33028 15200 33040
rect 13679 33000 15200 33028
rect 13679 32997 13691 33000
rect 13633 32991 13691 32997
rect 15194 32988 15200 33000
rect 15252 32988 15258 33040
rect 2961 32963 3019 32969
rect 2961 32929 2973 32963
rect 3007 32929 3019 32963
rect 2961 32923 3019 32929
rect 3694 32920 3700 32972
rect 3752 32960 3758 32972
rect 4065 32963 4123 32969
rect 4065 32960 4077 32963
rect 3752 32932 4077 32960
rect 3752 32920 3758 32932
rect 4065 32929 4077 32932
rect 4111 32929 4123 32963
rect 4065 32923 4123 32929
rect 5902 32920 5908 32972
rect 5960 32960 5966 32972
rect 8573 32963 8631 32969
rect 5960 32932 6005 32960
rect 5960 32920 5966 32932
rect 8573 32929 8585 32963
rect 8619 32929 8631 32963
rect 8573 32923 8631 32929
rect 9677 32963 9735 32969
rect 9677 32929 9689 32963
rect 9723 32960 9735 32963
rect 9766 32960 9772 32972
rect 9723 32932 9772 32960
rect 9723 32929 9735 32932
rect 9677 32923 9735 32929
rect 4522 32852 4528 32904
rect 4580 32892 4586 32904
rect 4706 32892 4712 32904
rect 4580 32864 4712 32892
rect 4580 32852 4586 32864
rect 4706 32852 4712 32864
rect 4764 32852 4770 32904
rect 5997 32895 6055 32901
rect 5997 32861 6009 32895
rect 6043 32892 6055 32895
rect 6178 32892 6184 32904
rect 6043 32864 6184 32892
rect 6043 32861 6055 32864
rect 5997 32855 6055 32861
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 6273 32895 6331 32901
rect 6273 32861 6285 32895
rect 6319 32892 6331 32895
rect 6454 32892 6460 32904
rect 6319 32864 6460 32892
rect 6319 32861 6331 32864
rect 6273 32855 6331 32861
rect 6454 32852 6460 32864
rect 6512 32852 6518 32904
rect 8588 32892 8616 32923
rect 9766 32920 9772 32932
rect 9824 32920 9830 32972
rect 9861 32963 9919 32969
rect 9861 32929 9873 32963
rect 9907 32960 9919 32963
rect 9907 32932 10180 32960
rect 9907 32929 9919 32932
rect 9861 32923 9919 32929
rect 9950 32892 9956 32904
rect 8588 32864 9956 32892
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 10152 32892 10180 32932
rect 10226 32920 10232 32972
rect 10284 32960 10290 32972
rect 10686 32960 10692 32972
rect 10284 32932 10692 32960
rect 10284 32920 10290 32932
rect 10686 32920 10692 32932
rect 10744 32960 10750 32972
rect 11149 32963 11207 32969
rect 11149 32960 11161 32963
rect 10744 32932 11161 32960
rect 10744 32920 10750 32932
rect 11149 32929 11161 32932
rect 11195 32929 11207 32963
rect 11330 32960 11336 32972
rect 11243 32932 11336 32960
rect 11149 32923 11207 32929
rect 11330 32920 11336 32932
rect 11388 32960 11394 32972
rect 11885 32963 11943 32969
rect 11885 32960 11897 32963
rect 11388 32932 11897 32960
rect 11388 32920 11394 32932
rect 11885 32929 11897 32932
rect 11931 32929 11943 32963
rect 11885 32923 11943 32929
rect 12069 32963 12127 32969
rect 12069 32929 12081 32963
rect 12115 32960 12127 32963
rect 12434 32960 12440 32972
rect 12115 32932 12440 32960
rect 12115 32929 12127 32932
rect 12069 32923 12127 32929
rect 12434 32920 12440 32932
rect 12492 32920 12498 32972
rect 13538 32960 13544 32972
rect 13499 32932 13544 32960
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 14182 32960 14188 32972
rect 14016 32932 14188 32960
rect 10962 32892 10968 32904
rect 10152 32864 10968 32892
rect 10962 32852 10968 32864
rect 11020 32852 11026 32904
rect 14016 32901 14044 32932
rect 14182 32920 14188 32932
rect 14240 32920 14246 32972
rect 15010 32920 15016 32972
rect 15068 32960 15074 32972
rect 15933 32963 15991 32969
rect 15933 32960 15945 32963
rect 15068 32932 15945 32960
rect 15068 32920 15074 32932
rect 15933 32929 15945 32932
rect 15979 32929 15991 32963
rect 15933 32923 15991 32929
rect 16301 32963 16359 32969
rect 16301 32929 16313 32963
rect 16347 32929 16359 32963
rect 16301 32923 16359 32929
rect 16485 32963 16543 32969
rect 16485 32929 16497 32963
rect 16531 32960 16543 32963
rect 16666 32960 16672 32972
rect 16531 32932 16672 32960
rect 16531 32929 16543 32932
rect 16485 32923 16543 32929
rect 14001 32895 14059 32901
rect 14001 32861 14013 32895
rect 14047 32861 14059 32895
rect 14001 32855 14059 32861
rect 14090 32852 14096 32904
rect 14148 32892 14154 32904
rect 15378 32892 15384 32904
rect 14148 32864 14193 32892
rect 14936 32864 15384 32892
rect 14148 32852 14154 32864
rect 13906 32824 13912 32836
rect 13867 32796 13912 32824
rect 13906 32784 13912 32796
rect 13964 32784 13970 32836
rect 14936 32824 14964 32864
rect 15378 32852 15384 32864
rect 15436 32852 15442 32904
rect 15838 32892 15844 32904
rect 15799 32864 15844 32892
rect 15838 32852 15844 32864
rect 15896 32852 15902 32904
rect 16316 32892 16344 32923
rect 16666 32920 16672 32932
rect 16724 32920 16730 32972
rect 16574 32892 16580 32904
rect 16316 32864 16580 32892
rect 16574 32852 16580 32864
rect 16632 32852 16638 32904
rect 14016 32796 14964 32824
rect 5718 32756 5724 32768
rect 5679 32728 5724 32756
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 9858 32716 9864 32768
rect 9916 32756 9922 32768
rect 9953 32759 10011 32765
rect 9953 32756 9965 32759
rect 9916 32728 9965 32756
rect 9916 32716 9922 32728
rect 9953 32725 9965 32728
rect 9999 32725 10011 32759
rect 13354 32756 13360 32768
rect 13315 32728 13360 32756
rect 9953 32719 10011 32725
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13814 32765 13820 32768
rect 13798 32759 13820 32765
rect 13798 32725 13810 32759
rect 13872 32756 13878 32768
rect 14016 32756 14044 32796
rect 15378 32756 15384 32768
rect 13872 32728 14044 32756
rect 15339 32728 15384 32756
rect 13798 32719 13820 32725
rect 13814 32716 13820 32719
rect 13872 32716 13878 32728
rect 15378 32716 15384 32728
rect 15436 32716 15442 32768
rect 1104 32666 24840 32688
rect 1104 32614 4947 32666
rect 4999 32614 5011 32666
rect 5063 32614 5075 32666
rect 5127 32614 5139 32666
rect 5191 32614 12878 32666
rect 12930 32614 12942 32666
rect 12994 32614 13006 32666
rect 13058 32614 13070 32666
rect 13122 32614 20808 32666
rect 20860 32614 20872 32666
rect 20924 32614 20936 32666
rect 20988 32614 21000 32666
rect 21052 32614 24840 32666
rect 1104 32592 24840 32614
rect 14090 32552 14096 32564
rect 1504 32524 14096 32552
rect 1504 32357 1532 32524
rect 14090 32512 14096 32524
rect 14148 32512 14154 32564
rect 3970 32484 3976 32496
rect 3931 32456 3976 32484
rect 3970 32444 3976 32456
rect 4028 32444 4034 32496
rect 5810 32444 5816 32496
rect 5868 32484 5874 32496
rect 6181 32487 6239 32493
rect 6181 32484 6193 32487
rect 5868 32456 6193 32484
rect 5868 32444 5874 32456
rect 6181 32453 6193 32456
rect 6227 32453 6239 32487
rect 6181 32447 6239 32453
rect 7466 32376 7472 32428
rect 7524 32416 7530 32428
rect 7653 32419 7711 32425
rect 7653 32416 7665 32419
rect 7524 32388 7665 32416
rect 7524 32376 7530 32388
rect 7653 32385 7665 32388
rect 7699 32385 7711 32419
rect 7653 32379 7711 32385
rect 8018 32376 8024 32428
rect 8076 32416 8082 32428
rect 9217 32419 9275 32425
rect 9217 32416 9229 32419
rect 8076 32388 9229 32416
rect 8076 32376 8082 32388
rect 9217 32385 9229 32388
rect 9263 32385 9275 32419
rect 9217 32379 9275 32385
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32416 9551 32419
rect 9674 32416 9680 32428
rect 9539 32388 9680 32416
rect 9539 32385 9551 32388
rect 9493 32379 9551 32385
rect 9674 32376 9680 32388
rect 9732 32376 9738 32428
rect 9950 32376 9956 32428
rect 10008 32416 10014 32428
rect 10318 32416 10324 32428
rect 10008 32388 10324 32416
rect 10008 32376 10014 32388
rect 10318 32376 10324 32388
rect 10376 32416 10382 32428
rect 10597 32419 10655 32425
rect 10597 32416 10609 32419
rect 10376 32388 10609 32416
rect 10376 32376 10382 32388
rect 10597 32385 10609 32388
rect 10643 32385 10655 32419
rect 10597 32379 10655 32385
rect 12526 32376 12532 32428
rect 12584 32416 12590 32428
rect 13538 32416 13544 32428
rect 12584 32388 13544 32416
rect 12584 32376 12590 32388
rect 13538 32376 13544 32388
rect 13596 32416 13602 32428
rect 13633 32419 13691 32425
rect 13633 32416 13645 32419
rect 13596 32388 13645 32416
rect 13596 32376 13602 32388
rect 13633 32385 13645 32388
rect 13679 32385 13691 32419
rect 13633 32379 13691 32385
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32416 13967 32419
rect 15378 32416 15384 32428
rect 13955 32388 15384 32416
rect 13955 32385 13967 32388
rect 13909 32379 13967 32385
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 1489 32351 1547 32357
rect 1489 32317 1501 32351
rect 1535 32317 1547 32351
rect 1489 32311 1547 32317
rect 2869 32351 2927 32357
rect 2869 32317 2881 32351
rect 2915 32317 2927 32351
rect 3050 32348 3056 32360
rect 3011 32320 3056 32348
rect 2869 32311 2927 32317
rect 1578 32212 1584 32224
rect 1539 32184 1584 32212
rect 1578 32172 1584 32184
rect 1636 32172 1642 32224
rect 2884 32212 2912 32311
rect 3050 32308 3056 32320
rect 3108 32308 3114 32360
rect 3605 32351 3663 32357
rect 3605 32317 3617 32351
rect 3651 32317 3663 32351
rect 3786 32348 3792 32360
rect 3699 32320 3792 32348
rect 3605 32311 3663 32317
rect 3068 32280 3096 32308
rect 3620 32280 3648 32311
rect 3786 32308 3792 32320
rect 3844 32348 3850 32360
rect 4062 32348 4068 32360
rect 3844 32320 4068 32348
rect 3844 32308 3850 32320
rect 4062 32308 4068 32320
rect 4120 32308 4126 32360
rect 4798 32308 4804 32360
rect 4856 32348 4862 32360
rect 5077 32351 5135 32357
rect 5077 32348 5089 32351
rect 4856 32320 5089 32348
rect 4856 32308 4862 32320
rect 5077 32317 5089 32320
rect 5123 32317 5135 32351
rect 5077 32311 5135 32317
rect 5718 32308 5724 32360
rect 5776 32348 5782 32360
rect 6365 32351 6423 32357
rect 6365 32348 6377 32351
rect 5776 32320 6377 32348
rect 5776 32308 5782 32320
rect 6365 32317 6377 32320
rect 6411 32348 6423 32351
rect 6454 32348 6460 32360
rect 6411 32320 6460 32348
rect 6411 32317 6423 32320
rect 6365 32311 6423 32317
rect 6454 32308 6460 32320
rect 6512 32308 6518 32360
rect 7837 32351 7895 32357
rect 7837 32317 7849 32351
rect 7883 32317 7895 32351
rect 7837 32311 7895 32317
rect 3068 32252 3648 32280
rect 7098 32240 7104 32292
rect 7156 32280 7162 32292
rect 7852 32280 7880 32311
rect 8110 32308 8116 32360
rect 8168 32348 8174 32360
rect 8205 32351 8263 32357
rect 8205 32348 8217 32351
rect 8168 32320 8217 32348
rect 8168 32308 8174 32320
rect 8205 32317 8217 32320
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 8389 32351 8447 32357
rect 8389 32317 8401 32351
rect 8435 32348 8447 32351
rect 10134 32348 10140 32360
rect 8435 32320 10140 32348
rect 8435 32317 8447 32320
rect 8389 32311 8447 32317
rect 10134 32308 10140 32320
rect 10192 32308 10198 32360
rect 10410 32308 10416 32360
rect 10468 32348 10474 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 10468 32320 12449 32348
rect 10468 32308 10474 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 16298 32348 16304 32360
rect 16259 32320 16304 32348
rect 12437 32311 12495 32317
rect 16298 32308 16304 32320
rect 16356 32308 16362 32360
rect 7156 32252 7880 32280
rect 7156 32240 7162 32252
rect 7926 32240 7932 32292
rect 7984 32280 7990 32292
rect 16117 32283 16175 32289
rect 7984 32252 9352 32280
rect 7984 32240 7990 32252
rect 4706 32212 4712 32224
rect 2884 32184 4712 32212
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 5258 32212 5264 32224
rect 5219 32184 5264 32212
rect 5258 32172 5264 32184
rect 5316 32172 5322 32224
rect 7469 32215 7527 32221
rect 7469 32181 7481 32215
rect 7515 32212 7527 32215
rect 9214 32212 9220 32224
rect 7515 32184 9220 32212
rect 7515 32181 7527 32184
rect 7469 32175 7527 32181
rect 9214 32172 9220 32184
rect 9272 32172 9278 32224
rect 9324 32212 9352 32252
rect 16117 32249 16129 32283
rect 16163 32280 16175 32283
rect 16206 32280 16212 32292
rect 16163 32252 16212 32280
rect 16163 32249 16175 32252
rect 16117 32243 16175 32249
rect 16206 32240 16212 32252
rect 16264 32240 16270 32292
rect 16482 32240 16488 32292
rect 16540 32280 16546 32292
rect 16669 32283 16727 32289
rect 16669 32280 16681 32283
rect 16540 32252 16681 32280
rect 16540 32240 16546 32252
rect 16669 32249 16681 32252
rect 16715 32249 16727 32283
rect 16669 32243 16727 32249
rect 10594 32212 10600 32224
rect 9324 32184 10600 32212
rect 10594 32172 10600 32184
rect 10652 32172 10658 32224
rect 11698 32172 11704 32224
rect 11756 32212 11762 32224
rect 12621 32215 12679 32221
rect 12621 32212 12633 32215
rect 11756 32184 12633 32212
rect 11756 32172 11762 32184
rect 12621 32181 12633 32184
rect 12667 32181 12679 32215
rect 12621 32175 12679 32181
rect 14182 32172 14188 32224
rect 14240 32212 14246 32224
rect 15197 32215 15255 32221
rect 15197 32212 15209 32215
rect 14240 32184 15209 32212
rect 14240 32172 14246 32184
rect 15197 32181 15209 32184
rect 15243 32212 15255 32215
rect 16574 32212 16580 32224
rect 15243 32184 16580 32212
rect 15243 32181 15255 32184
rect 15197 32175 15255 32181
rect 16574 32172 16580 32184
rect 16632 32172 16638 32224
rect 1104 32122 24840 32144
rect 1104 32070 8912 32122
rect 8964 32070 8976 32122
rect 9028 32070 9040 32122
rect 9092 32070 9104 32122
rect 9156 32070 16843 32122
rect 16895 32070 16907 32122
rect 16959 32070 16971 32122
rect 17023 32070 17035 32122
rect 17087 32070 24840 32122
rect 1104 32048 24840 32070
rect 4985 32011 5043 32017
rect 4985 31977 4997 32011
rect 5031 32008 5043 32011
rect 5718 32008 5724 32020
rect 5031 31980 5724 32008
rect 5031 31977 5043 31980
rect 4985 31971 5043 31977
rect 5718 31968 5724 31980
rect 5776 31968 5782 32020
rect 7285 32011 7343 32017
rect 7285 32008 7297 32011
rect 6012 31980 7297 32008
rect 2774 31900 2780 31952
rect 2832 31940 2838 31952
rect 3053 31943 3111 31949
rect 3053 31940 3065 31943
rect 2832 31912 3065 31940
rect 2832 31900 2838 31912
rect 3053 31909 3065 31912
rect 3099 31909 3111 31943
rect 6012 31940 6040 31980
rect 7285 31977 7297 31980
rect 7331 32008 7343 32011
rect 7926 32008 7932 32020
rect 7331 31980 7932 32008
rect 7331 31977 7343 31980
rect 7285 31971 7343 31977
rect 7926 31968 7932 31980
rect 7984 31968 7990 32020
rect 8665 32011 8723 32017
rect 8665 31977 8677 32011
rect 8711 32008 8723 32011
rect 10042 32008 10048 32020
rect 8711 31980 10048 32008
rect 8711 31977 8723 31980
rect 8665 31971 8723 31977
rect 10042 31968 10048 31980
rect 10100 31968 10106 32020
rect 10962 31968 10968 32020
rect 11020 31968 11026 32020
rect 13357 32011 13415 32017
rect 13357 31977 13369 32011
rect 13403 32008 13415 32011
rect 15286 32008 15292 32020
rect 13403 31980 15292 32008
rect 13403 31977 13415 31980
rect 13357 31971 13415 31977
rect 15286 31968 15292 31980
rect 15344 31968 15350 32020
rect 16022 31968 16028 32020
rect 16080 32008 16086 32020
rect 16298 32008 16304 32020
rect 16080 31980 16304 32008
rect 16080 31968 16086 31980
rect 16298 31968 16304 31980
rect 16356 32008 16362 32020
rect 16669 32011 16727 32017
rect 16669 32008 16681 32011
rect 16356 31980 16681 32008
rect 16356 31968 16362 31980
rect 16669 31977 16681 31980
rect 16715 31977 16727 32011
rect 16669 31971 16727 31977
rect 3053 31903 3111 31909
rect 5736 31912 6040 31940
rect 1949 31875 2007 31881
rect 1949 31841 1961 31875
rect 1995 31872 2007 31875
rect 1995 31844 2912 31872
rect 1995 31841 2007 31844
rect 1949 31835 2007 31841
rect 2884 31736 2912 31844
rect 2958 31832 2964 31884
rect 3016 31872 3022 31884
rect 4798 31872 4804 31884
rect 3016 31844 3061 31872
rect 4759 31844 4804 31872
rect 3016 31832 3022 31844
rect 4798 31832 4804 31844
rect 4856 31832 4862 31884
rect 5736 31804 5764 31912
rect 7374 31900 7380 31952
rect 7432 31940 7438 31952
rect 9677 31943 9735 31949
rect 9677 31940 9689 31943
rect 7432 31912 9689 31940
rect 7432 31900 7438 31912
rect 9677 31909 9689 31912
rect 9723 31909 9735 31943
rect 10980 31940 11008 31968
rect 13446 31940 13452 31952
rect 9677 31903 9735 31909
rect 9876 31912 13452 31940
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 5905 31875 5963 31881
rect 5905 31872 5917 31875
rect 5868 31844 5917 31872
rect 5868 31832 5874 31844
rect 5905 31841 5917 31844
rect 5951 31872 5963 31875
rect 6270 31872 6276 31884
rect 5951 31844 6276 31872
rect 5951 31841 5963 31844
rect 5905 31835 5963 31841
rect 6270 31832 6276 31844
rect 6328 31832 6334 31884
rect 8294 31832 8300 31884
rect 8352 31872 8358 31884
rect 9876 31881 9904 31912
rect 13446 31900 13452 31912
rect 13504 31900 13510 31952
rect 8481 31875 8539 31881
rect 8481 31872 8493 31875
rect 8352 31844 8493 31872
rect 8352 31832 8358 31844
rect 8481 31841 8493 31844
rect 8527 31841 8539 31875
rect 8481 31835 8539 31841
rect 9861 31875 9919 31881
rect 9861 31841 9873 31875
rect 9907 31841 9919 31875
rect 11330 31872 11336 31884
rect 11291 31844 11336 31872
rect 9861 31835 9919 31841
rect 6178 31804 6184 31816
rect 4448 31776 5764 31804
rect 6139 31776 6184 31804
rect 4448 31736 4476 31776
rect 6178 31764 6184 31776
rect 6236 31764 6242 31816
rect 8496 31804 8524 31835
rect 11330 31832 11336 31844
rect 11388 31872 11394 31884
rect 11698 31872 11704 31884
rect 11388 31844 11704 31872
rect 11388 31832 11394 31844
rect 11698 31832 11704 31844
rect 11756 31872 11762 31884
rect 11885 31875 11943 31881
rect 11885 31872 11897 31875
rect 11756 31844 11897 31872
rect 11756 31832 11762 31844
rect 11885 31841 11897 31844
rect 11931 31841 11943 31875
rect 12066 31872 12072 31884
rect 12027 31844 12072 31872
rect 11885 31835 11943 31841
rect 12066 31832 12072 31844
rect 12124 31832 12130 31884
rect 12526 31832 12532 31884
rect 12584 31872 12590 31884
rect 13354 31872 13360 31884
rect 12584 31844 13360 31872
rect 12584 31832 12590 31844
rect 13354 31832 13360 31844
rect 13412 31872 13418 31884
rect 13541 31875 13599 31881
rect 13541 31872 13553 31875
rect 13412 31844 13553 31872
rect 13412 31832 13418 31844
rect 13541 31841 13553 31844
rect 13587 31841 13599 31875
rect 13541 31835 13599 31841
rect 13630 31832 13636 31884
rect 13688 31872 13694 31884
rect 14369 31875 14427 31881
rect 13688 31844 13733 31872
rect 13688 31832 13694 31844
rect 14369 31841 14381 31875
rect 14415 31872 14427 31875
rect 14918 31872 14924 31884
rect 14415 31844 14924 31872
rect 14415 31841 14427 31844
rect 14369 31835 14427 31841
rect 14918 31832 14924 31844
rect 14976 31872 14982 31884
rect 16206 31872 16212 31884
rect 14976 31844 16212 31872
rect 14976 31832 14982 31844
rect 16206 31832 16212 31844
rect 16264 31832 16270 31884
rect 16298 31832 16304 31884
rect 16356 31872 16362 31884
rect 16482 31872 16488 31884
rect 16356 31844 16488 31872
rect 16356 31832 16362 31844
rect 16482 31832 16488 31844
rect 16540 31872 16546 31884
rect 17773 31875 17831 31881
rect 17773 31872 17785 31875
rect 16540 31844 17785 31872
rect 16540 31832 16546 31844
rect 17773 31841 17785 31844
rect 17819 31841 17831 31875
rect 17773 31835 17831 31841
rect 8496 31776 8708 31804
rect 2884 31708 4476 31736
rect 4522 31696 4528 31748
rect 4580 31736 4586 31748
rect 5442 31736 5448 31748
rect 4580 31708 5448 31736
rect 4580 31696 4586 31708
rect 5442 31696 5448 31708
rect 5500 31696 5506 31748
rect 8680 31736 8708 31776
rect 8754 31764 8760 31816
rect 8812 31804 8818 31816
rect 10137 31807 10195 31813
rect 10137 31804 10149 31807
rect 8812 31776 10149 31804
rect 8812 31764 8818 31776
rect 10137 31773 10149 31776
rect 10183 31773 10195 31807
rect 10318 31804 10324 31816
rect 10137 31767 10195 31773
rect 10244 31776 10324 31804
rect 9490 31736 9496 31748
rect 8680 31708 9496 31736
rect 9490 31696 9496 31708
rect 9548 31696 9554 31748
rect 10244 31680 10272 31776
rect 10318 31764 10324 31776
rect 10376 31764 10382 31816
rect 11149 31807 11207 31813
rect 11149 31773 11161 31807
rect 11195 31773 11207 31807
rect 11149 31767 11207 31773
rect 14001 31807 14059 31813
rect 14001 31773 14013 31807
rect 14047 31804 14059 31807
rect 14182 31804 14188 31816
rect 14047 31776 14188 31804
rect 14047 31773 14059 31776
rect 14001 31767 14059 31773
rect 11054 31696 11060 31748
rect 11112 31736 11118 31748
rect 11164 31736 11192 31767
rect 14182 31764 14188 31776
rect 14240 31764 14246 31816
rect 15286 31804 15292 31816
rect 15247 31776 15292 31804
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 15562 31804 15568 31816
rect 15523 31776 15568 31804
rect 15562 31764 15568 31776
rect 15620 31764 15626 31816
rect 13814 31745 13820 31748
rect 11112 31708 11192 31736
rect 13798 31739 13820 31745
rect 11112 31696 11118 31708
rect 13798 31705 13810 31739
rect 13798 31699 13820 31705
rect 13814 31696 13820 31699
rect 13872 31696 13878 31748
rect 13906 31696 13912 31748
rect 13964 31736 13970 31748
rect 13964 31708 14009 31736
rect 13964 31696 13970 31708
rect 2041 31671 2099 31677
rect 2041 31637 2053 31671
rect 2087 31668 2099 31671
rect 5350 31668 5356 31680
rect 2087 31640 5356 31668
rect 2087 31637 2099 31640
rect 2041 31631 2099 31637
rect 5350 31628 5356 31640
rect 5408 31628 5414 31680
rect 5810 31628 5816 31680
rect 5868 31668 5874 31680
rect 8018 31668 8024 31680
rect 5868 31640 8024 31668
rect 5868 31628 5874 31640
rect 8018 31628 8024 31640
rect 8076 31628 8082 31680
rect 10226 31628 10232 31680
rect 10284 31628 10290 31680
rect 12342 31668 12348 31680
rect 12303 31640 12348 31668
rect 12342 31628 12348 31640
rect 12400 31628 12406 31680
rect 17862 31668 17868 31680
rect 17823 31640 17868 31668
rect 17862 31628 17868 31640
rect 17920 31628 17926 31680
rect 1104 31578 24840 31600
rect 1104 31526 4947 31578
rect 4999 31526 5011 31578
rect 5063 31526 5075 31578
rect 5127 31526 5139 31578
rect 5191 31526 12878 31578
rect 12930 31526 12942 31578
rect 12994 31526 13006 31578
rect 13058 31526 13070 31578
rect 13122 31526 20808 31578
rect 20860 31526 20872 31578
rect 20924 31526 20936 31578
rect 20988 31526 21000 31578
rect 21052 31526 24840 31578
rect 1104 31504 24840 31526
rect 4430 31424 4436 31476
rect 4488 31424 4494 31476
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 10410 31464 10416 31476
rect 9732 31436 10416 31464
rect 9732 31424 9738 31436
rect 10410 31424 10416 31436
rect 10468 31424 10474 31476
rect 11977 31467 12035 31473
rect 11977 31433 11989 31467
rect 12023 31464 12035 31467
rect 13538 31464 13544 31476
rect 12023 31436 13544 31464
rect 12023 31433 12035 31436
rect 11977 31427 12035 31433
rect 4448 31396 4476 31424
rect 5166 31396 5172 31408
rect 4080 31368 5172 31396
rect 1486 31328 1492 31340
rect 1447 31300 1492 31328
rect 1486 31288 1492 31300
rect 1544 31288 1550 31340
rect 4080 31337 4108 31368
rect 5166 31356 5172 31368
rect 5224 31356 5230 31408
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 4065 31331 4123 31337
rect 1811 31300 3004 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 1762 31084 1768 31136
rect 1820 31124 1826 31136
rect 2869 31127 2927 31133
rect 2869 31124 2881 31127
rect 1820 31096 2881 31124
rect 1820 31084 1826 31096
rect 2869 31093 2881 31096
rect 2915 31093 2927 31127
rect 2976 31124 3004 31300
rect 4065 31297 4077 31331
rect 4111 31297 4123 31331
rect 9677 31331 9735 31337
rect 9677 31328 9689 31331
rect 4065 31291 4123 31297
rect 7116 31300 9689 31328
rect 3050 31220 3056 31272
rect 3108 31260 3114 31272
rect 4157 31263 4215 31269
rect 4157 31260 4169 31263
rect 3108 31232 4169 31260
rect 3108 31220 3114 31232
rect 4157 31229 4169 31232
rect 4203 31229 4215 31263
rect 4157 31223 4215 31229
rect 4709 31263 4767 31269
rect 4709 31229 4721 31263
rect 4755 31229 4767 31263
rect 4890 31260 4896 31272
rect 4851 31232 4896 31260
rect 4709 31223 4767 31229
rect 4172 31192 4200 31223
rect 4724 31192 4752 31223
rect 4890 31220 4896 31232
rect 4948 31220 4954 31272
rect 7116 31269 7144 31300
rect 9677 31297 9689 31300
rect 9723 31328 9735 31331
rect 9766 31328 9772 31340
rect 9723 31300 9772 31328
rect 9723 31297 9735 31300
rect 9677 31291 9735 31297
rect 9766 31288 9772 31300
rect 9824 31288 9830 31340
rect 10318 31288 10324 31340
rect 10376 31328 10382 31340
rect 10376 31300 10824 31328
rect 10376 31288 10382 31300
rect 7101 31263 7159 31269
rect 7101 31229 7113 31263
rect 7147 31229 7159 31263
rect 7101 31223 7159 31229
rect 8018 31220 8024 31272
rect 8076 31260 8082 31272
rect 8113 31263 8171 31269
rect 8113 31260 8125 31263
rect 8076 31232 8125 31260
rect 8076 31220 8082 31232
rect 8113 31229 8125 31232
rect 8159 31229 8171 31263
rect 8113 31223 8171 31229
rect 8389 31263 8447 31269
rect 8389 31229 8401 31263
rect 8435 31260 8447 31263
rect 10410 31260 10416 31272
rect 8435 31232 10416 31260
rect 8435 31229 8447 31232
rect 8389 31223 8447 31229
rect 10410 31220 10416 31232
rect 10468 31220 10474 31272
rect 10594 31260 10600 31272
rect 10555 31232 10600 31260
rect 10594 31220 10600 31232
rect 10652 31220 10658 31272
rect 10796 31269 10824 31300
rect 10781 31263 10839 31269
rect 10781 31229 10793 31263
rect 10827 31260 10839 31263
rect 12161 31263 12219 31269
rect 10827 31232 11008 31260
rect 10827 31229 10839 31232
rect 10781 31223 10839 31229
rect 4172 31164 4752 31192
rect 9214 31152 9220 31204
rect 9272 31192 9278 31204
rect 9272 31164 10916 31192
rect 9272 31152 9278 31164
rect 5169 31127 5227 31133
rect 5169 31124 5181 31127
rect 2976 31096 5181 31124
rect 2869 31087 2927 31093
rect 5169 31093 5181 31096
rect 5215 31093 5227 31127
rect 5169 31087 5227 31093
rect 7193 31127 7251 31133
rect 7193 31093 7205 31127
rect 7239 31124 7251 31127
rect 9398 31124 9404 31136
rect 7239 31096 9404 31124
rect 7239 31093 7251 31096
rect 7193 31087 7251 31093
rect 9398 31084 9404 31096
rect 9456 31084 9462 31136
rect 10888 31133 10916 31164
rect 10873 31127 10931 31133
rect 10873 31093 10885 31127
rect 10919 31093 10931 31127
rect 10980 31124 11008 31232
rect 12161 31229 12173 31263
rect 12207 31229 12219 31263
rect 12268 31260 12296 31436
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 14001 31467 14059 31473
rect 14001 31433 14013 31467
rect 14047 31464 14059 31467
rect 14182 31464 14188 31476
rect 14047 31436 14188 31464
rect 14047 31433 14059 31436
rect 14001 31427 14059 31433
rect 14182 31424 14188 31436
rect 14240 31424 14246 31476
rect 15197 31467 15255 31473
rect 15197 31433 15209 31467
rect 15243 31464 15255 31467
rect 15562 31464 15568 31476
rect 15243 31436 15568 31464
rect 15243 31433 15255 31436
rect 15197 31427 15255 31433
rect 15562 31424 15568 31436
rect 15620 31424 15626 31476
rect 17862 31396 17868 31408
rect 15764 31368 17868 31396
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 12713 31331 12771 31337
rect 12713 31328 12725 31331
rect 12400 31300 12725 31328
rect 12400 31288 12406 31300
rect 12713 31297 12725 31300
rect 12759 31297 12771 31331
rect 12713 31291 12771 31297
rect 12434 31260 12440 31272
rect 12268 31232 12440 31260
rect 12161 31223 12219 31229
rect 12176 31192 12204 31223
rect 12434 31220 12440 31232
rect 12492 31260 12498 31272
rect 15764 31269 15792 31368
rect 17862 31356 17868 31368
rect 17920 31356 17926 31408
rect 16206 31328 16212 31340
rect 16167 31300 16212 31328
rect 16206 31288 16212 31300
rect 16264 31288 16270 31340
rect 15749 31263 15807 31269
rect 12492 31232 12585 31260
rect 12492 31220 12498 31232
rect 15749 31229 15761 31263
rect 15795 31229 15807 31263
rect 15749 31223 15807 31229
rect 15838 31220 15844 31272
rect 15896 31260 15902 31272
rect 16117 31263 16175 31269
rect 15896 31232 15941 31260
rect 15896 31220 15902 31232
rect 16117 31229 16129 31263
rect 16163 31229 16175 31263
rect 16117 31223 16175 31229
rect 12526 31192 12532 31204
rect 12176 31164 12532 31192
rect 12526 31152 12532 31164
rect 12584 31152 12590 31204
rect 15378 31152 15384 31204
rect 15436 31192 15442 31204
rect 16022 31192 16028 31204
rect 15436 31164 16028 31192
rect 15436 31152 15442 31164
rect 16022 31152 16028 31164
rect 16080 31192 16086 31204
rect 16132 31192 16160 31223
rect 16080 31164 16160 31192
rect 16080 31152 16086 31164
rect 13906 31124 13912 31136
rect 10980 31096 13912 31124
rect 10873 31087 10931 31093
rect 13906 31084 13912 31096
rect 13964 31084 13970 31136
rect 1104 31034 24840 31056
rect 1104 30982 8912 31034
rect 8964 30982 8976 31034
rect 9028 30982 9040 31034
rect 9092 30982 9104 31034
rect 9156 30982 16843 31034
rect 16895 30982 16907 31034
rect 16959 30982 16971 31034
rect 17023 30982 17035 31034
rect 17087 30982 24840 31034
rect 1104 30960 24840 30982
rect 3050 30920 3056 30932
rect 3011 30892 3056 30920
rect 3050 30880 3056 30892
rect 3108 30880 3114 30932
rect 3602 30880 3608 30932
rect 3660 30920 3666 30932
rect 4798 30920 4804 30932
rect 3660 30892 4804 30920
rect 3660 30880 3666 30892
rect 4798 30880 4804 30892
rect 4856 30880 4862 30932
rect 6178 30920 6184 30932
rect 6139 30892 6184 30920
rect 6178 30880 6184 30892
rect 6236 30880 6242 30932
rect 10318 30920 10324 30932
rect 7668 30892 10324 30920
rect 5810 30852 5816 30864
rect 1872 30824 5816 30852
rect 1872 30793 1900 30824
rect 5810 30812 5816 30824
rect 5868 30812 5874 30864
rect 7190 30812 7196 30864
rect 7248 30852 7254 30864
rect 7469 30855 7527 30861
rect 7469 30852 7481 30855
rect 7248 30824 7481 30852
rect 7248 30812 7254 30824
rect 7469 30821 7481 30824
rect 7515 30821 7527 30855
rect 7469 30815 7527 30821
rect 1849 30787 1907 30793
rect 1849 30753 1861 30787
rect 1895 30753 1907 30787
rect 1849 30747 1907 30753
rect 2869 30787 2927 30793
rect 2869 30753 2881 30787
rect 2915 30784 2927 30787
rect 2958 30784 2964 30796
rect 2915 30756 2964 30784
rect 2915 30753 2927 30756
rect 2869 30747 2927 30753
rect 2958 30744 2964 30756
rect 3016 30744 3022 30796
rect 5169 30787 5227 30793
rect 5169 30753 5181 30787
rect 5215 30784 5227 30787
rect 5258 30784 5264 30796
rect 5215 30756 5264 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 5258 30744 5264 30756
rect 5316 30744 5322 30796
rect 5350 30744 5356 30796
rect 5408 30784 5414 30796
rect 5629 30787 5687 30793
rect 5629 30784 5641 30787
rect 5408 30756 5641 30784
rect 5408 30744 5414 30756
rect 5629 30753 5641 30756
rect 5675 30753 5687 30787
rect 5629 30747 5687 30753
rect 5718 30744 5724 30796
rect 5776 30784 5782 30796
rect 5776 30756 6408 30784
rect 5776 30744 5782 30756
rect 4430 30676 4436 30728
rect 4488 30716 4494 30728
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4488 30688 4997 30716
rect 4488 30676 4494 30688
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 6380 30716 6408 30756
rect 6454 30744 6460 30796
rect 6512 30784 6518 30796
rect 7668 30793 7696 30892
rect 10318 30880 10324 30892
rect 10376 30880 10382 30932
rect 10410 30880 10416 30932
rect 10468 30920 10474 30932
rect 10965 30923 11023 30929
rect 10965 30920 10977 30923
rect 10468 30892 10977 30920
rect 10468 30880 10474 30892
rect 10965 30889 10977 30892
rect 11011 30889 11023 30923
rect 10965 30883 11023 30889
rect 11422 30880 11428 30932
rect 11480 30920 11486 30932
rect 11480 30892 13032 30920
rect 11480 30880 11486 30892
rect 9398 30812 9404 30864
rect 9456 30852 9462 30864
rect 9456 30824 10732 30852
rect 9456 30812 9462 30824
rect 7377 30787 7435 30793
rect 7377 30784 7389 30787
rect 6512 30756 7389 30784
rect 6512 30744 6518 30756
rect 7377 30753 7389 30756
rect 7423 30753 7435 30787
rect 7377 30747 7435 30753
rect 7653 30787 7711 30793
rect 7653 30753 7665 30787
rect 7699 30753 7711 30787
rect 9950 30784 9956 30796
rect 9911 30756 9956 30784
rect 7653 30747 7711 30753
rect 9950 30744 9956 30756
rect 10008 30784 10014 30796
rect 10318 30784 10324 30796
rect 10008 30756 10324 30784
rect 10008 30744 10014 30756
rect 10318 30744 10324 30756
rect 10376 30784 10382 30796
rect 10704 30793 10732 30824
rect 11790 30812 11796 30864
rect 11848 30852 11854 30864
rect 11977 30855 12035 30861
rect 11977 30852 11989 30855
rect 11848 30824 11989 30852
rect 11848 30812 11854 30824
rect 11977 30821 11989 30824
rect 12023 30821 12035 30855
rect 11977 30815 12035 30821
rect 12158 30812 12164 30864
rect 12216 30852 12222 30864
rect 12216 30824 12664 30852
rect 12216 30812 12222 30824
rect 12636 30793 12664 30824
rect 13004 30793 13032 30892
rect 14458 30880 14464 30932
rect 14516 30920 14522 30932
rect 14642 30920 14648 30932
rect 14516 30892 14648 30920
rect 14516 30880 14522 30892
rect 14642 30880 14648 30892
rect 14700 30880 14706 30932
rect 15194 30880 15200 30932
rect 15252 30920 15258 30932
rect 15933 30923 15991 30929
rect 15933 30920 15945 30923
rect 15252 30892 15945 30920
rect 15252 30880 15258 30892
rect 15933 30889 15945 30892
rect 15979 30889 15991 30923
rect 15933 30883 15991 30889
rect 10505 30787 10563 30793
rect 10505 30784 10517 30787
rect 10376 30756 10517 30784
rect 10376 30744 10382 30756
rect 10505 30753 10517 30756
rect 10551 30753 10563 30787
rect 10505 30747 10563 30753
rect 10689 30787 10747 30793
rect 10689 30753 10701 30787
rect 10735 30784 10747 30787
rect 12437 30787 12495 30793
rect 12437 30784 12449 30787
rect 10735 30756 12449 30784
rect 10735 30753 10747 30756
rect 10689 30747 10747 30753
rect 12437 30753 12449 30756
rect 12483 30753 12495 30787
rect 12437 30747 12495 30753
rect 12621 30787 12679 30793
rect 12621 30753 12633 30787
rect 12667 30753 12679 30787
rect 12621 30747 12679 30753
rect 12989 30787 13047 30793
rect 12989 30753 13001 30787
rect 13035 30753 13047 30787
rect 12989 30747 13047 30753
rect 13173 30787 13231 30793
rect 13173 30753 13185 30787
rect 13219 30753 13231 30787
rect 13998 30784 14004 30796
rect 13959 30756 14004 30784
rect 13173 30747 13231 30753
rect 7006 30716 7012 30728
rect 6380 30688 7012 30716
rect 4985 30679 5043 30685
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 9907 30688 9996 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 9968 30660 9996 30688
rect 12066 30676 12072 30728
rect 12124 30716 12130 30728
rect 13188 30716 13216 30747
rect 13998 30744 14004 30756
rect 14056 30744 14062 30796
rect 15013 30787 15071 30793
rect 15013 30753 15025 30787
rect 15059 30784 15071 30787
rect 15289 30787 15347 30793
rect 15289 30784 15301 30787
rect 15059 30756 15301 30784
rect 15059 30753 15071 30756
rect 15013 30747 15071 30753
rect 15289 30753 15301 30756
rect 15335 30753 15347 30787
rect 15289 30747 15347 30753
rect 16574 30744 16580 30796
rect 16632 30784 16638 30796
rect 16853 30787 16911 30793
rect 16853 30784 16865 30787
rect 16632 30756 16865 30784
rect 16632 30744 16638 30756
rect 16853 30753 16865 30756
rect 16899 30753 16911 30787
rect 16853 30747 16911 30753
rect 15657 30719 15715 30725
rect 12124 30688 15332 30716
rect 12124 30676 12130 30688
rect 15304 30660 15332 30688
rect 15657 30685 15669 30719
rect 15703 30716 15715 30719
rect 16022 30716 16028 30728
rect 15703 30688 16028 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 16022 30676 16028 30688
rect 16080 30676 16086 30728
rect 1949 30651 2007 30657
rect 1949 30617 1961 30651
rect 1995 30648 2007 30651
rect 3970 30648 3976 30660
rect 1995 30620 3976 30648
rect 1995 30617 2007 30620
rect 1949 30611 2007 30617
rect 3970 30608 3976 30620
rect 4028 30608 4034 30660
rect 5350 30608 5356 30660
rect 5408 30648 5414 30660
rect 5902 30648 5908 30660
rect 5408 30620 5908 30648
rect 5408 30608 5414 30620
rect 5902 30608 5908 30620
rect 5960 30608 5966 30660
rect 8018 30648 8024 30660
rect 7668 30620 8024 30648
rect 7190 30580 7196 30592
rect 7151 30552 7196 30580
rect 7190 30540 7196 30552
rect 7248 30580 7254 30592
rect 7668 30580 7696 30620
rect 8018 30608 8024 30620
rect 8076 30608 8082 30660
rect 9950 30608 9956 30660
rect 10008 30648 10014 30660
rect 11054 30648 11060 30660
rect 10008 30620 11060 30648
rect 10008 30608 10014 30620
rect 11054 30608 11060 30620
rect 11112 30608 11118 30660
rect 11514 30608 11520 30660
rect 11572 30648 11578 30660
rect 13446 30648 13452 30660
rect 11572 30620 13452 30648
rect 11572 30608 11578 30620
rect 13446 30608 13452 30620
rect 13504 30608 13510 30660
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 16945 30651 17003 30657
rect 16945 30648 16957 30651
rect 15344 30620 16957 30648
rect 15344 30608 15350 30620
rect 16945 30617 16957 30620
rect 16991 30617 17003 30651
rect 16945 30611 17003 30617
rect 7248 30552 7696 30580
rect 7745 30583 7803 30589
rect 7248 30540 7254 30552
rect 7745 30549 7757 30583
rect 7791 30580 7803 30583
rect 7834 30580 7840 30592
rect 7791 30552 7840 30580
rect 7791 30549 7803 30552
rect 7745 30543 7803 30549
rect 7834 30540 7840 30552
rect 7892 30540 7898 30592
rect 14090 30580 14096 30592
rect 14051 30552 14096 30580
rect 14090 30540 14096 30552
rect 14148 30580 14154 30592
rect 15013 30583 15071 30589
rect 15013 30580 15025 30583
rect 14148 30552 15025 30580
rect 14148 30540 14154 30552
rect 15013 30549 15025 30552
rect 15059 30549 15071 30583
rect 15013 30543 15071 30549
rect 15378 30540 15384 30592
rect 15436 30589 15442 30592
rect 15436 30583 15485 30589
rect 15436 30549 15439 30583
rect 15473 30549 15485 30583
rect 15436 30543 15485 30549
rect 15565 30583 15623 30589
rect 15565 30549 15577 30583
rect 15611 30580 15623 30583
rect 16482 30580 16488 30592
rect 15611 30552 16488 30580
rect 15611 30549 15623 30552
rect 15565 30543 15623 30549
rect 15436 30540 15442 30543
rect 16482 30540 16488 30552
rect 16540 30540 16546 30592
rect 1104 30490 24840 30512
rect 1104 30438 4947 30490
rect 4999 30438 5011 30490
rect 5063 30438 5075 30490
rect 5127 30438 5139 30490
rect 5191 30438 12878 30490
rect 12930 30438 12942 30490
rect 12994 30438 13006 30490
rect 13058 30438 13070 30490
rect 13122 30438 20808 30490
rect 20860 30438 20872 30490
rect 20924 30438 20936 30490
rect 20988 30438 21000 30490
rect 21052 30438 24840 30490
rect 1104 30416 24840 30438
rect 3510 30336 3516 30388
rect 3568 30376 3574 30388
rect 5534 30376 5540 30388
rect 3568 30348 5540 30376
rect 3568 30336 3574 30348
rect 5534 30336 5540 30348
rect 5592 30336 5598 30388
rect 2866 30268 2872 30320
rect 2924 30308 2930 30320
rect 10597 30311 10655 30317
rect 2924 30280 4292 30308
rect 2924 30268 2930 30280
rect 1949 30175 2007 30181
rect 1949 30141 1961 30175
rect 1995 30172 2007 30175
rect 2498 30172 2504 30184
rect 1995 30144 2504 30172
rect 1995 30141 2007 30144
rect 1949 30135 2007 30141
rect 2498 30132 2504 30144
rect 2556 30132 2562 30184
rect 3050 30132 3056 30184
rect 3108 30172 3114 30184
rect 3145 30175 3203 30181
rect 3145 30172 3157 30175
rect 3108 30144 3157 30172
rect 3108 30132 3114 30144
rect 3145 30141 3157 30144
rect 3191 30141 3203 30175
rect 3145 30135 3203 30141
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30172 3295 30175
rect 3510 30172 3516 30184
rect 3283 30144 3516 30172
rect 3283 30141 3295 30144
rect 3237 30135 3295 30141
rect 3510 30132 3516 30144
rect 3568 30132 3574 30184
rect 3605 30175 3663 30181
rect 3605 30141 3617 30175
rect 3651 30141 3663 30175
rect 3605 30135 3663 30141
rect 3697 30175 3755 30181
rect 3697 30141 3709 30175
rect 3743 30172 3755 30175
rect 4062 30172 4068 30184
rect 3743 30144 4068 30172
rect 3743 30141 3755 30144
rect 3697 30135 3755 30141
rect 2041 30107 2099 30113
rect 2041 30073 2053 30107
rect 2087 30104 2099 30107
rect 3620 30104 3648 30135
rect 4062 30132 4068 30144
rect 4120 30132 4126 30184
rect 4154 30132 4160 30184
rect 4212 30132 4218 30184
rect 4264 30172 4292 30280
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 11146 30308 11152 30320
rect 10643 30280 11152 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 11146 30268 11152 30280
rect 11204 30268 11210 30320
rect 11790 30268 11796 30320
rect 11848 30308 11854 30320
rect 13998 30308 14004 30320
rect 11848 30280 14004 30308
rect 11848 30268 11854 30280
rect 8754 30240 8760 30252
rect 8128 30212 8760 30240
rect 5353 30175 5411 30181
rect 5353 30172 5365 30175
rect 4264 30144 5365 30172
rect 5353 30141 5365 30144
rect 5399 30141 5411 30175
rect 5353 30135 5411 30141
rect 5537 30175 5595 30181
rect 5537 30141 5549 30175
rect 5583 30172 5595 30175
rect 5583 30144 6408 30172
rect 5583 30141 5595 30144
rect 5537 30135 5595 30141
rect 4172 30104 4200 30132
rect 4338 30104 4344 30116
rect 2087 30076 4344 30104
rect 2087 30073 2099 30076
rect 2041 30067 2099 30073
rect 4338 30064 4344 30076
rect 4396 30064 4402 30116
rect 5368 30104 5396 30135
rect 5718 30104 5724 30116
rect 5368 30076 5724 30104
rect 5718 30064 5724 30076
rect 5776 30064 5782 30116
rect 5902 30104 5908 30116
rect 5863 30076 5908 30104
rect 5902 30064 5908 30076
rect 5960 30064 5966 30116
rect 6380 30104 6408 30144
rect 6454 30132 6460 30184
rect 6512 30172 6518 30184
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 6512 30144 6837 30172
rect 6512 30132 6518 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 8018 30172 8024 30184
rect 7979 30144 8024 30172
rect 6825 30135 6883 30141
rect 8018 30132 8024 30144
rect 8076 30132 8082 30184
rect 8128 30181 8156 30212
rect 8754 30200 8760 30212
rect 8812 30200 8818 30252
rect 12618 30240 12624 30252
rect 12579 30212 12624 30240
rect 12618 30200 12624 30212
rect 12676 30200 12682 30252
rect 8113 30175 8171 30181
rect 8113 30141 8125 30175
rect 8159 30141 8171 30175
rect 8113 30135 8171 30141
rect 8205 30175 8263 30181
rect 8205 30141 8217 30175
rect 8251 30172 8263 30175
rect 9214 30172 9220 30184
rect 8251 30144 9220 30172
rect 8251 30141 8263 30144
rect 8205 30135 8263 30141
rect 9214 30132 9220 30144
rect 9272 30132 9278 30184
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30172 10839 30175
rect 10965 30175 11023 30181
rect 10827 30144 10916 30172
rect 10827 30141 10839 30144
rect 10781 30135 10839 30141
rect 7374 30104 7380 30116
rect 6380 30076 7380 30104
rect 7374 30064 7380 30076
rect 7432 30064 7438 30116
rect 8662 30104 8668 30116
rect 8623 30076 8668 30104
rect 8662 30064 8668 30076
rect 8720 30064 8726 30116
rect 4154 30036 4160 30048
rect 4115 30008 4160 30036
rect 4154 29996 4160 30008
rect 4212 29996 4218 30048
rect 6914 30036 6920 30048
rect 6875 30008 6920 30036
rect 6914 29996 6920 30008
rect 6972 29996 6978 30048
rect 10888 30036 10916 30144
rect 10965 30141 10977 30175
rect 11011 30141 11023 30175
rect 10965 30135 11023 30141
rect 11333 30175 11391 30181
rect 11333 30141 11345 30175
rect 11379 30172 11391 30175
rect 11422 30172 11428 30184
rect 11379 30144 11428 30172
rect 11379 30141 11391 30144
rect 11333 30135 11391 30141
rect 10980 30104 11008 30135
rect 11422 30132 11428 30144
rect 11480 30132 11486 30184
rect 11517 30175 11575 30181
rect 11517 30141 11529 30175
rect 11563 30172 11575 30175
rect 12158 30172 12164 30184
rect 11563 30144 12164 30172
rect 11563 30141 11575 30144
rect 11517 30135 11575 30141
rect 12158 30132 12164 30144
rect 12216 30132 12222 30184
rect 12989 30175 13047 30181
rect 12989 30141 13001 30175
rect 13035 30172 13047 30175
rect 13170 30172 13176 30184
rect 13035 30144 13176 30172
rect 13035 30141 13047 30144
rect 12989 30135 13047 30141
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 13280 30181 13308 30280
rect 13998 30268 14004 30280
rect 14056 30268 14062 30320
rect 13541 30243 13599 30249
rect 13541 30209 13553 30243
rect 13587 30240 13599 30243
rect 13630 30240 13636 30252
rect 13587 30212 13636 30240
rect 13587 30209 13599 30212
rect 13541 30203 13599 30209
rect 13630 30200 13636 30212
rect 13688 30200 13694 30252
rect 15838 30240 15844 30252
rect 15799 30212 15844 30240
rect 15838 30200 15844 30212
rect 15896 30200 15902 30252
rect 16206 30200 16212 30252
rect 16264 30240 16270 30252
rect 16393 30243 16451 30249
rect 16393 30240 16405 30243
rect 16264 30212 16405 30240
rect 16264 30200 16270 30212
rect 16393 30209 16405 30212
rect 16439 30209 16451 30243
rect 16393 30203 16451 30209
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30141 13323 30175
rect 15930 30172 15936 30184
rect 15891 30144 15936 30172
rect 13265 30135 13323 30141
rect 15930 30132 15936 30144
rect 15988 30132 15994 30184
rect 16301 30175 16359 30181
rect 16301 30141 16313 30175
rect 16347 30172 16359 30175
rect 16482 30172 16488 30184
rect 16347 30144 16488 30172
rect 16347 30141 16359 30144
rect 16301 30135 16359 30141
rect 16482 30132 16488 30144
rect 16540 30132 16546 30184
rect 12066 30104 12072 30116
rect 10980 30076 12072 30104
rect 12066 30064 12072 30076
rect 12124 30064 12130 30116
rect 15289 30107 15347 30113
rect 15289 30073 15301 30107
rect 15335 30104 15347 30107
rect 15562 30104 15568 30116
rect 15335 30076 15568 30104
rect 15335 30073 15347 30076
rect 15289 30067 15347 30073
rect 15562 30064 15568 30076
rect 15620 30064 15626 30116
rect 11054 30036 11060 30048
rect 10888 30008 11060 30036
rect 11054 29996 11060 30008
rect 11112 30036 11118 30048
rect 17586 30036 17592 30048
rect 11112 30008 17592 30036
rect 11112 29996 11118 30008
rect 17586 29996 17592 30008
rect 17644 29996 17650 30048
rect 1104 29946 24840 29968
rect 1104 29894 8912 29946
rect 8964 29894 8976 29946
rect 9028 29894 9040 29946
rect 9092 29894 9104 29946
rect 9156 29894 16843 29946
rect 16895 29894 16907 29946
rect 16959 29894 16971 29946
rect 17023 29894 17035 29946
rect 17087 29894 24840 29946
rect 1104 29872 24840 29894
rect 3510 29792 3516 29844
rect 3568 29832 3574 29844
rect 4430 29832 4436 29844
rect 3568 29804 4436 29832
rect 3568 29792 3574 29804
rect 4430 29792 4436 29804
rect 4488 29792 4494 29844
rect 4893 29835 4951 29841
rect 4893 29801 4905 29835
rect 4939 29832 4951 29835
rect 5350 29832 5356 29844
rect 4939 29804 5356 29832
rect 4939 29801 4951 29804
rect 4893 29795 4951 29801
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 5718 29792 5724 29844
rect 5776 29832 5782 29844
rect 7193 29835 7251 29841
rect 7193 29832 7205 29835
rect 5776 29804 7205 29832
rect 5776 29792 5782 29804
rect 7193 29801 7205 29804
rect 7239 29801 7251 29835
rect 11514 29832 11520 29844
rect 7193 29795 7251 29801
rect 9692 29804 11520 29832
rect 3142 29724 3148 29776
rect 3200 29764 3206 29776
rect 3418 29764 3424 29776
rect 3200 29736 3424 29764
rect 3200 29724 3206 29736
rect 3418 29724 3424 29736
rect 3476 29724 3482 29776
rect 8018 29724 8024 29776
rect 8076 29764 8082 29776
rect 9692 29764 9720 29804
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 9858 29764 9864 29776
rect 8076 29736 9720 29764
rect 9819 29736 9864 29764
rect 8076 29724 8082 29736
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 1486 29696 1492 29708
rect 1443 29668 1492 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 1486 29656 1492 29668
rect 1544 29656 1550 29708
rect 1673 29699 1731 29705
rect 1673 29665 1685 29699
rect 1719 29696 1731 29699
rect 4154 29696 4160 29708
rect 1719 29668 4160 29696
rect 1719 29665 1731 29668
rect 1673 29659 1731 29665
rect 4154 29656 4160 29668
rect 4212 29656 4218 29708
rect 4709 29699 4767 29705
rect 4709 29665 4721 29699
rect 4755 29696 4767 29699
rect 5813 29699 5871 29705
rect 4755 29668 5028 29696
rect 4755 29665 4767 29668
rect 4709 29659 4767 29665
rect 3418 29588 3424 29640
rect 3476 29628 3482 29640
rect 3602 29628 3608 29640
rect 3476 29600 3608 29628
rect 3476 29588 3482 29600
rect 3602 29588 3608 29600
rect 3660 29588 3666 29640
rect 2498 29452 2504 29504
rect 2556 29492 2562 29504
rect 2777 29495 2835 29501
rect 2777 29492 2789 29495
rect 2556 29464 2789 29492
rect 2556 29452 2562 29464
rect 2777 29461 2789 29464
rect 2823 29461 2835 29495
rect 5000 29492 5028 29668
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 7190 29696 7196 29708
rect 5859 29668 7196 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 7190 29656 7196 29668
rect 7248 29656 7254 29708
rect 8481 29699 8539 29705
rect 8481 29665 8493 29699
rect 8527 29696 8539 29699
rect 9398 29696 9404 29708
rect 8527 29668 9404 29696
rect 8527 29665 8539 29668
rect 8481 29659 8539 29665
rect 9398 29656 9404 29668
rect 9456 29656 9462 29708
rect 9692 29705 9720 29736
rect 9858 29724 9864 29736
rect 9916 29724 9922 29776
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 9953 29699 10011 29705
rect 9953 29665 9965 29699
rect 9999 29696 10011 29699
rect 11698 29696 11704 29708
rect 9999 29668 10088 29696
rect 11659 29668 11704 29696
rect 9999 29665 10011 29668
rect 9953 29659 10011 29665
rect 6089 29631 6147 29637
rect 6089 29597 6101 29631
rect 6135 29628 6147 29631
rect 8018 29628 8024 29640
rect 6135 29600 8024 29628
rect 6135 29597 6147 29600
rect 6089 29591 6147 29597
rect 8018 29588 8024 29600
rect 8076 29588 8082 29640
rect 10060 29560 10088 29668
rect 11698 29656 11704 29668
rect 11756 29656 11762 29708
rect 12158 29696 12164 29708
rect 12119 29668 12164 29696
rect 12158 29656 12164 29668
rect 12216 29656 12222 29708
rect 12253 29699 12311 29705
rect 12253 29665 12265 29699
rect 12299 29696 12311 29699
rect 12618 29696 12624 29708
rect 12299 29668 12624 29696
rect 12299 29665 12311 29668
rect 12253 29659 12311 29665
rect 12618 29656 12624 29668
rect 12676 29656 12682 29708
rect 13722 29696 13728 29708
rect 13683 29668 13728 29696
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 13906 29696 13912 29708
rect 13867 29668 13912 29696
rect 13906 29656 13912 29668
rect 13964 29656 13970 29708
rect 15194 29656 15200 29708
rect 15252 29696 15258 29708
rect 15289 29699 15347 29705
rect 15289 29696 15301 29699
rect 15252 29668 15301 29696
rect 15252 29656 15258 29668
rect 15289 29665 15301 29668
rect 15335 29665 15347 29699
rect 15562 29696 15568 29708
rect 15523 29668 15568 29696
rect 15289 29659 15347 29665
rect 15562 29656 15568 29668
rect 15620 29656 15626 29708
rect 10134 29588 10140 29640
rect 10192 29628 10198 29640
rect 11517 29631 11575 29637
rect 11517 29628 11529 29631
rect 10192 29600 11529 29628
rect 10192 29588 10198 29600
rect 11517 29597 11529 29600
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 10060 29532 14044 29560
rect 6178 29492 6184 29504
rect 5000 29464 6184 29492
rect 2777 29455 2835 29461
rect 6178 29452 6184 29464
rect 6236 29452 6242 29504
rect 8570 29452 8576 29504
rect 8628 29492 8634 29504
rect 8665 29495 8723 29501
rect 8665 29492 8677 29495
rect 8628 29464 8677 29492
rect 8628 29452 8634 29464
rect 8665 29461 8677 29464
rect 8711 29461 8723 29495
rect 8665 29455 8723 29461
rect 9766 29452 9772 29504
rect 9824 29492 9830 29504
rect 10137 29495 10195 29501
rect 10137 29492 10149 29495
rect 9824 29464 10149 29492
rect 9824 29452 9830 29464
rect 10137 29461 10149 29464
rect 10183 29461 10195 29495
rect 12710 29492 12716 29504
rect 12671 29464 12716 29492
rect 10137 29455 10195 29461
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 14016 29501 14044 29532
rect 14001 29495 14059 29501
rect 14001 29461 14013 29495
rect 14047 29461 14059 29495
rect 14001 29455 14059 29461
rect 16482 29452 16488 29504
rect 16540 29492 16546 29504
rect 16669 29495 16727 29501
rect 16669 29492 16681 29495
rect 16540 29464 16681 29492
rect 16540 29452 16546 29464
rect 16669 29461 16681 29464
rect 16715 29461 16727 29495
rect 16669 29455 16727 29461
rect 1104 29402 24840 29424
rect 1104 29350 4947 29402
rect 4999 29350 5011 29402
rect 5063 29350 5075 29402
rect 5127 29350 5139 29402
rect 5191 29350 12878 29402
rect 12930 29350 12942 29402
rect 12994 29350 13006 29402
rect 13058 29350 13070 29402
rect 13122 29350 20808 29402
rect 20860 29350 20872 29402
rect 20924 29350 20936 29402
rect 20988 29350 21000 29402
rect 21052 29350 24840 29402
rect 1104 29328 24840 29350
rect 8018 29288 8024 29300
rect 7979 29260 8024 29288
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 15362 29291 15420 29297
rect 15362 29288 15374 29291
rect 12216 29260 15374 29288
rect 12216 29248 12222 29260
rect 15362 29257 15374 29260
rect 15408 29288 15420 29291
rect 18141 29291 18199 29297
rect 18141 29288 18153 29291
rect 15408 29260 18153 29288
rect 15408 29257 15420 29260
rect 15362 29251 15420 29257
rect 18141 29257 18153 29260
rect 18187 29257 18199 29291
rect 18141 29251 18199 29257
rect 4985 29223 5043 29229
rect 4985 29220 4997 29223
rect 2700 29192 4997 29220
rect 1397 29087 1455 29093
rect 1397 29053 1409 29087
rect 1443 29084 1455 29087
rect 1486 29084 1492 29096
rect 1443 29056 1492 29084
rect 1443 29053 1455 29056
rect 1397 29047 1455 29053
rect 1486 29044 1492 29056
rect 1544 29044 1550 29096
rect 1673 29087 1731 29093
rect 1673 29053 1685 29087
rect 1719 29084 1731 29087
rect 2700 29084 2728 29192
rect 4985 29189 4997 29192
rect 5031 29189 5043 29223
rect 4985 29183 5043 29189
rect 9217 29223 9275 29229
rect 9217 29189 9229 29223
rect 9263 29220 9275 29223
rect 9674 29220 9680 29232
rect 9263 29192 9680 29220
rect 9263 29189 9275 29192
rect 9217 29183 9275 29189
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 12710 29180 12716 29232
rect 12768 29180 12774 29232
rect 15194 29180 15200 29232
rect 15252 29220 15258 29232
rect 15473 29223 15531 29229
rect 15473 29220 15485 29223
rect 15252 29192 15485 29220
rect 15252 29180 15258 29192
rect 15473 29189 15485 29192
rect 15519 29220 15531 29223
rect 16853 29223 16911 29229
rect 16853 29220 16865 29223
rect 15519 29192 16865 29220
rect 15519 29189 15531 29192
rect 15473 29183 15531 29189
rect 16853 29189 16865 29192
rect 16899 29189 16911 29223
rect 16853 29183 16911 29189
rect 3973 29155 4031 29161
rect 3973 29121 3985 29155
rect 4019 29152 4031 29155
rect 4154 29152 4160 29164
rect 4019 29124 4160 29152
rect 4019 29121 4031 29124
rect 3973 29115 4031 29121
rect 4154 29112 4160 29124
rect 4212 29112 4218 29164
rect 12728 29152 12756 29180
rect 12989 29155 13047 29161
rect 12989 29152 13001 29155
rect 12728 29124 13001 29152
rect 12989 29121 13001 29124
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 13170 29112 13176 29164
rect 13228 29112 13234 29164
rect 15565 29155 15623 29161
rect 15565 29121 15577 29155
rect 15611 29152 15623 29155
rect 16298 29152 16304 29164
rect 15611 29124 16304 29152
rect 15611 29121 15623 29124
rect 15565 29115 15623 29121
rect 16298 29112 16304 29124
rect 16356 29112 16362 29164
rect 4062 29084 4068 29096
rect 1719 29056 2728 29084
rect 4023 29056 4068 29084
rect 1719 29053 1731 29056
rect 1673 29047 1731 29053
rect 4062 29044 4068 29056
rect 4120 29044 4126 29096
rect 4522 29084 4528 29096
rect 4483 29056 4528 29084
rect 4522 29044 4528 29056
rect 4580 29044 4586 29096
rect 4617 29087 4675 29093
rect 4617 29053 4629 29087
rect 4663 29053 4675 29087
rect 4617 29047 4675 29053
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 7006 29084 7012 29096
rect 6967 29056 7012 29084
rect 6825 29047 6883 29053
rect 3050 28976 3056 29028
rect 3108 29016 3114 29028
rect 3602 29016 3608 29028
rect 3108 28988 3608 29016
rect 3108 28976 3114 28988
rect 3602 28976 3608 28988
rect 3660 28976 3666 29028
rect 4080 29016 4108 29044
rect 4632 29016 4660 29047
rect 4080 28988 4660 29016
rect 4798 28976 4804 29028
rect 4856 29016 4862 29028
rect 6840 29016 6868 29047
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7190 29044 7196 29096
rect 7248 29084 7254 29096
rect 7469 29087 7527 29093
rect 7469 29084 7481 29087
rect 7248 29056 7481 29084
rect 7248 29044 7254 29056
rect 7469 29053 7481 29056
rect 7515 29053 7527 29087
rect 7469 29047 7527 29053
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29053 7619 29087
rect 7561 29047 7619 29053
rect 4856 28988 6868 29016
rect 7024 29016 7052 29044
rect 7576 29016 7604 29047
rect 8754 29044 8760 29096
rect 8812 29084 8818 29096
rect 9033 29087 9091 29093
rect 9033 29084 9045 29087
rect 8812 29056 9045 29084
rect 8812 29044 8818 29056
rect 9033 29053 9045 29056
rect 9079 29053 9091 29087
rect 10134 29084 10140 29096
rect 10095 29056 10140 29084
rect 9033 29047 9091 29053
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 10318 29084 10324 29096
rect 10279 29056 10324 29084
rect 10318 29044 10324 29056
rect 10376 29044 10382 29096
rect 10873 29087 10931 29093
rect 10873 29053 10885 29087
rect 10919 29053 10931 29087
rect 11054 29084 11060 29096
rect 11015 29056 11060 29084
rect 10873 29047 10931 29053
rect 7024 28988 7604 29016
rect 10888 29016 10916 29047
rect 11054 29044 11060 29056
rect 11112 29044 11118 29096
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 12713 29087 12771 29093
rect 12713 29084 12725 29087
rect 12584 29056 12725 29084
rect 12584 29044 12590 29056
rect 12713 29053 12725 29056
rect 12759 29053 12771 29087
rect 13188 29084 13216 29112
rect 15933 29087 15991 29093
rect 15933 29084 15945 29087
rect 13188 29056 15945 29084
rect 12713 29047 12771 29053
rect 15933 29053 15945 29056
rect 15979 29053 15991 29087
rect 15933 29047 15991 29053
rect 16482 29044 16488 29096
rect 16540 29084 16546 29096
rect 16761 29087 16819 29093
rect 16761 29084 16773 29087
rect 16540 29056 16773 29084
rect 16540 29044 16546 29056
rect 16761 29053 16773 29056
rect 16807 29053 16819 29087
rect 16761 29047 16819 29053
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29053 18107 29087
rect 18049 29047 18107 29053
rect 11238 29016 11244 29028
rect 10888 28988 11244 29016
rect 4856 28976 4862 28988
rect 11238 28976 11244 28988
rect 11296 28976 11302 29028
rect 14369 29019 14427 29025
rect 14369 28985 14381 29019
rect 14415 29016 14427 29019
rect 15197 29019 15255 29025
rect 14415 28988 15148 29016
rect 14415 28985 14427 28988
rect 14369 28979 14427 28985
rect 2774 28908 2780 28960
rect 2832 28948 2838 28960
rect 11330 28948 11336 28960
rect 2832 28920 2877 28948
rect 11291 28920 11336 28948
rect 2832 28908 2838 28920
rect 11330 28908 11336 28920
rect 11388 28908 11394 28960
rect 15120 28948 15148 28988
rect 15197 28985 15209 29019
rect 15243 29016 15255 29019
rect 15286 29016 15292 29028
rect 15243 28988 15292 29016
rect 15243 28985 15255 28988
rect 15197 28979 15255 28985
rect 15286 28976 15292 28988
rect 15344 28976 15350 29028
rect 15378 28976 15384 29028
rect 15436 29016 15442 29028
rect 18064 29016 18092 29047
rect 15436 28988 18092 29016
rect 15436 28976 15442 28988
rect 15396 28948 15424 28976
rect 15120 28920 15424 28948
rect 1104 28858 24840 28880
rect 1104 28806 8912 28858
rect 8964 28806 8976 28858
rect 9028 28806 9040 28858
rect 9092 28806 9104 28858
rect 9156 28806 16843 28858
rect 16895 28806 16907 28858
rect 16959 28806 16971 28858
rect 17023 28806 17035 28858
rect 17087 28806 24840 28858
rect 1104 28784 24840 28806
rect 3053 28747 3111 28753
rect 3053 28713 3065 28747
rect 3099 28744 3111 28747
rect 4062 28744 4068 28756
rect 3099 28716 4068 28744
rect 3099 28713 3111 28716
rect 3053 28707 3111 28713
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 4157 28747 4215 28753
rect 4157 28713 4169 28747
rect 4203 28744 4215 28747
rect 4203 28716 4568 28744
rect 4203 28713 4215 28716
rect 4157 28707 4215 28713
rect 3786 28636 3792 28688
rect 3844 28676 3850 28688
rect 4249 28679 4307 28685
rect 4249 28676 4261 28679
rect 3844 28648 4261 28676
rect 3844 28636 3850 28648
rect 4249 28645 4261 28648
rect 4295 28645 4307 28679
rect 4249 28639 4307 28645
rect 4338 28636 4344 28688
rect 4396 28676 4402 28688
rect 4396 28648 4476 28676
rect 4396 28636 4402 28648
rect 1857 28611 1915 28617
rect 1857 28577 1869 28611
rect 1903 28608 1915 28611
rect 2682 28608 2688 28620
rect 1903 28580 2688 28608
rect 1903 28577 1915 28580
rect 1857 28571 1915 28577
rect 2682 28568 2688 28580
rect 2740 28568 2746 28620
rect 2869 28611 2927 28617
rect 2869 28577 2881 28611
rect 2915 28608 2927 28611
rect 2958 28608 2964 28620
rect 2915 28580 2964 28608
rect 2915 28577 2927 28580
rect 2869 28571 2927 28577
rect 2958 28568 2964 28580
rect 3016 28568 3022 28620
rect 1486 28500 1492 28552
rect 1544 28540 1550 28552
rect 3050 28540 3056 28552
rect 1544 28512 3056 28540
rect 1544 28500 1550 28512
rect 3050 28500 3056 28512
rect 3108 28540 3114 28552
rect 4448 28549 4476 28648
rect 4540 28608 4568 28716
rect 5810 28704 5816 28756
rect 5868 28744 5874 28756
rect 6822 28744 6828 28756
rect 5868 28716 6828 28744
rect 5868 28704 5874 28716
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 15102 28704 15108 28756
rect 15160 28744 15166 28756
rect 15378 28744 15384 28756
rect 15160 28716 15384 28744
rect 15160 28704 15166 28716
rect 15378 28704 15384 28716
rect 15436 28704 15442 28756
rect 17586 28744 17592 28756
rect 17547 28716 17592 28744
rect 17586 28704 17592 28716
rect 17644 28704 17650 28756
rect 11701 28679 11759 28685
rect 11701 28645 11713 28679
rect 11747 28676 11759 28679
rect 13722 28676 13728 28688
rect 11747 28648 13728 28676
rect 11747 28645 11759 28648
rect 11701 28639 11759 28645
rect 13722 28636 13728 28648
rect 13780 28676 13786 28688
rect 13780 28648 17540 28676
rect 13780 28636 13786 28648
rect 5813 28611 5871 28617
rect 5813 28608 5825 28611
rect 4540 28580 5825 28608
rect 5813 28577 5825 28580
rect 5859 28577 5871 28611
rect 5813 28571 5871 28577
rect 6178 28568 6184 28620
rect 6236 28608 6242 28620
rect 8294 28608 8300 28620
rect 6236 28580 8300 28608
rect 6236 28568 6242 28580
rect 8294 28568 8300 28580
rect 8352 28568 8358 28620
rect 10321 28611 10379 28617
rect 10321 28577 10333 28611
rect 10367 28608 10379 28611
rect 11330 28608 11336 28620
rect 10367 28580 11336 28608
rect 10367 28577 10379 28580
rect 10321 28571 10379 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 12618 28568 12624 28620
rect 12676 28608 12682 28620
rect 12713 28611 12771 28617
rect 12713 28608 12725 28611
rect 12676 28580 12725 28608
rect 12676 28568 12682 28580
rect 12713 28577 12725 28580
rect 12759 28608 12771 28611
rect 13265 28611 13323 28617
rect 13265 28608 13277 28611
rect 12759 28580 13277 28608
rect 12759 28577 12771 28580
rect 12713 28571 12771 28577
rect 13265 28577 13277 28580
rect 13311 28577 13323 28611
rect 13265 28571 13323 28577
rect 13449 28611 13507 28617
rect 13449 28577 13461 28611
rect 13495 28608 13507 28611
rect 15194 28608 15200 28620
rect 13495 28580 15200 28608
rect 13495 28577 13507 28580
rect 13449 28571 13507 28577
rect 15194 28568 15200 28580
rect 15252 28568 15258 28620
rect 16114 28608 16120 28620
rect 16075 28580 16120 28608
rect 16114 28568 16120 28580
rect 16172 28568 16178 28620
rect 17512 28617 17540 28648
rect 16485 28611 16543 28617
rect 16485 28608 16497 28611
rect 16316 28580 16497 28608
rect 4157 28543 4215 28549
rect 4157 28540 4169 28543
rect 3108 28512 4169 28540
rect 3108 28500 3114 28512
rect 4157 28509 4169 28512
rect 4203 28509 4215 28543
rect 4157 28503 4215 28509
rect 4396 28543 4476 28549
rect 4396 28509 4408 28543
rect 4442 28512 4476 28543
rect 4617 28543 4675 28549
rect 4442 28509 4454 28512
rect 4396 28503 4454 28509
rect 4617 28509 4629 28543
rect 4663 28540 4675 28543
rect 4798 28540 4804 28552
rect 4663 28512 4804 28540
rect 4663 28509 4675 28512
rect 4617 28503 4675 28509
rect 4798 28500 4804 28512
rect 4856 28500 4862 28552
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28540 6147 28543
rect 6822 28540 6828 28552
rect 6135 28512 6828 28540
rect 6135 28509 6147 28512
rect 6089 28503 6147 28509
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28540 10103 28543
rect 12342 28540 12348 28552
rect 10091 28512 12348 28540
rect 10091 28509 10103 28512
rect 10045 28503 10103 28509
rect 12342 28500 12348 28512
rect 12400 28500 12406 28552
rect 12526 28540 12532 28552
rect 12487 28512 12532 28540
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 16209 28543 16267 28549
rect 16209 28540 16221 28543
rect 15896 28512 16221 28540
rect 15896 28500 15902 28512
rect 16209 28509 16221 28512
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 1949 28475 2007 28481
rect 1949 28441 1961 28475
rect 1995 28472 2007 28475
rect 4522 28472 4528 28484
rect 1995 28444 4528 28472
rect 1995 28441 2007 28444
rect 1949 28435 2007 28441
rect 4522 28432 4528 28444
rect 4580 28472 4586 28484
rect 5258 28472 5264 28484
rect 4580 28444 5264 28472
rect 4580 28432 4586 28444
rect 5258 28432 5264 28444
rect 5316 28432 5322 28484
rect 16022 28432 16028 28484
rect 16080 28472 16086 28484
rect 16316 28472 16344 28580
rect 16485 28577 16497 28580
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 17497 28611 17555 28617
rect 17497 28577 17509 28611
rect 17543 28577 17555 28611
rect 17497 28571 17555 28577
rect 16574 28540 16580 28552
rect 16535 28512 16580 28540
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 16080 28444 16344 28472
rect 16080 28432 16086 28444
rect 3970 28364 3976 28416
rect 4028 28404 4034 28416
rect 4338 28404 4344 28416
rect 4028 28376 4344 28404
rect 4028 28364 4034 28376
rect 4338 28364 4344 28376
rect 4396 28364 4402 28416
rect 4709 28407 4767 28413
rect 4709 28373 4721 28407
rect 4755 28404 4767 28407
rect 4798 28404 4804 28416
rect 4755 28376 4804 28404
rect 4755 28373 4767 28376
rect 4709 28367 4767 28373
rect 4798 28364 4804 28376
rect 4856 28364 4862 28416
rect 6454 28364 6460 28416
rect 6512 28404 6518 28416
rect 7193 28407 7251 28413
rect 7193 28404 7205 28407
rect 6512 28376 7205 28404
rect 6512 28364 6518 28376
rect 7193 28373 7205 28376
rect 7239 28373 7251 28407
rect 7193 28367 7251 28373
rect 7282 28364 7288 28416
rect 7340 28404 7346 28416
rect 8481 28407 8539 28413
rect 8481 28404 8493 28407
rect 7340 28376 8493 28404
rect 7340 28364 7346 28376
rect 8481 28373 8493 28376
rect 8527 28373 8539 28407
rect 8481 28367 8539 28373
rect 13725 28407 13783 28413
rect 13725 28373 13737 28407
rect 13771 28404 13783 28407
rect 13906 28404 13912 28416
rect 13771 28376 13912 28404
rect 13771 28373 13783 28376
rect 13725 28367 13783 28373
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 15562 28404 15568 28416
rect 15523 28376 15568 28404
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 1104 28314 24840 28336
rect 1104 28262 4947 28314
rect 4999 28262 5011 28314
rect 5063 28262 5075 28314
rect 5127 28262 5139 28314
rect 5191 28262 12878 28314
rect 12930 28262 12942 28314
rect 12994 28262 13006 28314
rect 13058 28262 13070 28314
rect 13122 28262 20808 28314
rect 20860 28262 20872 28314
rect 20924 28262 20936 28314
rect 20988 28262 21000 28314
rect 21052 28262 24840 28314
rect 1104 28240 24840 28262
rect 2774 28160 2780 28212
rect 2832 28200 2838 28212
rect 2832 28172 2877 28200
rect 2832 28160 2838 28172
rect 3142 28160 3148 28212
rect 3200 28200 3206 28212
rect 11057 28203 11115 28209
rect 11057 28200 11069 28203
rect 3200 28172 11069 28200
rect 3200 28160 3206 28172
rect 11057 28169 11069 28172
rect 11103 28169 11115 28203
rect 12618 28200 12624 28212
rect 12579 28172 12624 28200
rect 11057 28163 11115 28169
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 15930 28160 15936 28212
rect 15988 28200 15994 28212
rect 18141 28203 18199 28209
rect 18141 28200 18153 28203
rect 15988 28172 18153 28200
rect 15988 28160 15994 28172
rect 18141 28169 18153 28172
rect 18187 28169 18199 28203
rect 18141 28163 18199 28169
rect 7190 28132 7196 28144
rect 5000 28104 7196 28132
rect 4614 28064 4620 28076
rect 4575 28036 4620 28064
rect 4614 28024 4620 28036
rect 4672 28024 4678 28076
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27996 1455 27999
rect 1486 27996 1492 28008
rect 1443 27968 1492 27996
rect 1443 27965 1455 27968
rect 1397 27959 1455 27965
rect 1486 27956 1492 27968
rect 1544 27956 1550 28008
rect 1670 27996 1676 28008
rect 1631 27968 1676 27996
rect 1670 27956 1676 27968
rect 1728 27956 1734 28008
rect 2866 27956 2872 28008
rect 2924 27996 2930 28008
rect 5000 28005 5028 28104
rect 7190 28092 7196 28104
rect 7248 28092 7254 28144
rect 8662 28092 8668 28144
rect 8720 28132 8726 28144
rect 9125 28135 9183 28141
rect 9125 28132 9137 28135
rect 8720 28104 9137 28132
rect 8720 28092 8726 28104
rect 9125 28101 9137 28104
rect 9171 28101 9183 28135
rect 9125 28095 9183 28101
rect 9674 28092 9680 28144
rect 9732 28132 9738 28144
rect 9732 28104 12480 28132
rect 9732 28092 9738 28104
rect 5258 28024 5264 28076
rect 5316 28064 5322 28076
rect 5445 28067 5503 28073
rect 5445 28064 5457 28067
rect 5316 28036 5457 28064
rect 5316 28024 5322 28036
rect 5445 28033 5457 28036
rect 5491 28033 5503 28067
rect 5445 28027 5503 28033
rect 8018 28024 8024 28076
rect 8076 28064 8082 28076
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 8076 28036 10609 28064
rect 8076 28024 8082 28036
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 10597 28027 10655 28033
rect 4985 27999 5043 28005
rect 4985 27996 4997 27999
rect 2924 27968 4997 27996
rect 2924 27956 2930 27968
rect 4985 27965 4997 27968
rect 5031 27965 5043 27999
rect 4985 27959 5043 27965
rect 5169 27999 5227 28005
rect 5169 27965 5181 27999
rect 5215 27996 5227 27999
rect 5350 27996 5356 28008
rect 5215 27968 5356 27996
rect 5215 27965 5227 27968
rect 5169 27959 5227 27965
rect 5350 27956 5356 27968
rect 5408 27956 5414 28008
rect 5537 27999 5595 28005
rect 5537 27965 5549 27999
rect 5583 27996 5595 27999
rect 5626 27996 5632 28008
rect 5583 27968 5632 27996
rect 5583 27965 5595 27968
rect 5537 27959 5595 27965
rect 5626 27956 5632 27968
rect 5684 27956 5690 28008
rect 7558 27996 7564 28008
rect 7519 27968 7564 27996
rect 7558 27956 7564 27968
rect 7616 27956 7622 28008
rect 7742 27996 7748 28008
rect 7703 27968 7748 27996
rect 7742 27956 7748 27968
rect 7800 27956 7806 28008
rect 8205 27999 8263 28005
rect 8205 27965 8217 27999
rect 8251 27996 8263 27999
rect 9033 27999 9091 28005
rect 9033 27996 9045 27999
rect 8251 27968 9045 27996
rect 8251 27965 8263 27968
rect 8205 27959 8263 27965
rect 9033 27965 9045 27968
rect 9079 27965 9091 27999
rect 9033 27959 9091 27965
rect 9309 27999 9367 28005
rect 9309 27965 9321 27999
rect 9355 27996 9367 27999
rect 9858 27996 9864 28008
rect 9355 27968 9864 27996
rect 9355 27965 9367 27968
rect 9309 27959 9367 27965
rect 9858 27956 9864 27968
rect 9916 27956 9922 28008
rect 10870 27996 10876 28008
rect 10831 27968 10876 27996
rect 10870 27956 10876 27968
rect 10928 27956 10934 28008
rect 12452 28005 12480 28104
rect 13906 28064 13912 28076
rect 13867 28036 13912 28064
rect 13906 28024 13912 28036
rect 13964 28024 13970 28076
rect 12437 27999 12495 28005
rect 12437 27965 12449 27999
rect 12483 27965 12495 27999
rect 12437 27959 12495 27965
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 15378 27996 15384 28008
rect 13679 27968 15384 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 16206 27996 16212 28008
rect 16167 27968 16212 27996
rect 16206 27956 16212 27968
rect 16264 27956 16270 28008
rect 16393 27999 16451 28005
rect 16393 27965 16405 27999
rect 16439 27996 16451 27999
rect 16482 27996 16488 28008
rect 16439 27968 16488 27996
rect 16439 27965 16451 27968
rect 16393 27959 16451 27965
rect 5902 27888 5908 27940
rect 5960 27928 5966 27940
rect 7653 27931 7711 27937
rect 7653 27928 7665 27931
rect 5960 27900 7665 27928
rect 5960 27888 5966 27900
rect 7653 27897 7665 27900
rect 7699 27897 7711 27931
rect 7653 27891 7711 27897
rect 10410 27888 10416 27940
rect 10468 27928 10474 27940
rect 10781 27931 10839 27937
rect 10781 27928 10793 27931
rect 10468 27900 10793 27928
rect 10468 27888 10474 27900
rect 10781 27897 10793 27900
rect 10827 27897 10839 27931
rect 10781 27891 10839 27897
rect 15289 27931 15347 27937
rect 15289 27897 15301 27931
rect 15335 27928 15347 27931
rect 16408 27928 16436 27959
rect 16482 27956 16488 27968
rect 16540 27956 16546 28008
rect 16574 27956 16580 28008
rect 16632 27996 16638 28008
rect 16761 27999 16819 28005
rect 16761 27996 16773 27999
rect 16632 27968 16773 27996
rect 16632 27956 16638 27968
rect 16761 27965 16773 27968
rect 16807 27996 16819 27999
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 16807 27968 18061 27996
rect 16807 27965 16819 27968
rect 16761 27959 16819 27965
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 15335 27900 16436 27928
rect 15335 27897 15347 27900
rect 15289 27891 15347 27897
rect 2406 27820 2412 27872
rect 2464 27860 2470 27872
rect 2774 27860 2780 27872
rect 2464 27832 2780 27860
rect 2464 27820 2470 27832
rect 2774 27820 2780 27832
rect 2832 27820 2838 27872
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 9493 27863 9551 27869
rect 9493 27860 9505 27863
rect 8352 27832 9505 27860
rect 8352 27820 8358 27832
rect 9493 27829 9505 27832
rect 9539 27829 9551 27863
rect 9493 27823 9551 27829
rect 1104 27770 24840 27792
rect 1104 27718 8912 27770
rect 8964 27718 8976 27770
rect 9028 27718 9040 27770
rect 9092 27718 9104 27770
rect 9156 27718 16843 27770
rect 16895 27718 16907 27770
rect 16959 27718 16971 27770
rect 17023 27718 17035 27770
rect 17087 27718 24840 27770
rect 1104 27696 24840 27718
rect 1673 27659 1731 27665
rect 1673 27625 1685 27659
rect 1719 27656 1731 27659
rect 4890 27656 4896 27668
rect 1719 27628 4896 27656
rect 1719 27625 1731 27628
rect 1673 27619 1731 27625
rect 4890 27616 4896 27628
rect 4948 27616 4954 27668
rect 7006 27656 7012 27668
rect 6748 27628 7012 27656
rect 4062 27548 4068 27600
rect 4120 27588 4126 27600
rect 4120 27560 4292 27588
rect 4120 27548 4126 27560
rect 1581 27523 1639 27529
rect 1581 27489 1593 27523
rect 1627 27489 1639 27523
rect 1581 27483 1639 27489
rect 2593 27523 2651 27529
rect 2593 27489 2605 27523
rect 2639 27489 2651 27523
rect 2593 27483 2651 27489
rect 2777 27523 2835 27529
rect 2777 27489 2789 27523
rect 2823 27520 2835 27523
rect 3786 27520 3792 27532
rect 2823 27492 3792 27520
rect 2823 27489 2835 27492
rect 2777 27483 2835 27489
rect 1596 27384 1624 27483
rect 2608 27384 2636 27483
rect 3786 27480 3792 27492
rect 3844 27480 3850 27532
rect 4264 27529 4292 27560
rect 4249 27523 4307 27529
rect 4249 27489 4261 27523
rect 4295 27520 4307 27523
rect 4801 27523 4859 27529
rect 4801 27520 4813 27523
rect 4295 27492 4813 27520
rect 4295 27489 4307 27492
rect 4249 27483 4307 27489
rect 4801 27489 4813 27492
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 4985 27523 5043 27529
rect 4985 27520 4997 27523
rect 4948 27492 4997 27520
rect 4948 27480 4954 27492
rect 4985 27489 4997 27492
rect 5031 27520 5043 27523
rect 5258 27520 5264 27532
rect 5031 27492 5264 27520
rect 5031 27489 5043 27492
rect 4985 27483 5043 27489
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 6457 27523 6515 27529
rect 6457 27489 6469 27523
rect 6503 27520 6515 27523
rect 6748 27520 6776 27628
rect 7006 27616 7012 27628
rect 7064 27616 7070 27668
rect 8202 27616 8208 27668
rect 8260 27656 8266 27668
rect 8478 27656 8484 27668
rect 8260 27628 8484 27656
rect 8260 27616 8266 27628
rect 8478 27616 8484 27628
rect 8536 27616 8542 27668
rect 6822 27548 6828 27600
rect 6880 27588 6886 27600
rect 7561 27591 7619 27597
rect 7561 27588 7573 27591
rect 6880 27560 7573 27588
rect 6880 27548 6886 27560
rect 7561 27557 7573 27560
rect 7607 27557 7619 27591
rect 10413 27591 10471 27597
rect 7561 27551 7619 27557
rect 8496 27560 10088 27588
rect 6914 27520 6920 27532
rect 6503 27492 6776 27520
rect 6875 27492 6920 27520
rect 6503 27489 6515 27492
rect 6457 27483 6515 27489
rect 6914 27480 6920 27492
rect 6972 27480 6978 27532
rect 7006 27480 7012 27532
rect 7064 27520 7070 27532
rect 8496 27529 8524 27560
rect 8481 27523 8539 27529
rect 7064 27492 7109 27520
rect 7064 27480 7070 27492
rect 8481 27489 8493 27523
rect 8527 27489 8539 27523
rect 9674 27520 9680 27532
rect 9635 27492 9680 27520
rect 8481 27483 8539 27489
rect 9674 27480 9680 27492
rect 9732 27480 9738 27532
rect 9766 27480 9772 27532
rect 9824 27520 9830 27532
rect 9953 27523 10011 27529
rect 9824 27492 9869 27520
rect 9824 27480 9830 27492
rect 9953 27489 9965 27523
rect 9999 27489 10011 27523
rect 9953 27483 10011 27489
rect 3145 27455 3203 27461
rect 3145 27421 3157 27455
rect 3191 27452 3203 27455
rect 3970 27452 3976 27464
rect 3191 27424 3976 27452
rect 3191 27421 3203 27424
rect 3145 27415 3203 27421
rect 3970 27412 3976 27424
rect 4028 27412 4034 27464
rect 4154 27452 4160 27464
rect 4115 27424 4160 27452
rect 4154 27412 4160 27424
rect 4212 27412 4218 27464
rect 6270 27452 6276 27464
rect 6231 27424 6276 27452
rect 6270 27412 6276 27424
rect 6328 27412 6334 27464
rect 8386 27412 8392 27464
rect 8444 27452 8450 27464
rect 8938 27452 8944 27464
rect 8444 27424 8944 27452
rect 8444 27412 8450 27424
rect 8938 27412 8944 27424
rect 8996 27412 9002 27464
rect 9858 27412 9864 27464
rect 9916 27452 9922 27464
rect 9968 27452 9996 27483
rect 9916 27424 9996 27452
rect 10060 27452 10088 27560
rect 10413 27557 10425 27591
rect 10459 27588 10471 27591
rect 10870 27588 10876 27600
rect 10459 27560 10876 27588
rect 10459 27557 10471 27560
rect 10413 27551 10471 27557
rect 10870 27548 10876 27560
rect 10928 27548 10934 27600
rect 13173 27591 13231 27597
rect 13173 27557 13185 27591
rect 13219 27588 13231 27591
rect 13262 27588 13268 27600
rect 13219 27560 13268 27588
rect 13219 27557 13231 27560
rect 13173 27551 13231 27557
rect 13262 27548 13268 27560
rect 13320 27548 13326 27600
rect 15286 27588 15292 27600
rect 13832 27560 15292 27588
rect 10226 27480 10232 27532
rect 10284 27520 10290 27532
rect 11241 27523 11299 27529
rect 11241 27520 11253 27523
rect 10284 27492 11253 27520
rect 10284 27480 10290 27492
rect 11241 27489 11253 27492
rect 11287 27489 11299 27523
rect 11241 27483 11299 27489
rect 11330 27480 11336 27532
rect 11388 27520 11394 27532
rect 13832 27529 13860 27560
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 11425 27523 11483 27529
rect 11425 27520 11437 27523
rect 11388 27492 11437 27520
rect 11388 27480 11394 27492
rect 11425 27489 11437 27492
rect 11471 27489 11483 27523
rect 11425 27483 11483 27489
rect 13817 27523 13875 27529
rect 13817 27489 13829 27523
rect 13863 27489 13875 27523
rect 13817 27483 13875 27489
rect 14185 27523 14243 27529
rect 14185 27489 14197 27523
rect 14231 27520 14243 27523
rect 14369 27523 14427 27529
rect 14231 27492 14320 27520
rect 14231 27489 14243 27492
rect 14185 27483 14243 27489
rect 11348 27452 11376 27480
rect 10060 27424 11376 27452
rect 9916 27412 9922 27424
rect 11606 27412 11612 27464
rect 11664 27452 11670 27464
rect 13262 27452 13268 27464
rect 11664 27424 13268 27452
rect 11664 27412 11670 27424
rect 13262 27412 13268 27424
rect 13320 27412 13326 27464
rect 13909 27455 13967 27461
rect 13909 27452 13921 27455
rect 13832 27424 13921 27452
rect 13832 27396 13860 27424
rect 13909 27421 13921 27424
rect 13955 27421 13967 27455
rect 13909 27415 13967 27421
rect 12710 27384 12716 27396
rect 1596 27356 2176 27384
rect 2608 27356 12716 27384
rect 2148 27316 2176 27356
rect 12710 27344 12716 27356
rect 12768 27344 12774 27396
rect 13814 27344 13820 27396
rect 13872 27344 13878 27396
rect 2774 27316 2780 27328
rect 2148 27288 2780 27316
rect 2774 27276 2780 27288
rect 2832 27276 2838 27328
rect 3142 27276 3148 27328
rect 3200 27316 3206 27328
rect 5261 27319 5319 27325
rect 5261 27316 5273 27319
rect 3200 27288 5273 27316
rect 3200 27276 3206 27288
rect 5261 27285 5273 27288
rect 5307 27285 5319 27319
rect 5261 27279 5319 27285
rect 5534 27276 5540 27328
rect 5592 27316 5598 27328
rect 6822 27316 6828 27328
rect 5592 27288 6828 27316
rect 5592 27276 5598 27288
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 7650 27276 7656 27328
rect 7708 27316 7714 27328
rect 8662 27316 8668 27328
rect 7708 27288 8668 27316
rect 7708 27276 7714 27288
rect 8662 27276 8668 27288
rect 8720 27276 8726 27328
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 11112 27288 11529 27316
rect 11112 27276 11118 27288
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 14292 27316 14320 27492
rect 14369 27489 14381 27523
rect 14415 27520 14427 27523
rect 15194 27520 15200 27532
rect 14415 27492 15200 27520
rect 14415 27489 14427 27492
rect 14369 27483 14427 27489
rect 15194 27480 15200 27492
rect 15252 27480 15258 27532
rect 15378 27480 15384 27532
rect 15436 27480 15442 27532
rect 15562 27520 15568 27532
rect 15523 27492 15568 27520
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 17773 27523 17831 27529
rect 17773 27489 17785 27523
rect 17819 27489 17831 27523
rect 17773 27483 17831 27489
rect 15289 27455 15347 27461
rect 15289 27421 15301 27455
rect 15335 27452 15347 27455
rect 15396 27452 15424 27480
rect 15335 27424 15424 27452
rect 15335 27421 15347 27424
rect 15289 27415 15347 27421
rect 16022 27412 16028 27464
rect 16080 27452 16086 27464
rect 16669 27455 16727 27461
rect 16669 27452 16681 27455
rect 16080 27424 16681 27452
rect 16080 27412 16086 27424
rect 16669 27421 16681 27424
rect 16715 27452 16727 27455
rect 17788 27452 17816 27483
rect 16715 27424 17816 27452
rect 16715 27421 16727 27424
rect 16669 27415 16727 27421
rect 15562 27316 15568 27328
rect 14292 27288 15568 27316
rect 11517 27279 11575 27285
rect 15562 27276 15568 27288
rect 15620 27276 15626 27328
rect 16206 27276 16212 27328
rect 16264 27316 16270 27328
rect 17865 27319 17923 27325
rect 17865 27316 17877 27319
rect 16264 27288 17877 27316
rect 16264 27276 16270 27288
rect 17865 27285 17877 27288
rect 17911 27285 17923 27319
rect 17865 27279 17923 27285
rect 1104 27226 24840 27248
rect 1104 27174 4947 27226
rect 4999 27174 5011 27226
rect 5063 27174 5075 27226
rect 5127 27174 5139 27226
rect 5191 27174 12878 27226
rect 12930 27174 12942 27226
rect 12994 27174 13006 27226
rect 13058 27174 13070 27226
rect 13122 27174 20808 27226
rect 20860 27174 20872 27226
rect 20924 27174 20936 27226
rect 20988 27174 21000 27226
rect 21052 27174 24840 27226
rect 1104 27152 24840 27174
rect 3050 27112 3056 27124
rect 2884 27084 3056 27112
rect 2884 26988 2912 27084
rect 3050 27072 3056 27084
rect 3108 27072 3114 27124
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 6270 27112 6276 27124
rect 4212 27084 6276 27112
rect 4212 27072 4218 27084
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 6822 27072 6828 27124
rect 6880 27112 6886 27124
rect 8846 27112 8852 27124
rect 6880 27084 8852 27112
rect 6880 27072 6886 27084
rect 8846 27072 8852 27084
rect 8904 27072 8910 27124
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 10045 27115 10103 27121
rect 10045 27112 10057 27115
rect 9732 27084 10057 27112
rect 9732 27072 9738 27084
rect 10045 27081 10057 27084
rect 10091 27081 10103 27115
rect 11422 27112 11428 27124
rect 11383 27084 11428 27112
rect 10045 27075 10103 27081
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 11974 27072 11980 27124
rect 12032 27112 12038 27124
rect 12342 27112 12348 27124
rect 12032 27084 12348 27112
rect 12032 27072 12038 27084
rect 12342 27072 12348 27084
rect 12400 27072 12406 27124
rect 15289 27115 15347 27121
rect 15289 27081 15301 27115
rect 15335 27112 15347 27115
rect 16022 27112 16028 27124
rect 15335 27084 16028 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 16022 27072 16028 27084
rect 16080 27072 16086 27124
rect 16114 27072 16120 27124
rect 16172 27112 16178 27124
rect 16485 27115 16543 27121
rect 16485 27112 16497 27115
rect 16172 27084 16497 27112
rect 16172 27072 16178 27084
rect 16485 27081 16497 27084
rect 16531 27081 16543 27115
rect 16485 27075 16543 27081
rect 3970 27004 3976 27056
rect 4028 27044 4034 27056
rect 8294 27044 8300 27056
rect 4028 27016 8300 27044
rect 4028 27004 4034 27016
rect 8294 27004 8300 27016
rect 8352 27004 8358 27056
rect 12066 27004 12072 27056
rect 12124 27044 12130 27056
rect 12621 27047 12679 27053
rect 12621 27044 12633 27047
rect 12124 27016 12633 27044
rect 12124 27004 12130 27016
rect 12621 27013 12633 27016
rect 12667 27013 12679 27047
rect 12621 27007 12679 27013
rect 2866 26936 2872 26988
rect 2924 26976 2930 26988
rect 3142 26976 3148 26988
rect 2924 26948 3017 26976
rect 3103 26948 3148 26976
rect 2924 26936 2930 26948
rect 3142 26936 3148 26948
rect 3200 26936 3206 26988
rect 3786 26936 3792 26988
rect 3844 26976 3850 26988
rect 4062 26976 4068 26988
rect 3844 26948 4068 26976
rect 3844 26936 3850 26948
rect 4062 26936 4068 26948
rect 4120 26936 4126 26988
rect 4154 26936 4160 26988
rect 4212 26976 4218 26988
rect 4522 26976 4528 26988
rect 4212 26948 4528 26976
rect 4212 26936 4218 26948
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 5905 26979 5963 26985
rect 5000 26948 5672 26976
rect 1765 26911 1823 26917
rect 1765 26877 1777 26911
rect 1811 26908 1823 26911
rect 5000 26908 5028 26948
rect 5537 26911 5595 26917
rect 5537 26908 5549 26911
rect 1811 26880 5028 26908
rect 5276 26880 5549 26908
rect 1811 26877 1823 26880
rect 1765 26871 1823 26877
rect 4062 26800 4068 26852
rect 4120 26840 4126 26852
rect 5276 26840 5304 26880
rect 5537 26877 5549 26880
rect 5583 26877 5595 26911
rect 5644 26908 5672 26948
rect 5905 26945 5917 26979
rect 5951 26976 5963 26979
rect 7742 26976 7748 26988
rect 5951 26948 7748 26976
rect 5951 26945 5963 26948
rect 5905 26939 5963 26945
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 7852 26948 8432 26976
rect 6822 26908 6828 26920
rect 5644 26880 6828 26908
rect 5537 26871 5595 26877
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7650 26908 7656 26920
rect 6932 26880 7656 26908
rect 4120 26812 5304 26840
rect 4120 26800 4126 26812
rect 1946 26772 1952 26784
rect 1907 26744 1952 26772
rect 1946 26732 1952 26744
rect 2004 26732 2010 26784
rect 3142 26732 3148 26784
rect 3200 26772 3206 26784
rect 4249 26775 4307 26781
rect 4249 26772 4261 26775
rect 3200 26744 4261 26772
rect 3200 26732 3206 26744
rect 4249 26741 4261 26744
rect 4295 26741 4307 26775
rect 4249 26735 4307 26741
rect 4430 26732 4436 26784
rect 4488 26772 4494 26784
rect 4614 26772 4620 26784
rect 4488 26744 4620 26772
rect 4488 26732 4494 26744
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 5276 26772 5304 26812
rect 5353 26843 5411 26849
rect 5353 26809 5365 26843
rect 5399 26840 5411 26843
rect 6454 26840 6460 26852
rect 5399 26812 6460 26840
rect 5399 26809 5411 26812
rect 5353 26803 5411 26809
rect 6454 26800 6460 26812
rect 6512 26800 6518 26852
rect 6932 26840 6960 26880
rect 7650 26868 7656 26880
rect 7708 26868 7714 26920
rect 7852 26840 7880 26948
rect 8018 26908 8024 26920
rect 7979 26880 8024 26908
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 8294 26868 8300 26920
rect 8352 26917 8358 26920
rect 8352 26911 8375 26917
rect 8363 26877 8375 26911
rect 8404 26908 8432 26948
rect 8588 26948 9170 26976
rect 8588 26908 8616 26948
rect 8404 26880 8616 26908
rect 8757 26911 8815 26917
rect 8352 26871 8375 26877
rect 8757 26877 8769 26911
rect 8803 26908 8815 26911
rect 8846 26908 8852 26920
rect 8803 26880 8852 26908
rect 8803 26877 8815 26880
rect 8757 26871 8815 26877
rect 8352 26868 8358 26871
rect 8846 26868 8852 26880
rect 8904 26868 8910 26920
rect 8202 26840 8208 26852
rect 6840 26812 6960 26840
rect 7024 26812 7880 26840
rect 8163 26812 8208 26840
rect 6840 26772 6868 26812
rect 7024 26784 7052 26812
rect 8202 26800 8208 26812
rect 8260 26800 8266 26852
rect 8938 26840 8944 26852
rect 8404 26812 8944 26840
rect 8404 26784 8432 26812
rect 8938 26800 8944 26812
rect 8996 26800 9002 26852
rect 9142 26840 9170 26948
rect 9674 26936 9680 26988
rect 9732 26976 9738 26988
rect 13725 26979 13783 26985
rect 9732 26948 9904 26976
rect 9732 26936 9738 26948
rect 9214 26868 9220 26920
rect 9272 26908 9278 26920
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 9272 26880 9597 26908
rect 9272 26868 9278 26880
rect 9585 26877 9597 26880
rect 9631 26877 9643 26911
rect 9766 26908 9772 26920
rect 9727 26880 9772 26908
rect 9585 26871 9643 26877
rect 9766 26868 9772 26880
rect 9824 26868 9830 26920
rect 9876 26917 9904 26948
rect 13725 26945 13737 26979
rect 13771 26976 13783 26979
rect 14182 26976 14188 26988
rect 13771 26948 14188 26976
rect 13771 26945 13783 26948
rect 13725 26939 13783 26945
rect 14182 26936 14188 26948
rect 14240 26976 14246 26988
rect 15378 26976 15384 26988
rect 14240 26948 15384 26976
rect 14240 26936 14246 26948
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 15930 26936 15936 26988
rect 15988 26976 15994 26988
rect 15988 26948 16344 26976
rect 15988 26936 15994 26948
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26877 9919 26911
rect 9861 26871 9919 26877
rect 11241 26911 11299 26917
rect 11241 26877 11253 26911
rect 11287 26877 11299 26911
rect 12434 26908 12440 26920
rect 12395 26880 12440 26908
rect 11241 26871 11299 26877
rect 11256 26840 11284 26871
rect 12434 26868 12440 26880
rect 12492 26868 12498 26920
rect 13998 26908 14004 26920
rect 13959 26880 14004 26908
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 16206 26908 16212 26920
rect 16167 26880 16212 26908
rect 16206 26868 16212 26880
rect 16264 26868 16270 26920
rect 16316 26917 16344 26948
rect 16301 26911 16359 26917
rect 16301 26877 16313 26911
rect 16347 26877 16359 26911
rect 16301 26871 16359 26877
rect 16482 26868 16488 26920
rect 16540 26908 16546 26920
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 16540 26880 18061 26908
rect 16540 26868 16546 26880
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 9142 26812 11284 26840
rect 7006 26772 7012 26784
rect 5276 26744 6868 26772
rect 6919 26744 7012 26772
rect 7006 26732 7012 26744
rect 7064 26732 7070 26784
rect 7558 26732 7564 26784
rect 7616 26772 7622 26784
rect 8294 26772 8300 26784
rect 7616 26744 8300 26772
rect 7616 26732 7622 26744
rect 8294 26732 8300 26744
rect 8352 26732 8358 26784
rect 8386 26732 8392 26784
rect 8444 26732 8450 26784
rect 11256 26772 11284 26812
rect 15194 26772 15200 26784
rect 11256 26744 15200 26772
rect 15194 26732 15200 26744
rect 15252 26732 15258 26784
rect 18138 26772 18144 26784
rect 18099 26744 18144 26772
rect 18138 26732 18144 26744
rect 18196 26732 18202 26784
rect 1104 26682 24840 26704
rect 1104 26630 8912 26682
rect 8964 26630 8976 26682
rect 9028 26630 9040 26682
rect 9092 26630 9104 26682
rect 9156 26630 16843 26682
rect 16895 26630 16907 26682
rect 16959 26630 16971 26682
rect 17023 26630 17035 26682
rect 17087 26630 24840 26682
rect 1104 26608 24840 26630
rect 1486 26528 1492 26580
rect 1544 26568 1550 26580
rect 1762 26568 1768 26580
rect 1544 26540 1768 26568
rect 1544 26528 1550 26540
rect 1762 26528 1768 26540
rect 1820 26528 1826 26580
rect 3326 26528 3332 26580
rect 3384 26568 3390 26580
rect 3970 26568 3976 26580
rect 3384 26540 3976 26568
rect 3384 26528 3390 26540
rect 3970 26528 3976 26540
rect 4028 26528 4034 26580
rect 5994 26568 6000 26580
rect 5955 26540 6000 26568
rect 5994 26528 6000 26540
rect 6052 26528 6058 26580
rect 6914 26568 6920 26580
rect 6472 26540 6920 26568
rect 3786 26460 3792 26512
rect 3844 26500 3850 26512
rect 4617 26503 4675 26509
rect 4617 26500 4629 26503
rect 3844 26472 4629 26500
rect 3844 26460 3850 26472
rect 4617 26469 4629 26472
rect 4663 26469 4675 26503
rect 4617 26463 4675 26469
rect 2409 26435 2467 26441
rect 2409 26401 2421 26435
rect 2455 26432 2467 26435
rect 2590 26432 2596 26444
rect 2455 26404 2596 26432
rect 2455 26401 2467 26404
rect 2409 26395 2467 26401
rect 2590 26392 2596 26404
rect 2648 26392 2654 26444
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 3142 26432 3148 26444
rect 2832 26404 3148 26432
rect 2832 26392 2838 26404
rect 3142 26392 3148 26404
rect 3200 26392 3206 26444
rect 4062 26432 4068 26444
rect 4023 26404 4068 26432
rect 4062 26392 4068 26404
rect 4120 26392 4126 26444
rect 4157 26435 4215 26441
rect 4157 26401 4169 26435
rect 4203 26401 4215 26435
rect 4157 26395 4215 26401
rect 2222 26324 2228 26376
rect 2280 26364 2286 26376
rect 2317 26367 2375 26373
rect 2317 26364 2329 26367
rect 2280 26336 2329 26364
rect 2280 26324 2286 26336
rect 2317 26333 2329 26336
rect 2363 26333 2375 26367
rect 2317 26327 2375 26333
rect 2682 26324 2688 26376
rect 2740 26364 2746 26376
rect 2869 26367 2927 26373
rect 2869 26364 2881 26367
rect 2740 26336 2881 26364
rect 2740 26324 2746 26336
rect 2869 26333 2881 26336
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 3050 26324 3056 26376
rect 3108 26364 3114 26376
rect 4172 26364 4200 26395
rect 5810 26392 5816 26444
rect 5868 26432 5874 26444
rect 5994 26432 6000 26444
rect 5868 26404 6000 26432
rect 5868 26392 5874 26404
rect 5994 26392 6000 26404
rect 6052 26392 6058 26444
rect 6365 26435 6423 26441
rect 6365 26401 6377 26435
rect 6411 26432 6423 26435
rect 6472 26432 6500 26540
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 8202 26528 8208 26580
rect 8260 26568 8266 26580
rect 8389 26571 8447 26577
rect 8389 26568 8401 26571
rect 8260 26540 8401 26568
rect 8260 26528 8266 26540
rect 8389 26537 8401 26540
rect 8435 26537 8447 26571
rect 8389 26531 8447 26537
rect 8662 26528 8668 26580
rect 8720 26568 8726 26580
rect 9214 26568 9220 26580
rect 8720 26540 9220 26568
rect 8720 26528 8726 26540
rect 9214 26528 9220 26540
rect 9272 26528 9278 26580
rect 9766 26528 9772 26580
rect 9824 26568 9830 26580
rect 14001 26571 14059 26577
rect 14001 26568 14013 26571
rect 9824 26540 14013 26568
rect 9824 26528 9830 26540
rect 14001 26537 14013 26540
rect 14047 26537 14059 26571
rect 14001 26531 14059 26537
rect 7282 26500 7288 26512
rect 6564 26472 7288 26500
rect 6564 26441 6592 26472
rect 7282 26460 7288 26472
rect 7340 26460 7346 26512
rect 10410 26500 10416 26512
rect 10371 26472 10416 26500
rect 10410 26460 10416 26472
rect 10468 26460 10474 26512
rect 12710 26460 12716 26512
rect 12768 26500 12774 26512
rect 12897 26503 12955 26509
rect 12897 26500 12909 26503
rect 12768 26472 12909 26500
rect 12768 26460 12774 26472
rect 12897 26469 12909 26472
rect 12943 26500 12955 26503
rect 16482 26500 16488 26512
rect 12943 26472 16488 26500
rect 12943 26469 12955 26472
rect 12897 26463 12955 26469
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 6411 26404 6500 26432
rect 6549 26435 6607 26441
rect 6411 26401 6423 26404
rect 6365 26395 6423 26401
rect 6549 26401 6561 26435
rect 6595 26401 6607 26435
rect 6549 26395 6607 26401
rect 6917 26435 6975 26441
rect 6917 26401 6929 26435
rect 6963 26432 6975 26435
rect 7558 26432 7564 26444
rect 6963 26404 7564 26432
rect 6963 26401 6975 26404
rect 6917 26395 6975 26401
rect 7558 26392 7564 26404
rect 7616 26392 7622 26444
rect 7650 26392 7656 26444
rect 7708 26432 7714 26444
rect 7929 26435 7987 26441
rect 7929 26432 7941 26435
rect 7708 26404 7941 26432
rect 7708 26392 7714 26404
rect 7929 26401 7941 26404
rect 7975 26401 7987 26435
rect 7929 26395 7987 26401
rect 8205 26435 8263 26441
rect 8205 26401 8217 26435
rect 8251 26401 8263 26435
rect 8205 26395 8263 26401
rect 9677 26435 9735 26441
rect 9677 26401 9689 26435
rect 9723 26432 9735 26435
rect 9766 26432 9772 26444
rect 9723 26404 9772 26432
rect 9723 26401 9735 26404
rect 9677 26395 9735 26401
rect 3108 26336 4200 26364
rect 6825 26367 6883 26373
rect 3108 26324 3114 26336
rect 6825 26333 6837 26367
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 5258 26296 5264 26308
rect 4120 26268 5264 26296
rect 4120 26256 4126 26268
rect 5258 26256 5264 26268
rect 5316 26296 5322 26308
rect 6840 26296 6868 26327
rect 7006 26324 7012 26376
rect 7064 26364 7070 26376
rect 8220 26364 8248 26395
rect 9766 26392 9772 26404
rect 9824 26392 9830 26444
rect 9953 26435 10011 26441
rect 9953 26401 9965 26435
rect 9999 26401 10011 26435
rect 9953 26395 10011 26401
rect 11241 26435 11299 26441
rect 11241 26401 11253 26435
rect 11287 26432 11299 26435
rect 11974 26432 11980 26444
rect 11287 26404 11980 26432
rect 11287 26401 11299 26404
rect 11241 26395 11299 26401
rect 9968 26364 9996 26395
rect 11974 26392 11980 26404
rect 12032 26392 12038 26444
rect 13722 26432 13728 26444
rect 13683 26404 13728 26432
rect 13722 26392 13728 26404
rect 13780 26392 13786 26444
rect 13909 26435 13967 26441
rect 13909 26401 13921 26435
rect 13955 26401 13967 26435
rect 13909 26395 13967 26401
rect 11514 26364 11520 26376
rect 7064 26336 9996 26364
rect 11475 26336 11520 26364
rect 7064 26324 7070 26336
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 12710 26324 12716 26376
rect 12768 26364 12774 26376
rect 13924 26364 13952 26395
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 15289 26435 15347 26441
rect 15289 26432 15301 26435
rect 15252 26404 15301 26432
rect 15252 26392 15258 26404
rect 15289 26401 15301 26404
rect 15335 26432 15347 26435
rect 18046 26432 18052 26444
rect 15335 26404 18052 26432
rect 15335 26401 15347 26404
rect 15289 26395 15347 26401
rect 18046 26392 18052 26404
rect 18104 26392 18110 26444
rect 12768 26336 13952 26364
rect 12768 26324 12774 26336
rect 15378 26324 15384 26376
rect 15436 26364 15442 26376
rect 16022 26364 16028 26376
rect 15436 26336 16028 26364
rect 15436 26324 15442 26336
rect 16022 26324 16028 26336
rect 16080 26364 16086 26376
rect 16393 26367 16451 26373
rect 16393 26364 16405 26367
rect 16080 26336 16405 26364
rect 16080 26324 16086 26336
rect 16393 26333 16405 26336
rect 16439 26333 16451 26367
rect 16666 26364 16672 26376
rect 16627 26336 16672 26364
rect 16393 26327 16451 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 8018 26296 8024 26308
rect 5316 26268 6868 26296
rect 7979 26268 8024 26296
rect 5316 26256 5322 26268
rect 8018 26256 8024 26268
rect 8076 26256 8082 26308
rect 9769 26299 9827 26305
rect 9769 26265 9781 26299
rect 9815 26296 9827 26299
rect 10594 26296 10600 26308
rect 9815 26268 10600 26296
rect 9815 26265 9827 26268
rect 9769 26259 9827 26265
rect 10594 26256 10600 26268
rect 10652 26256 10658 26308
rect 1854 26228 1860 26240
rect 1815 26200 1860 26228
rect 1854 26188 1860 26200
rect 1912 26188 1918 26240
rect 3510 26188 3516 26240
rect 3568 26228 3574 26240
rect 4430 26228 4436 26240
rect 3568 26200 4436 26228
rect 3568 26188 3574 26200
rect 4430 26188 4436 26200
rect 4488 26188 4494 26240
rect 6454 26188 6460 26240
rect 6512 26228 6518 26240
rect 6822 26228 6828 26240
rect 6512 26200 6828 26228
rect 6512 26188 6518 26200
rect 6822 26188 6828 26200
rect 6880 26188 6886 26240
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 10410 26228 10416 26240
rect 9916 26200 10416 26228
rect 9916 26188 9922 26200
rect 10410 26188 10416 26200
rect 10468 26188 10474 26240
rect 15473 26231 15531 26237
rect 15473 26197 15485 26231
rect 15519 26228 15531 26231
rect 15562 26228 15568 26240
rect 15519 26200 15568 26228
rect 15519 26197 15531 26200
rect 15473 26191 15531 26197
rect 15562 26188 15568 26200
rect 15620 26188 15626 26240
rect 17954 26228 17960 26240
rect 17915 26200 17960 26228
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 1104 26138 24840 26160
rect 1104 26086 4947 26138
rect 4999 26086 5011 26138
rect 5063 26086 5075 26138
rect 5127 26086 5139 26138
rect 5191 26086 12878 26138
rect 12930 26086 12942 26138
rect 12994 26086 13006 26138
rect 13058 26086 13070 26138
rect 13122 26086 20808 26138
rect 20860 26086 20872 26138
rect 20924 26086 20936 26138
rect 20988 26086 21000 26138
rect 21052 26086 24840 26138
rect 1104 26064 24840 26086
rect 8018 26024 8024 26036
rect 7979 25996 8024 26024
rect 8018 25984 8024 25996
rect 8076 25984 8082 26036
rect 9490 25984 9496 26036
rect 9548 25984 9554 26036
rect 10594 26024 10600 26036
rect 10555 25996 10600 26024
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 13633 26027 13691 26033
rect 13633 25993 13645 26027
rect 13679 26024 13691 26027
rect 13998 26024 14004 26036
rect 13679 25996 14004 26024
rect 13679 25993 13691 25996
rect 13633 25987 13691 25993
rect 13998 25984 14004 25996
rect 14056 25984 14062 26036
rect 9508 25956 9536 25984
rect 12066 25956 12072 25968
rect 9508 25928 12072 25956
rect 12066 25916 12072 25928
rect 12124 25916 12130 25968
rect 18138 25956 18144 25968
rect 15396 25928 18144 25956
rect 15396 25900 15424 25928
rect 18138 25916 18144 25928
rect 18196 25916 18202 25968
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 1854 25888 1860 25900
rect 1719 25860 1860 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 1854 25848 1860 25860
rect 1912 25848 1918 25900
rect 3878 25848 3884 25900
rect 3936 25888 3942 25900
rect 3973 25891 4031 25897
rect 3973 25888 3985 25891
rect 3936 25860 3985 25888
rect 3936 25848 3942 25860
rect 3973 25857 3985 25860
rect 4019 25857 4031 25891
rect 3973 25851 4031 25857
rect 4338 25848 4344 25900
rect 4396 25888 4402 25900
rect 4433 25891 4491 25897
rect 4433 25888 4445 25891
rect 4396 25860 4445 25888
rect 4396 25848 4402 25860
rect 4433 25857 4445 25860
rect 4479 25857 4491 25891
rect 5350 25888 5356 25900
rect 4433 25851 4491 25857
rect 4632 25860 5356 25888
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25820 1455 25823
rect 2866 25820 2872 25832
rect 1443 25792 2872 25820
rect 1443 25789 1455 25792
rect 1397 25783 1455 25789
rect 2866 25780 2872 25792
rect 2924 25780 2930 25832
rect 4632 25829 4660 25860
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 7561 25891 7619 25897
rect 7561 25857 7573 25891
rect 7607 25888 7619 25891
rect 10137 25891 10195 25897
rect 10137 25888 10149 25891
rect 7607 25860 10149 25888
rect 7607 25857 7619 25860
rect 7561 25851 7619 25857
rect 10137 25857 10149 25860
rect 10183 25888 10195 25891
rect 11146 25888 11152 25900
rect 10183 25860 11152 25888
rect 10183 25857 10195 25860
rect 10137 25851 10195 25857
rect 11146 25848 11152 25860
rect 11204 25848 11210 25900
rect 14550 25848 14556 25900
rect 14608 25888 14614 25900
rect 14645 25891 14703 25897
rect 14645 25888 14657 25891
rect 14608 25860 14657 25888
rect 14608 25848 14614 25860
rect 14645 25857 14657 25860
rect 14691 25857 14703 25891
rect 15378 25888 15384 25900
rect 15291 25860 15384 25888
rect 14645 25851 14703 25857
rect 15378 25848 15384 25860
rect 15436 25848 15442 25900
rect 16206 25888 16212 25900
rect 15488 25860 16212 25888
rect 4617 25823 4675 25829
rect 4617 25789 4629 25823
rect 4663 25789 4675 25823
rect 4617 25783 4675 25789
rect 4985 25823 5043 25829
rect 4985 25789 4997 25823
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 5169 25823 5227 25829
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 5258 25820 5264 25832
rect 5215 25792 5264 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 3053 25755 3111 25761
rect 3053 25721 3065 25755
rect 3099 25752 3111 25755
rect 3142 25752 3148 25764
rect 3099 25724 3148 25752
rect 3099 25721 3111 25724
rect 3053 25715 3111 25721
rect 3142 25712 3148 25724
rect 3200 25712 3206 25764
rect 5000 25752 5028 25783
rect 5258 25780 5264 25792
rect 5316 25780 5322 25832
rect 7834 25820 7840 25832
rect 7795 25792 7840 25820
rect 7834 25780 7840 25792
rect 7892 25780 7898 25832
rect 8662 25780 8668 25832
rect 8720 25820 8726 25832
rect 9125 25823 9183 25829
rect 9125 25820 9137 25823
rect 8720 25792 9137 25820
rect 8720 25780 8726 25792
rect 9125 25789 9137 25792
rect 9171 25820 9183 25823
rect 9398 25820 9404 25832
rect 9171 25792 9404 25820
rect 9171 25789 9183 25792
rect 9125 25783 9183 25789
rect 9398 25780 9404 25792
rect 9456 25780 9462 25832
rect 10413 25823 10471 25829
rect 10413 25789 10425 25823
rect 10459 25820 10471 25823
rect 11054 25820 11060 25832
rect 10459 25792 11060 25820
rect 10459 25789 10471 25792
rect 10413 25783 10471 25789
rect 11054 25780 11060 25792
rect 11112 25780 11118 25832
rect 11422 25780 11428 25832
rect 11480 25820 11486 25832
rect 12437 25823 12495 25829
rect 12437 25820 12449 25823
rect 11480 25792 12449 25820
rect 11480 25780 11486 25792
rect 12437 25789 12449 25792
rect 12483 25789 12495 25823
rect 12618 25820 12624 25832
rect 12579 25792 12624 25820
rect 12437 25783 12495 25789
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25789 13231 25823
rect 13173 25783 13231 25789
rect 13357 25823 13415 25829
rect 13357 25789 13369 25823
rect 13403 25789 13415 25823
rect 15286 25820 15292 25832
rect 15247 25792 15292 25820
rect 13357 25783 13415 25789
rect 5626 25752 5632 25764
rect 5000 25724 5632 25752
rect 1946 25644 1952 25696
rect 2004 25684 2010 25696
rect 5000 25684 5028 25724
rect 5626 25712 5632 25724
rect 5684 25712 5690 25764
rect 7742 25752 7748 25764
rect 7703 25724 7748 25752
rect 7742 25712 7748 25724
rect 7800 25712 7806 25764
rect 8570 25712 8576 25764
rect 8628 25752 8634 25764
rect 9490 25752 9496 25764
rect 8628 25724 9496 25752
rect 8628 25712 8634 25724
rect 9490 25712 9496 25724
rect 9548 25712 9554 25764
rect 10321 25755 10379 25761
rect 10321 25721 10333 25755
rect 10367 25752 10379 25755
rect 10686 25752 10692 25764
rect 10367 25724 10692 25752
rect 10367 25721 10379 25724
rect 10321 25715 10379 25721
rect 10686 25712 10692 25724
rect 10744 25712 10750 25764
rect 12636 25752 12664 25780
rect 13188 25752 13216 25783
rect 12636 25724 13216 25752
rect 13372 25752 13400 25783
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 15488 25752 15516 25860
rect 15562 25780 15568 25832
rect 15620 25820 15626 25832
rect 15764 25829 15792 25860
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 15657 25823 15715 25829
rect 15657 25820 15669 25823
rect 15620 25792 15669 25820
rect 15620 25780 15626 25792
rect 15657 25789 15669 25792
rect 15703 25789 15715 25823
rect 15657 25783 15715 25789
rect 15749 25823 15807 25829
rect 15749 25789 15761 25823
rect 15795 25789 15807 25823
rect 15749 25783 15807 25789
rect 13372 25724 15516 25752
rect 15672 25752 15700 25783
rect 16574 25780 16580 25832
rect 16632 25820 16638 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16632 25792 16681 25820
rect 16632 25780 16638 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16669 25783 16727 25789
rect 16114 25752 16120 25764
rect 15672 25724 16120 25752
rect 16114 25712 16120 25724
rect 16172 25712 16178 25764
rect 2004 25656 5028 25684
rect 2004 25644 2010 25656
rect 7098 25644 7104 25696
rect 7156 25684 7162 25696
rect 8018 25684 8024 25696
rect 7156 25656 8024 25684
rect 7156 25644 7162 25656
rect 8018 25644 8024 25656
rect 8076 25644 8082 25696
rect 9214 25684 9220 25696
rect 9127 25656 9220 25684
rect 9214 25644 9220 25656
rect 9272 25684 9278 25696
rect 15194 25684 15200 25696
rect 9272 25656 15200 25684
rect 9272 25644 9278 25656
rect 15194 25644 15200 25656
rect 15252 25644 15258 25696
rect 16206 25644 16212 25696
rect 16264 25684 16270 25696
rect 16761 25687 16819 25693
rect 16761 25684 16773 25687
rect 16264 25656 16773 25684
rect 16264 25644 16270 25656
rect 16761 25653 16773 25656
rect 16807 25653 16819 25687
rect 16761 25647 16819 25653
rect 1104 25594 24840 25616
rect 1104 25542 8912 25594
rect 8964 25542 8976 25594
rect 9028 25542 9040 25594
rect 9092 25542 9104 25594
rect 9156 25542 16843 25594
rect 16895 25542 16907 25594
rect 16959 25542 16971 25594
rect 17023 25542 17035 25594
rect 17087 25542 24840 25594
rect 1104 25520 24840 25542
rect 5718 25440 5724 25492
rect 5776 25480 5782 25492
rect 5813 25483 5871 25489
rect 5813 25480 5825 25483
rect 5776 25452 5825 25480
rect 5776 25440 5782 25452
rect 5813 25449 5825 25452
rect 5859 25449 5871 25483
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 5813 25443 5871 25449
rect 7208 25452 9965 25480
rect 1397 25415 1455 25421
rect 1397 25381 1409 25415
rect 1443 25412 1455 25415
rect 1670 25412 1676 25424
rect 1443 25384 1676 25412
rect 1443 25381 1455 25384
rect 1397 25375 1455 25381
rect 1670 25372 1676 25384
rect 1728 25372 1734 25424
rect 3050 25412 3056 25424
rect 2056 25384 3056 25412
rect 1762 25304 1768 25356
rect 1820 25344 1826 25356
rect 2056 25353 2084 25384
rect 3050 25372 3056 25384
rect 3108 25372 3114 25424
rect 2041 25347 2099 25353
rect 2041 25344 2053 25347
rect 1820 25316 2053 25344
rect 1820 25304 1826 25316
rect 2041 25313 2053 25316
rect 2087 25313 2099 25347
rect 2406 25344 2412 25356
rect 2367 25316 2412 25344
rect 2041 25307 2099 25313
rect 2406 25304 2412 25316
rect 2464 25304 2470 25356
rect 2866 25304 2872 25356
rect 2924 25344 2930 25356
rect 4433 25347 4491 25353
rect 4433 25344 4445 25347
rect 2924 25316 4445 25344
rect 2924 25304 2930 25316
rect 4433 25313 4445 25316
rect 4479 25313 4491 25347
rect 7098 25344 7104 25356
rect 7059 25316 7104 25344
rect 4433 25307 4491 25313
rect 7098 25304 7104 25316
rect 7156 25304 7162 25356
rect 7208 25353 7236 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 9953 25443 10011 25449
rect 11514 25440 11520 25492
rect 11572 25480 11578 25492
rect 12253 25483 12311 25489
rect 12253 25480 12265 25483
rect 11572 25452 12265 25480
rect 11572 25440 11578 25452
rect 12253 25449 12265 25452
rect 12299 25449 12311 25483
rect 15930 25480 15936 25492
rect 12253 25443 12311 25449
rect 13096 25452 15936 25480
rect 7650 25412 7656 25424
rect 7611 25384 7656 25412
rect 7650 25372 7656 25384
rect 7708 25372 7714 25424
rect 13096 25412 13124 25452
rect 15930 25440 15936 25452
rect 15988 25440 15994 25492
rect 13262 25412 13268 25424
rect 11256 25384 13124 25412
rect 13223 25384 13268 25412
rect 11256 25356 11284 25384
rect 7193 25347 7251 25353
rect 7193 25313 7205 25347
rect 7239 25313 7251 25347
rect 7193 25307 7251 25313
rect 8481 25347 8539 25353
rect 8481 25313 8493 25347
rect 8527 25344 8539 25347
rect 8570 25344 8576 25356
rect 8527 25316 8576 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 8570 25304 8576 25316
rect 8628 25304 8634 25356
rect 9674 25344 9680 25356
rect 9635 25316 9680 25344
rect 9674 25304 9680 25316
rect 9732 25304 9738 25356
rect 9861 25347 9919 25353
rect 9861 25313 9873 25347
rect 9907 25313 9919 25347
rect 11238 25344 11244 25356
rect 11199 25316 11244 25344
rect 9861 25307 9919 25313
rect 2133 25279 2191 25285
rect 2133 25245 2145 25279
rect 2179 25276 2191 25279
rect 2222 25276 2228 25288
rect 2179 25248 2228 25276
rect 2179 25245 2191 25248
rect 2133 25239 2191 25245
rect 2222 25236 2228 25248
rect 2280 25236 2286 25288
rect 2501 25279 2559 25285
rect 2501 25245 2513 25279
rect 2547 25245 2559 25279
rect 4706 25276 4712 25288
rect 4667 25248 4712 25276
rect 2501 25239 2559 25245
rect 2406 25168 2412 25220
rect 2464 25208 2470 25220
rect 2516 25208 2544 25239
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 2464 25180 2544 25208
rect 6917 25211 6975 25217
rect 2464 25168 2470 25180
rect 6917 25177 6929 25211
rect 6963 25208 6975 25211
rect 8202 25208 8208 25220
rect 6963 25180 8208 25208
rect 6963 25177 6975 25180
rect 6917 25171 6975 25177
rect 8202 25168 8208 25180
rect 8260 25168 8266 25220
rect 9876 25208 9904 25307
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11333 25347 11391 25353
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11422 25344 11428 25356
rect 11379 25316 11428 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 11808 25353 11836 25384
rect 13262 25372 13268 25384
rect 13320 25372 13326 25424
rect 15378 25412 15384 25424
rect 13372 25384 15384 25412
rect 11793 25347 11851 25353
rect 11793 25313 11805 25347
rect 11839 25313 11851 25347
rect 11793 25307 11851 25313
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 13372 25344 13400 25384
rect 15378 25372 15384 25384
rect 15436 25372 15442 25424
rect 17681 25415 17739 25421
rect 17681 25381 17693 25415
rect 17727 25412 17739 25415
rect 17954 25412 17960 25424
rect 17727 25384 17960 25412
rect 17727 25381 17739 25384
rect 17681 25375 17739 25381
rect 17954 25372 17960 25384
rect 18012 25372 18018 25424
rect 12023 25316 13400 25344
rect 13449 25347 13507 25353
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 13449 25313 13461 25347
rect 13495 25344 13507 25347
rect 13630 25344 13636 25356
rect 13495 25316 13636 25344
rect 13495 25313 13507 25316
rect 13449 25307 13507 25313
rect 13464 25208 13492 25307
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 16022 25344 16028 25356
rect 15983 25316 16028 25344
rect 16022 25304 16028 25316
rect 16080 25304 16086 25356
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 15838 25276 15844 25288
rect 15436 25248 15844 25276
rect 15436 25236 15442 25248
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 16298 25276 16304 25288
rect 16259 25248 16304 25276
rect 16298 25236 16304 25248
rect 16356 25236 16362 25288
rect 9876 25180 13492 25208
rect 7374 25100 7380 25152
rect 7432 25140 7438 25152
rect 8665 25143 8723 25149
rect 8665 25140 8677 25143
rect 7432 25112 8677 25140
rect 7432 25100 7438 25112
rect 8665 25109 8677 25112
rect 8711 25109 8723 25143
rect 8665 25103 8723 25109
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 13541 25143 13599 25149
rect 13541 25140 13553 25143
rect 11112 25112 13553 25140
rect 11112 25100 11118 25112
rect 13541 25109 13553 25112
rect 13587 25109 13599 25143
rect 13541 25103 13599 25109
rect 1104 25050 24840 25072
rect 1104 24998 4947 25050
rect 4999 24998 5011 25050
rect 5063 24998 5075 25050
rect 5127 24998 5139 25050
rect 5191 24998 12878 25050
rect 12930 24998 12942 25050
rect 12994 24998 13006 25050
rect 13058 24998 13070 25050
rect 13122 24998 20808 25050
rect 20860 24998 20872 25050
rect 20924 24998 20936 25050
rect 20988 24998 21000 25050
rect 21052 24998 24840 25050
rect 1104 24976 24840 24998
rect 4706 24936 4712 24948
rect 4667 24908 4712 24936
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 17494 24936 17500 24948
rect 4816 24908 17500 24936
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 4816 24868 4844 24908
rect 17494 24896 17500 24908
rect 17552 24896 17558 24948
rect 4120 24840 4844 24868
rect 4120 24828 4126 24840
rect 5718 24828 5724 24880
rect 5776 24828 5782 24880
rect 5810 24828 5816 24880
rect 5868 24868 5874 24880
rect 9033 24871 9091 24877
rect 9033 24868 9045 24871
rect 5868 24840 9045 24868
rect 5868 24828 5874 24840
rect 9033 24837 9045 24840
rect 9079 24837 9091 24871
rect 9033 24831 9091 24837
rect 9858 24828 9864 24880
rect 9916 24868 9922 24880
rect 10597 24871 10655 24877
rect 10597 24868 10609 24871
rect 9916 24840 10609 24868
rect 9916 24828 9922 24840
rect 10597 24837 10609 24840
rect 10643 24868 10655 24871
rect 11882 24868 11888 24880
rect 10643 24840 11888 24868
rect 10643 24837 10655 24840
rect 10597 24831 10655 24837
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 15930 24828 15936 24880
rect 15988 24868 15994 24880
rect 16761 24871 16819 24877
rect 16761 24868 16773 24871
rect 15988 24840 16773 24868
rect 15988 24828 15994 24840
rect 16761 24837 16773 24840
rect 16807 24837 16819 24871
rect 16761 24831 16819 24837
rect 2682 24800 2688 24812
rect 2643 24772 2688 24800
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 5736 24800 5764 24828
rect 7742 24800 7748 24812
rect 3712 24772 3924 24800
rect 5736 24772 7328 24800
rect 7703 24772 7748 24800
rect 2314 24732 2320 24744
rect 2275 24704 2320 24732
rect 2314 24692 2320 24704
rect 2372 24692 2378 24744
rect 2406 24692 2412 24744
rect 2464 24692 2470 24744
rect 3510 24732 3516 24744
rect 3471 24704 3516 24732
rect 3510 24692 3516 24704
rect 3568 24692 3574 24744
rect 3712 24741 3740 24772
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3896 24732 3924 24772
rect 4062 24732 4068 24744
rect 3896 24704 4068 24732
rect 3697 24695 3755 24701
rect 4062 24692 4068 24704
rect 4120 24732 4126 24744
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 4120 24704 4261 24732
rect 4120 24692 4126 24704
rect 4249 24701 4261 24704
rect 4295 24701 4307 24735
rect 4249 24695 4307 24701
rect 4338 24692 4344 24744
rect 4396 24732 4402 24744
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 4396 24704 4445 24732
rect 4396 24692 4402 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 5721 24735 5779 24741
rect 5721 24701 5733 24735
rect 5767 24732 5779 24735
rect 7006 24732 7012 24744
rect 5767 24704 7012 24732
rect 5767 24701 5779 24704
rect 5721 24695 5779 24701
rect 7006 24692 7012 24704
rect 7064 24732 7070 24744
rect 7190 24732 7196 24744
rect 7064 24704 7196 24732
rect 7064 24692 7070 24704
rect 7190 24692 7196 24704
rect 7248 24692 7254 24744
rect 7300 24741 7328 24772
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 7834 24760 7840 24812
rect 7892 24800 7898 24812
rect 10410 24800 10416 24812
rect 7892 24772 10416 24800
rect 7892 24760 7898 24772
rect 10410 24760 10416 24772
rect 10468 24760 10474 24812
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 11425 24803 11483 24809
rect 11425 24800 11437 24803
rect 10744 24772 11437 24800
rect 10744 24760 10750 24772
rect 11425 24769 11437 24772
rect 11471 24769 11483 24803
rect 11425 24763 11483 24769
rect 11532 24772 18092 24800
rect 7285 24735 7343 24741
rect 7285 24701 7297 24735
rect 7331 24701 7343 24735
rect 7285 24695 7343 24701
rect 7469 24735 7527 24741
rect 7469 24701 7481 24735
rect 7515 24732 7527 24735
rect 8570 24732 8576 24744
rect 7515 24704 8576 24732
rect 7515 24701 7527 24704
rect 7469 24695 7527 24701
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 10870 24692 10876 24744
rect 10928 24732 10934 24744
rect 10962 24735 11020 24741
rect 10962 24732 10974 24735
rect 10928 24704 10974 24732
rect 10928 24692 10934 24704
rect 10962 24701 10974 24704
rect 11008 24701 11020 24735
rect 10962 24695 11020 24701
rect 11149 24735 11207 24741
rect 11149 24701 11161 24735
rect 11195 24701 11207 24735
rect 11149 24695 11207 24701
rect 2133 24667 2191 24673
rect 2133 24633 2145 24667
rect 2179 24664 2191 24667
rect 2424 24664 2452 24692
rect 2179 24636 2452 24664
rect 9127 24667 9185 24673
rect 2179 24633 2191 24636
rect 2133 24627 2191 24633
rect 9127 24633 9139 24667
rect 9173 24633 9185 24667
rect 9127 24627 9185 24633
rect 5813 24599 5871 24605
rect 5813 24565 5825 24599
rect 5859 24596 5871 24599
rect 7834 24596 7840 24608
rect 5859 24568 7840 24596
rect 5859 24565 5871 24568
rect 5813 24559 5871 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 9033 24599 9091 24605
rect 9033 24565 9045 24599
rect 9079 24596 9091 24599
rect 9140 24596 9168 24627
rect 9214 24624 9220 24676
rect 9272 24624 9278 24676
rect 11164 24664 11192 24695
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 11532 24732 11560 24772
rect 12618 24732 12624 24744
rect 11388 24704 11560 24732
rect 12579 24704 12624 24732
rect 11388 24692 11394 24704
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 14093 24735 14151 24741
rect 14093 24701 14105 24735
rect 14139 24732 14151 24735
rect 14182 24732 14188 24744
rect 14139 24704 14188 24732
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24732 14427 24735
rect 14642 24732 14648 24744
rect 14415 24704 14648 24732
rect 14415 24701 14427 24704
rect 14369 24695 14427 24701
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 18064 24741 18092 24772
rect 16577 24735 16635 24741
rect 16577 24732 16589 24735
rect 14792 24704 16589 24732
rect 14792 24692 14798 24704
rect 16577 24701 16589 24704
rect 16623 24701 16635 24735
rect 16577 24695 16635 24701
rect 18049 24735 18107 24741
rect 18049 24701 18061 24735
rect 18095 24701 18107 24735
rect 19150 24732 19156 24744
rect 19111 24704 19156 24732
rect 18049 24695 18107 24701
rect 19150 24692 19156 24704
rect 19208 24692 19214 24744
rect 9416 24636 11192 24664
rect 12437 24667 12495 24673
rect 9079 24568 9168 24596
rect 9232 24596 9260 24624
rect 9416 24596 9444 24636
rect 12437 24633 12449 24667
rect 12483 24664 12495 24667
rect 13446 24664 13452 24676
rect 12483 24636 13452 24664
rect 12483 24633 12495 24636
rect 12437 24627 12495 24633
rect 13446 24624 13452 24636
rect 13504 24624 13510 24676
rect 15749 24667 15807 24673
rect 15749 24633 15761 24667
rect 15795 24664 15807 24667
rect 16482 24664 16488 24676
rect 15795 24636 16488 24664
rect 15795 24633 15807 24636
rect 15749 24627 15807 24633
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 17586 24624 17592 24676
rect 17644 24664 17650 24676
rect 19245 24667 19303 24673
rect 19245 24664 19257 24667
rect 17644 24636 19257 24664
rect 17644 24624 17650 24636
rect 19245 24633 19257 24636
rect 19291 24633 19303 24667
rect 19245 24627 19303 24633
rect 9232 24568 9444 24596
rect 9079 24565 9091 24568
rect 9033 24559 9091 24565
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10226 24596 10232 24608
rect 10008 24568 10232 24596
rect 10008 24556 10014 24568
rect 10226 24556 10232 24568
rect 10284 24556 10290 24608
rect 11422 24556 11428 24608
rect 11480 24596 11486 24608
rect 12713 24599 12771 24605
rect 12713 24596 12725 24599
rect 11480 24568 12725 24596
rect 11480 24556 11486 24568
rect 12713 24565 12725 24568
rect 12759 24565 12771 24599
rect 18230 24596 18236 24608
rect 18191 24568 18236 24596
rect 12713 24559 12771 24565
rect 18230 24556 18236 24568
rect 18288 24556 18294 24608
rect 1104 24506 24840 24528
rect 1104 24454 8912 24506
rect 8964 24454 8976 24506
rect 9028 24454 9040 24506
rect 9092 24454 9104 24506
rect 9156 24454 16843 24506
rect 16895 24454 16907 24506
rect 16959 24454 16971 24506
rect 17023 24454 17035 24506
rect 17087 24454 24840 24506
rect 1104 24432 24840 24454
rect 1489 24395 1547 24401
rect 1489 24361 1501 24395
rect 1535 24392 1547 24395
rect 1762 24392 1768 24404
rect 1535 24364 1768 24392
rect 1535 24361 1547 24364
rect 1489 24355 1547 24361
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 6914 24392 6920 24404
rect 5592 24364 6920 24392
rect 5592 24352 5598 24364
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 8665 24395 8723 24401
rect 8665 24392 8677 24395
rect 8628 24364 8677 24392
rect 8628 24352 8634 24364
rect 8665 24361 8677 24364
rect 8711 24392 8723 24395
rect 9214 24392 9220 24404
rect 8711 24364 9220 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 9214 24352 9220 24364
rect 9272 24352 9278 24404
rect 9692 24364 15976 24392
rect 9692 24336 9720 24364
rect 2682 24324 2688 24336
rect 1412 24296 2688 24324
rect 1412 24265 1440 24296
rect 2682 24284 2688 24296
rect 2740 24284 2746 24336
rect 6273 24327 6331 24333
rect 6273 24293 6285 24327
rect 6319 24324 6331 24327
rect 9674 24324 9680 24336
rect 6319 24296 9680 24324
rect 6319 24293 6331 24296
rect 6273 24287 6331 24293
rect 9674 24284 9680 24296
rect 9732 24284 9738 24336
rect 9861 24327 9919 24333
rect 9861 24293 9873 24327
rect 9907 24324 9919 24327
rect 10134 24324 10140 24336
rect 9907 24296 10140 24324
rect 9907 24293 9919 24296
rect 9861 24287 9919 24293
rect 10134 24284 10140 24296
rect 10192 24284 10198 24336
rect 10505 24327 10563 24333
rect 10505 24293 10517 24327
rect 10551 24324 10563 24327
rect 11882 24324 11888 24336
rect 10551 24296 11888 24324
rect 10551 24293 10563 24296
rect 10505 24287 10563 24293
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 13633 24327 13691 24333
rect 13633 24293 13645 24327
rect 13679 24324 13691 24327
rect 13722 24324 13728 24336
rect 13679 24296 13728 24324
rect 13679 24293 13691 24296
rect 13633 24287 13691 24293
rect 13722 24284 13728 24296
rect 13780 24324 13786 24336
rect 15948 24324 15976 24364
rect 16298 24352 16304 24404
rect 16356 24392 16362 24404
rect 16485 24395 16543 24401
rect 16485 24392 16497 24395
rect 16356 24364 16497 24392
rect 16356 24352 16362 24364
rect 16485 24361 16497 24364
rect 16531 24361 16543 24395
rect 16485 24355 16543 24361
rect 16592 24364 19564 24392
rect 16592 24324 16620 24364
rect 13780 24296 15424 24324
rect 15948 24296 16620 24324
rect 13780 24284 13786 24296
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24225 1455 24259
rect 1397 24219 1455 24225
rect 2409 24259 2467 24265
rect 2409 24225 2421 24259
rect 2455 24256 2467 24259
rect 2498 24256 2504 24268
rect 2455 24228 2504 24256
rect 2455 24225 2467 24228
rect 2409 24219 2467 24225
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 2590 24216 2596 24268
rect 2648 24256 2654 24268
rect 2648 24228 2693 24256
rect 2648 24216 2654 24228
rect 6914 24216 6920 24268
rect 6972 24256 6978 24268
rect 7101 24259 7159 24265
rect 7101 24256 7113 24259
rect 6972 24228 7113 24256
rect 6972 24216 6978 24228
rect 7101 24225 7113 24228
rect 7147 24225 7159 24259
rect 7101 24219 7159 24225
rect 7285 24259 7343 24265
rect 7285 24225 7297 24259
rect 7331 24256 7343 24259
rect 7374 24256 7380 24268
rect 7331 24228 7380 24256
rect 7331 24225 7343 24228
rect 7285 24219 7343 24225
rect 2130 24148 2136 24200
rect 2188 24188 2194 24200
rect 2608 24188 2636 24216
rect 2188 24160 2636 24188
rect 2188 24148 2194 24160
rect 2682 24148 2688 24200
rect 2740 24188 2746 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 2740 24160 4629 24188
rect 2740 24148 2746 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 5350 24188 5356 24200
rect 4939 24160 5356 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 5350 24148 5356 24160
rect 5408 24148 5414 24200
rect 6822 24148 6828 24200
rect 6880 24188 6886 24200
rect 7300 24188 7328 24219
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 7558 24216 7564 24268
rect 7616 24256 7622 24268
rect 7834 24256 7840 24268
rect 7616 24228 7840 24256
rect 7616 24216 7622 24228
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 8294 24216 8300 24268
rect 8352 24256 8358 24268
rect 8481 24259 8539 24265
rect 8481 24256 8493 24259
rect 8352 24228 8493 24256
rect 8352 24216 8358 24228
rect 8481 24225 8493 24228
rect 8527 24256 8539 24259
rect 8662 24256 8668 24268
rect 8527 24228 8668 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 9953 24259 10011 24265
rect 9953 24225 9965 24259
rect 9999 24225 10011 24259
rect 10686 24256 10692 24268
rect 10647 24228 10692 24256
rect 9953 24219 10011 24225
rect 6880 24160 7328 24188
rect 6880 24148 6886 24160
rect 8018 24148 8024 24200
rect 8076 24188 8082 24200
rect 8202 24188 8208 24200
rect 8076 24160 8208 24188
rect 8076 24148 8082 24160
rect 8202 24148 8208 24160
rect 8260 24188 8266 24200
rect 9968 24188 9996 24219
rect 10686 24216 10692 24228
rect 10744 24216 10750 24268
rect 11238 24216 11244 24268
rect 11296 24256 11302 24268
rect 11422 24256 11428 24268
rect 11296 24228 11428 24256
rect 11296 24216 11302 24228
rect 11422 24216 11428 24228
rect 11480 24216 11486 24268
rect 11974 24256 11980 24268
rect 11935 24228 11980 24256
rect 11974 24216 11980 24228
rect 12032 24216 12038 24268
rect 12066 24216 12072 24268
rect 12124 24256 12130 24268
rect 14734 24256 14740 24268
rect 12124 24228 14740 24256
rect 12124 24216 12130 24228
rect 14734 24216 14740 24228
rect 14792 24216 14798 24268
rect 11054 24188 11060 24200
rect 8260 24160 9720 24188
rect 9968 24160 11060 24188
rect 8260 24148 8266 24160
rect 9692 24064 9720 24160
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 12247 24191 12305 24197
rect 12247 24188 12259 24191
rect 11998 24160 12259 24188
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 11998 24120 12026 24160
rect 12247 24157 12259 24160
rect 12293 24157 12305 24191
rect 12247 24151 12305 24157
rect 13906 24148 13912 24200
rect 13964 24188 13970 24200
rect 14918 24188 14924 24200
rect 13964 24160 14924 24188
rect 13964 24148 13970 24160
rect 14918 24148 14924 24160
rect 14976 24188 14982 24200
rect 15289 24191 15347 24197
rect 15289 24188 15301 24191
rect 14976 24160 15301 24188
rect 14976 24148 14982 24160
rect 15289 24157 15301 24160
rect 15335 24157 15347 24191
rect 15396 24188 15424 24296
rect 16666 24284 16672 24336
rect 16724 24324 16730 24336
rect 17497 24327 17555 24333
rect 17497 24324 17509 24327
rect 16724 24296 17509 24324
rect 16724 24284 16730 24296
rect 17497 24293 17509 24296
rect 17543 24293 17555 24327
rect 17497 24287 17555 24293
rect 17954 24284 17960 24336
rect 18012 24324 18018 24336
rect 18414 24324 18420 24336
rect 18012 24296 18420 24324
rect 18012 24284 18018 24296
rect 18414 24284 18420 24296
rect 18472 24324 18478 24336
rect 18472 24296 18552 24324
rect 18472 24284 18478 24296
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24256 15531 24259
rect 15838 24256 15844 24268
rect 15519 24228 15844 24256
rect 15519 24225 15531 24228
rect 15473 24219 15531 24225
rect 15838 24216 15844 24228
rect 15896 24256 15902 24268
rect 16025 24259 16083 24265
rect 16025 24256 16037 24259
rect 15896 24228 16037 24256
rect 15896 24216 15902 24228
rect 16025 24225 16037 24228
rect 16071 24225 16083 24259
rect 16025 24219 16083 24225
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 17126 24256 17132 24268
rect 16255 24228 17132 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 18138 24256 18144 24268
rect 18099 24228 18144 24256
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18524 24265 18552 24296
rect 19536 24265 19564 24364
rect 18509 24259 18567 24265
rect 18509 24225 18521 24259
rect 18555 24225 18567 24259
rect 18509 24219 18567 24225
rect 19521 24259 19579 24265
rect 19521 24225 19533 24259
rect 19567 24225 19579 24259
rect 19521 24219 19579 24225
rect 15396 24160 15700 24188
rect 15289 24151 15347 24157
rect 11296 24092 12026 24120
rect 15672 24120 15700 24160
rect 16482 24148 16488 24200
rect 16540 24188 16546 24200
rect 18049 24191 18107 24197
rect 18049 24188 18061 24191
rect 16540 24160 18061 24188
rect 16540 24148 16546 24160
rect 18049 24157 18061 24160
rect 18095 24157 18107 24191
rect 18598 24188 18604 24200
rect 18559 24160 18604 24188
rect 18049 24151 18107 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 19150 24120 19156 24132
rect 15672 24092 19156 24120
rect 11296 24080 11302 24092
rect 19150 24080 19156 24092
rect 19208 24080 19214 24132
rect 2406 24012 2412 24064
rect 2464 24052 2470 24064
rect 2685 24055 2743 24061
rect 2685 24052 2697 24055
rect 2464 24024 2697 24052
rect 2464 24012 2470 24024
rect 2685 24021 2697 24024
rect 2731 24021 2743 24055
rect 2685 24015 2743 24021
rect 7006 24012 7012 24064
rect 7064 24052 7070 24064
rect 7377 24055 7435 24061
rect 7377 24052 7389 24055
rect 7064 24024 7389 24052
rect 7064 24012 7070 24024
rect 7377 24021 7389 24024
rect 7423 24021 7435 24055
rect 7377 24015 7435 24021
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 10134 24052 10140 24064
rect 9732 24024 9777 24052
rect 10095 24024 10140 24052
rect 9732 24012 9738 24024
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10594 24012 10600 24064
rect 10652 24052 10658 24064
rect 10781 24055 10839 24061
rect 10781 24052 10793 24055
rect 10652 24024 10793 24052
rect 10652 24012 10658 24024
rect 10781 24021 10793 24024
rect 10827 24021 10839 24055
rect 10781 24015 10839 24021
rect 14366 24012 14372 24064
rect 14424 24052 14430 24064
rect 19613 24055 19671 24061
rect 19613 24052 19625 24055
rect 14424 24024 19625 24052
rect 14424 24012 14430 24024
rect 19613 24021 19625 24024
rect 19659 24021 19671 24055
rect 19613 24015 19671 24021
rect 1104 23962 24840 23984
rect 1104 23910 4947 23962
rect 4999 23910 5011 23962
rect 5063 23910 5075 23962
rect 5127 23910 5139 23962
rect 5191 23910 12878 23962
rect 12930 23910 12942 23962
rect 12994 23910 13006 23962
rect 13058 23910 13070 23962
rect 13122 23910 20808 23962
rect 20860 23910 20872 23962
rect 20924 23910 20936 23962
rect 20988 23910 21000 23962
rect 21052 23910 24840 23962
rect 1104 23888 24840 23910
rect 1302 23808 1308 23860
rect 1360 23848 1366 23860
rect 1360 23820 2268 23848
rect 1360 23808 1366 23820
rect 2130 23740 2136 23792
rect 2188 23740 2194 23792
rect 2240 23780 2268 23820
rect 2498 23808 2504 23860
rect 2556 23848 2562 23860
rect 2682 23848 2688 23860
rect 2556 23820 2688 23848
rect 2556 23808 2562 23820
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 7098 23808 7104 23860
rect 7156 23848 7162 23860
rect 8665 23851 8723 23857
rect 8665 23848 8677 23851
rect 7156 23820 8677 23848
rect 7156 23808 7162 23820
rect 8665 23817 8677 23820
rect 8711 23817 8723 23851
rect 8665 23811 8723 23817
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 10781 23851 10839 23857
rect 10781 23848 10793 23851
rect 10744 23820 10793 23848
rect 10744 23808 10750 23820
rect 10781 23817 10793 23820
rect 10827 23817 10839 23851
rect 10781 23811 10839 23817
rect 11790 23808 11796 23860
rect 11848 23848 11854 23860
rect 18506 23848 18512 23860
rect 11848 23820 18512 23848
rect 11848 23808 11854 23820
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 5810 23780 5816 23792
rect 2240 23752 5816 23780
rect 5810 23740 5816 23752
rect 5868 23740 5874 23792
rect 14366 23780 14372 23792
rect 7300 23752 14372 23780
rect 2148 23712 2176 23740
rect 2682 23712 2688 23724
rect 2148 23684 2688 23712
rect 1762 23604 1768 23656
rect 1820 23644 1826 23656
rect 2133 23647 2191 23653
rect 2133 23644 2145 23647
rect 1820 23616 2145 23644
rect 1820 23604 1826 23616
rect 2133 23613 2145 23616
rect 2179 23613 2191 23647
rect 2133 23607 2191 23613
rect 2222 23604 2228 23656
rect 2280 23644 2286 23656
rect 2516 23653 2544 23684
rect 2682 23672 2688 23684
rect 2740 23672 2746 23724
rect 4246 23712 4252 23724
rect 4207 23684 4252 23712
rect 4246 23672 4252 23684
rect 4304 23672 4310 23724
rect 4338 23672 4344 23724
rect 4396 23712 4402 23724
rect 5077 23715 5135 23721
rect 5077 23712 5089 23715
rect 4396 23684 5089 23712
rect 4396 23672 4402 23684
rect 5077 23681 5089 23684
rect 5123 23681 5135 23715
rect 5077 23675 5135 23681
rect 2501 23647 2559 23653
rect 2280 23616 2325 23644
rect 2280 23604 2286 23616
rect 2501 23613 2513 23647
rect 2547 23613 2559 23647
rect 2501 23607 2559 23613
rect 2590 23604 2596 23656
rect 2648 23644 2654 23656
rect 4617 23647 4675 23653
rect 2648 23616 2693 23644
rect 2648 23604 2654 23616
rect 4617 23613 4629 23647
rect 4663 23613 4675 23647
rect 4617 23607 4675 23613
rect 1489 23579 1547 23585
rect 1489 23545 1501 23579
rect 1535 23576 1547 23579
rect 1670 23576 1676 23588
rect 1535 23548 1676 23576
rect 1535 23545 1547 23548
rect 1489 23539 1547 23545
rect 1670 23536 1676 23548
rect 1728 23536 1734 23588
rect 4632 23576 4660 23607
rect 4706 23604 4712 23656
rect 4764 23644 4770 23656
rect 4801 23647 4859 23653
rect 4801 23644 4813 23647
rect 4764 23616 4813 23644
rect 4764 23604 4770 23616
rect 4801 23613 4813 23616
rect 4847 23613 4859 23647
rect 4801 23607 4859 23613
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23644 5227 23647
rect 5534 23644 5540 23656
rect 5215 23616 5540 23644
rect 5215 23613 5227 23616
rect 5169 23607 5227 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 5810 23604 5816 23656
rect 5868 23644 5874 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 5868 23616 6837 23644
rect 5868 23604 5874 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 7006 23644 7012 23656
rect 6967 23616 7012 23644
rect 6825 23607 6883 23613
rect 7006 23604 7012 23616
rect 7064 23604 7070 23656
rect 7098 23604 7104 23656
rect 7156 23644 7162 23656
rect 7156 23616 7201 23644
rect 7156 23604 7162 23616
rect 4982 23576 4988 23588
rect 4632 23548 4988 23576
rect 4982 23536 4988 23548
rect 5040 23576 5046 23588
rect 7300 23576 7328 23752
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 14642 23780 14648 23792
rect 14603 23752 14648 23780
rect 14642 23740 14648 23752
rect 14700 23740 14706 23792
rect 15102 23740 15108 23792
rect 15160 23780 15166 23792
rect 16482 23780 16488 23792
rect 15160 23752 16488 23780
rect 15160 23740 15166 23752
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23749 18291 23783
rect 18233 23743 18291 23749
rect 19337 23783 19395 23789
rect 19337 23749 19349 23783
rect 19383 23749 19395 23783
rect 19337 23743 19395 23749
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23712 10379 23715
rect 10870 23712 10876 23724
rect 10367 23684 10876 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 10870 23672 10876 23684
rect 10928 23712 10934 23724
rect 11146 23712 11152 23724
rect 10928 23684 11152 23712
rect 10928 23672 10934 23684
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 11606 23672 11612 23724
rect 11664 23712 11670 23724
rect 13633 23715 13691 23721
rect 11664 23684 12480 23712
rect 11664 23672 11670 23684
rect 8573 23647 8631 23653
rect 8573 23613 8585 23647
rect 8619 23644 8631 23647
rect 8662 23644 8668 23656
rect 8619 23616 8668 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 8662 23604 8668 23616
rect 8720 23644 8726 23656
rect 9490 23644 9496 23656
rect 8720 23616 9496 23644
rect 8720 23604 8726 23616
rect 9490 23604 9496 23616
rect 9548 23604 9554 23656
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23644 10655 23647
rect 12342 23644 12348 23656
rect 10643 23616 12348 23644
rect 10643 23613 10655 23616
rect 10597 23607 10655 23613
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12452 23653 12480 23684
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13906 23712 13912 23724
rect 13679 23684 13912 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 15746 23712 15752 23724
rect 15707 23684 15752 23712
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 16206 23712 16212 23724
rect 16167 23684 16212 23712
rect 16206 23672 16212 23684
rect 16264 23672 16270 23724
rect 18248 23712 18276 23743
rect 16776 23684 18276 23712
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23613 12495 23647
rect 13722 23644 13728 23656
rect 13635 23616 13728 23644
rect 12437 23607 12495 23613
rect 13722 23604 13728 23616
rect 13780 23644 13786 23656
rect 14277 23647 14335 23653
rect 14277 23644 14289 23647
rect 13780 23616 14289 23644
rect 13780 23604 13786 23616
rect 14277 23613 14289 23616
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 14461 23647 14519 23653
rect 14461 23613 14473 23647
rect 14507 23644 14519 23647
rect 16224 23644 16252 23672
rect 14507 23616 16252 23644
rect 16393 23647 16451 23653
rect 14507 23613 14519 23616
rect 14461 23607 14519 23613
rect 16393 23613 16405 23647
rect 16439 23644 16451 23647
rect 16482 23644 16488 23656
rect 16439 23616 16488 23644
rect 16439 23613 16451 23616
rect 16393 23607 16451 23613
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 16776 23653 16804 23684
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18380 23684 19288 23712
rect 18380 23672 18386 23684
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16724 23616 16773 23644
rect 16724 23604 16730 23616
rect 16761 23613 16773 23616
rect 16807 23613 16819 23647
rect 16761 23607 16819 23613
rect 16945 23647 17003 23653
rect 16945 23613 16957 23647
rect 16991 23644 17003 23647
rect 17126 23644 17132 23656
rect 16991 23616 17132 23644
rect 16991 23613 17003 23616
rect 16945 23607 17003 23613
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18506 23604 18512 23656
rect 18564 23644 18570 23656
rect 19141 23647 19199 23653
rect 19141 23644 19153 23647
rect 18564 23616 19153 23644
rect 18564 23604 18570 23616
rect 19141 23613 19153 23616
rect 19187 23613 19199 23647
rect 19260 23644 19288 23684
rect 19352 23644 19380 23743
rect 19260 23616 19380 23644
rect 20257 23647 20315 23653
rect 19141 23607 19199 23613
rect 20257 23613 20269 23647
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 5040 23548 7328 23576
rect 5040 23536 5046 23548
rect 7374 23536 7380 23588
rect 7432 23576 7438 23588
rect 7561 23579 7619 23585
rect 7561 23576 7573 23579
rect 7432 23548 7573 23576
rect 7432 23536 7438 23548
rect 7561 23545 7573 23548
rect 7607 23545 7619 23579
rect 7561 23539 7619 23545
rect 8389 23579 8447 23585
rect 8389 23545 8401 23579
rect 8435 23576 8447 23579
rect 9214 23576 9220 23588
rect 8435 23548 9220 23576
rect 8435 23545 8447 23548
rect 8389 23539 8447 23545
rect 9214 23536 9220 23548
rect 9272 23536 9278 23588
rect 10505 23579 10563 23585
rect 10505 23545 10517 23579
rect 10551 23576 10563 23579
rect 13078 23576 13084 23588
rect 10551 23548 13084 23576
rect 10551 23545 10563 23548
rect 10505 23539 10563 23545
rect 13078 23536 13084 23548
rect 13136 23536 13142 23588
rect 14550 23536 14556 23588
rect 14608 23576 14614 23588
rect 15102 23576 15108 23588
rect 14608 23548 15108 23576
rect 14608 23536 14614 23548
rect 15102 23536 15108 23548
rect 15160 23536 15166 23588
rect 18414 23536 18420 23588
rect 18472 23576 18478 23588
rect 20272 23576 20300 23607
rect 18472 23548 20300 23576
rect 18472 23536 18478 23548
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 3786 23508 3792 23520
rect 3568 23480 3792 23508
rect 3568 23468 3574 23480
rect 3786 23468 3792 23480
rect 3844 23468 3850 23520
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 7282 23508 7288 23520
rect 7064 23480 7288 23508
rect 7064 23468 7070 23480
rect 7282 23468 7288 23480
rect 7340 23468 7346 23520
rect 8294 23468 8300 23520
rect 8352 23508 8358 23520
rect 11790 23508 11796 23520
rect 8352 23480 11796 23508
rect 8352 23468 8358 23480
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 11882 23468 11888 23520
rect 11940 23508 11946 23520
rect 12342 23508 12348 23520
rect 11940 23480 12348 23508
rect 11940 23468 11946 23480
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 12618 23508 12624 23520
rect 12579 23480 12624 23508
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 13814 23508 13820 23520
rect 13412 23480 13820 23508
rect 13412 23468 13418 23480
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 17586 23508 17592 23520
rect 13872 23480 17592 23508
rect 13872 23468 13878 23480
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 17862 23468 17868 23520
rect 17920 23508 17926 23520
rect 20349 23511 20407 23517
rect 20349 23508 20361 23511
rect 17920 23480 20361 23508
rect 17920 23468 17926 23480
rect 20349 23477 20361 23480
rect 20395 23477 20407 23511
rect 20349 23471 20407 23477
rect 1104 23418 24840 23440
rect 1104 23366 8912 23418
rect 8964 23366 8976 23418
rect 9028 23366 9040 23418
rect 9092 23366 9104 23418
rect 9156 23366 16843 23418
rect 16895 23366 16907 23418
rect 16959 23366 16971 23418
rect 17023 23366 17035 23418
rect 17087 23366 24840 23418
rect 1104 23344 24840 23366
rect 2682 23264 2688 23316
rect 2740 23304 2746 23316
rect 2777 23307 2835 23313
rect 2777 23304 2789 23307
rect 2740 23276 2789 23304
rect 2740 23264 2746 23276
rect 2777 23273 2789 23276
rect 2823 23273 2835 23307
rect 2777 23267 2835 23273
rect 4062 23264 4068 23316
rect 4120 23264 4126 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 8352 23276 8493 23304
rect 8352 23264 8358 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 11790 23304 11796 23316
rect 8481 23267 8539 23273
rect 9968 23276 11796 23304
rect 1670 23168 1676 23180
rect 1631 23140 1676 23168
rect 1670 23128 1676 23140
rect 1728 23128 1734 23180
rect 3878 23128 3884 23180
rect 3936 23168 3942 23180
rect 4080 23168 4108 23264
rect 5350 23236 5356 23248
rect 5311 23208 5356 23236
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 9490 23196 9496 23248
rect 9548 23236 9554 23248
rect 9858 23236 9864 23248
rect 9548 23208 9864 23236
rect 9548 23196 9554 23208
rect 9858 23196 9864 23208
rect 9916 23196 9922 23248
rect 9968 23245 9996 23276
rect 11790 23264 11796 23276
rect 11848 23264 11854 23316
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 12529 23307 12587 23313
rect 12529 23304 12541 23307
rect 12308 23276 12541 23304
rect 12308 23264 12314 23276
rect 12529 23273 12541 23276
rect 12575 23273 12587 23307
rect 12529 23267 12587 23273
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 13817 23307 13875 23313
rect 13817 23304 13829 23307
rect 13136 23276 13829 23304
rect 13136 23264 13142 23276
rect 13817 23273 13829 23276
rect 13863 23273 13875 23307
rect 15565 23307 15623 23313
rect 15565 23304 15577 23307
rect 13817 23267 13875 23273
rect 13924 23276 15577 23304
rect 9953 23239 10011 23245
rect 9953 23205 9965 23239
rect 9999 23205 10011 23239
rect 11882 23236 11888 23248
rect 9953 23199 10011 23205
rect 11624 23208 11888 23236
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 3936 23140 4261 23168
rect 3936 23128 3942 23140
rect 4249 23137 4261 23140
rect 4295 23168 4307 23171
rect 4801 23171 4859 23177
rect 4801 23168 4813 23171
rect 4295 23140 4813 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4801 23137 4813 23140
rect 4847 23137 4859 23171
rect 4982 23168 4988 23180
rect 4943 23140 4988 23168
rect 4801 23131 4859 23137
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 7374 23168 7380 23180
rect 7335 23140 7380 23168
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 10134 23168 10140 23180
rect 10095 23140 10140 23168
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 11422 23128 11428 23180
rect 11480 23168 11486 23180
rect 11624 23177 11652 23208
rect 11882 23196 11888 23208
rect 11940 23196 11946 23248
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 13924 23236 13952 23276
rect 15565 23273 15577 23276
rect 15611 23273 15623 23307
rect 15565 23267 15623 23273
rect 16482 23264 16488 23316
rect 16540 23304 16546 23316
rect 18417 23307 18475 23313
rect 18417 23304 18429 23307
rect 16540 23276 18429 23304
rect 16540 23264 16546 23276
rect 18417 23273 18429 23276
rect 18463 23273 18475 23307
rect 18417 23267 18475 23273
rect 12492 23208 13952 23236
rect 15289 23239 15347 23245
rect 12492 23196 12498 23208
rect 15289 23205 15301 23239
rect 15335 23236 15347 23239
rect 16574 23236 16580 23248
rect 15335 23208 16580 23236
rect 15335 23205 15347 23208
rect 15289 23199 15347 23205
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 17405 23239 17463 23245
rect 16868 23208 17080 23236
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 11480 23140 11529 23168
rect 11480 23128 11486 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 11517 23131 11575 23137
rect 11609 23171 11667 23177
rect 11609 23137 11621 23171
rect 11655 23137 11667 23171
rect 11983 23171 12041 23177
rect 11983 23168 11995 23171
rect 11609 23131 11667 23137
rect 11716 23140 11995 23168
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23100 1455 23103
rect 2498 23100 2504 23112
rect 1443 23072 2504 23100
rect 1443 23069 1455 23072
rect 1397 23063 1455 23069
rect 2498 23060 2504 23072
rect 2556 23060 2562 23112
rect 4154 23100 4160 23112
rect 4115 23072 4160 23100
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 5902 23060 5908 23112
rect 5960 23100 5966 23112
rect 7101 23103 7159 23109
rect 7101 23100 7113 23103
rect 5960 23072 7113 23100
rect 5960 23060 5966 23072
rect 7101 23069 7113 23072
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 11716 23032 11744 23140
rect 11983 23137 11995 23140
rect 12029 23137 12041 23171
rect 11983 23131 12041 23137
rect 12069 23171 12127 23177
rect 12069 23137 12081 23171
rect 12115 23168 12127 23171
rect 12250 23168 12256 23180
rect 12115 23140 12256 23168
rect 12115 23137 12127 23140
rect 12069 23131 12127 23137
rect 12250 23128 12256 23140
rect 12308 23128 12314 23180
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 16868 23177 16896 23208
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23137 13783 23171
rect 15473 23171 15531 23177
rect 15473 23168 15485 23171
rect 13725 23131 13783 23137
rect 13813 23140 15485 23168
rect 12710 23060 12716 23112
rect 12768 23100 12774 23112
rect 13740 23100 13768 23131
rect 12768 23072 13768 23100
rect 12768 23060 12774 23072
rect 13354 23032 13360 23044
rect 11716 23004 13360 23032
rect 13354 22992 13360 23004
rect 13412 22992 13418 23044
rect 13446 22992 13452 23044
rect 13504 23032 13510 23044
rect 13630 23032 13636 23044
rect 13504 23004 13636 23032
rect 13504 22992 13510 23004
rect 13630 22992 13636 23004
rect 13688 23032 13694 23044
rect 13813 23032 13841 23140
rect 15473 23137 15485 23140
rect 15519 23168 15531 23171
rect 16669 23171 16727 23177
rect 16669 23168 16681 23171
rect 15519 23140 16681 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 16669 23137 16681 23140
rect 16715 23137 16727 23171
rect 16669 23131 16727 23137
rect 16853 23171 16911 23177
rect 16853 23137 16865 23171
rect 16899 23137 16911 23171
rect 16853 23131 16911 23137
rect 16945 23171 17003 23177
rect 16945 23137 16957 23171
rect 16991 23137 17003 23171
rect 17052 23168 17080 23208
rect 17405 23205 17417 23239
rect 17451 23236 17463 23239
rect 18138 23236 18144 23248
rect 17451 23208 18144 23236
rect 17451 23205 17463 23208
rect 17405 23199 17463 23205
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 17126 23168 17132 23180
rect 17039 23140 17132 23168
rect 16945 23131 17003 23137
rect 16960 23100 16988 23131
rect 17126 23128 17132 23140
rect 17184 23168 17190 23180
rect 17862 23168 17868 23180
rect 17184 23140 17868 23168
rect 17184 23128 17190 23140
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18233 23171 18291 23177
rect 18233 23168 18245 23171
rect 18012 23140 18245 23168
rect 18012 23128 18018 23140
rect 18233 23137 18245 23140
rect 18279 23168 18291 23171
rect 18690 23168 18696 23180
rect 18279 23140 18696 23168
rect 18279 23137 18291 23140
rect 18233 23131 18291 23137
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 19337 23171 19395 23177
rect 19337 23137 19349 23171
rect 19383 23137 19395 23171
rect 19337 23131 19395 23137
rect 19242 23100 19248 23112
rect 16960 23072 19248 23100
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 13688 23004 13841 23032
rect 13688 22992 13694 23004
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 19352 23032 19380 23131
rect 15252 23004 19380 23032
rect 15252 22992 15258 23004
rect 1854 22924 1860 22976
rect 1912 22964 1918 22976
rect 7558 22964 7564 22976
rect 1912 22936 7564 22964
rect 1912 22924 1918 22936
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10229 22967 10287 22973
rect 10229 22964 10241 22967
rect 10008 22936 10241 22964
rect 10008 22924 10014 22936
rect 10229 22933 10241 22936
rect 10275 22933 10287 22967
rect 10229 22927 10287 22933
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 18230 22964 18236 22976
rect 16715 22936 18236 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19521 22967 19579 22973
rect 19521 22964 19533 22967
rect 19484 22936 19533 22964
rect 19484 22924 19490 22936
rect 19521 22933 19533 22936
rect 19567 22933 19579 22967
rect 19521 22927 19579 22933
rect 1104 22874 24840 22896
rect 1104 22822 4947 22874
rect 4999 22822 5011 22874
rect 5063 22822 5075 22874
rect 5127 22822 5139 22874
rect 5191 22822 12878 22874
rect 12930 22822 12942 22874
rect 12994 22822 13006 22874
rect 13058 22822 13070 22874
rect 13122 22822 20808 22874
rect 20860 22822 20872 22874
rect 20924 22822 20936 22874
rect 20988 22822 21000 22874
rect 21052 22822 24840 22874
rect 1104 22800 24840 22822
rect 1854 22760 1860 22772
rect 1815 22732 1860 22760
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 2915 22763 2973 22769
rect 2915 22760 2927 22763
rect 2740 22732 2927 22760
rect 2740 22720 2746 22732
rect 2915 22729 2927 22732
rect 2961 22729 2973 22763
rect 2915 22723 2973 22729
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 7156 22732 8493 22760
rect 7156 22720 7162 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 11698 22760 11704 22772
rect 8481 22723 8539 22729
rect 9600 22732 11704 22760
rect 2314 22652 2320 22704
rect 2372 22692 2378 22704
rect 3053 22695 3111 22701
rect 3053 22692 3065 22695
rect 2372 22664 3065 22692
rect 2372 22652 2378 22664
rect 3053 22661 3065 22664
rect 3099 22661 3111 22695
rect 3053 22655 3111 22661
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 4430 22692 4436 22704
rect 4120 22664 4436 22692
rect 4120 22652 4126 22664
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 4706 22652 4712 22704
rect 4764 22692 4770 22704
rect 4982 22692 4988 22704
rect 4764 22664 4988 22692
rect 4764 22652 4770 22664
rect 4982 22652 4988 22664
rect 5040 22692 5046 22704
rect 5040 22664 8340 22692
rect 5040 22652 5046 22664
rect 3142 22584 3148 22636
rect 3200 22624 3206 22636
rect 4893 22627 4951 22633
rect 3200 22596 3245 22624
rect 3200 22584 3206 22596
rect 4893 22593 4905 22627
rect 4939 22624 4951 22627
rect 7926 22624 7932 22636
rect 4939 22596 7932 22624
rect 4939 22593 4951 22596
rect 4893 22587 4951 22593
rect 7926 22584 7932 22596
rect 7984 22624 7990 22636
rect 7984 22596 8248 22624
rect 7984 22584 7990 22596
rect 1670 22556 1676 22568
rect 1631 22528 1676 22556
rect 1670 22516 1676 22528
rect 1728 22516 1734 22568
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 5445 22559 5503 22565
rect 5445 22556 5457 22559
rect 2823 22528 5457 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 5445 22525 5457 22528
rect 5491 22556 5503 22559
rect 5491 22528 5580 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 2866 22380 2872 22432
rect 2924 22420 2930 22432
rect 3421 22423 3479 22429
rect 3421 22420 3433 22423
rect 2924 22392 3433 22420
rect 2924 22380 2930 22392
rect 3421 22389 3433 22392
rect 3467 22389 3479 22423
rect 5552 22420 5580 22528
rect 5626 22516 5632 22568
rect 5684 22556 5690 22568
rect 5721 22559 5779 22565
rect 5721 22556 5733 22559
rect 5684 22528 5733 22556
rect 5684 22516 5690 22528
rect 5721 22525 5733 22528
rect 5767 22525 5779 22559
rect 5721 22519 5779 22525
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 6178 22556 6184 22568
rect 5951 22528 6184 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 6178 22516 6184 22528
rect 6236 22516 6242 22568
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 7009 22559 7067 22565
rect 7009 22525 7021 22559
rect 7055 22556 7067 22559
rect 7650 22556 7656 22568
rect 7055 22528 7656 22556
rect 7055 22525 7067 22528
rect 7009 22519 7067 22525
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 8220 22565 8248 22596
rect 8205 22559 8263 22565
rect 8205 22525 8217 22559
rect 8251 22525 8263 22559
rect 8205 22519 8263 22525
rect 7558 22488 7564 22500
rect 6932 22460 7564 22488
rect 6932 22420 6960 22460
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8312 22488 8340 22664
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 8478 22556 8484 22568
rect 8435 22528 8484 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 8478 22516 8484 22528
rect 8536 22516 8542 22568
rect 9600 22565 9628 22732
rect 11698 22720 11704 22732
rect 11756 22720 11762 22772
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 13630 22760 13636 22772
rect 13320 22732 13636 22760
rect 13320 22720 13326 22732
rect 13630 22720 13636 22732
rect 13688 22760 13694 22772
rect 18322 22760 18328 22772
rect 13688 22732 18328 22760
rect 13688 22720 13694 22732
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 19242 22720 19248 22772
rect 19300 22760 19306 22772
rect 19521 22763 19579 22769
rect 19521 22760 19533 22763
rect 19300 22732 19533 22760
rect 19300 22720 19306 22732
rect 19521 22729 19533 22732
rect 19567 22729 19579 22763
rect 19521 22723 19579 22729
rect 10134 22652 10140 22704
rect 10192 22692 10198 22704
rect 13998 22692 14004 22704
rect 10192 22664 14004 22692
rect 10192 22652 10198 22664
rect 13998 22652 14004 22664
rect 14056 22692 14062 22704
rect 15562 22692 15568 22704
rect 14056 22664 15568 22692
rect 14056 22652 14062 22664
rect 15562 22652 15568 22664
rect 15620 22652 15626 22704
rect 16482 22692 16488 22704
rect 16040 22664 16488 22692
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 13170 22624 13176 22636
rect 10827 22596 13176 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 13372 22596 13584 22624
rect 9585 22559 9643 22565
rect 9585 22525 9597 22559
rect 9631 22525 9643 22559
rect 10686 22556 10692 22568
rect 10647 22528 10692 22556
rect 9585 22519 9643 22525
rect 10686 22516 10692 22528
rect 10744 22516 10750 22568
rect 10962 22556 10968 22568
rect 10923 22528 10968 22556
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 11606 22516 11612 22568
rect 11664 22556 11670 22568
rect 11882 22556 11888 22568
rect 11664 22528 11888 22556
rect 11664 22516 11670 22528
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 13372 22565 13400 22596
rect 13357 22559 13415 22565
rect 13357 22525 13369 22559
rect 13403 22525 13415 22559
rect 13357 22519 13415 22525
rect 13449 22559 13507 22565
rect 13449 22525 13461 22559
rect 13495 22525 13507 22559
rect 13556 22556 13584 22596
rect 14826 22584 14832 22636
rect 14884 22624 14890 22636
rect 15381 22627 15439 22633
rect 15381 22624 15393 22627
rect 14884 22596 15393 22624
rect 14884 22584 14890 22596
rect 15381 22593 15393 22596
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 13722 22556 13728 22568
rect 13556 22528 13728 22556
rect 13449 22519 13507 22525
rect 9674 22488 9680 22500
rect 8312 22460 9680 22488
rect 9674 22448 9680 22460
rect 9732 22448 9738 22500
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 10980 22488 11008 22516
rect 10468 22460 11008 22488
rect 13464 22488 13492 22519
rect 13722 22516 13728 22528
rect 13780 22556 13786 22568
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13780 22528 13921 22556
rect 13780 22516 13786 22528
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 14139 22528 15853 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 15841 22525 15853 22528
rect 15887 22525 15899 22559
rect 15841 22519 15899 22525
rect 14734 22488 14740 22500
rect 13464 22460 14740 22488
rect 10468 22448 10474 22460
rect 14734 22448 14740 22460
rect 14792 22448 14798 22500
rect 15856 22488 15884 22519
rect 15930 22516 15936 22568
rect 15988 22556 15994 22568
rect 16040 22565 16068 22664
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 17678 22652 17684 22704
rect 17736 22692 17742 22704
rect 19426 22692 19432 22704
rect 17736 22664 19432 22692
rect 17736 22652 17742 22664
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 16298 22624 16304 22636
rect 16259 22596 16304 22624
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 18598 22624 18604 22636
rect 18559 22596 18604 22624
rect 18598 22584 18604 22596
rect 18656 22624 18662 22636
rect 18656 22596 19472 22624
rect 18656 22584 18662 22596
rect 16025 22559 16083 22565
rect 16025 22556 16037 22559
rect 15988 22528 16037 22556
rect 15988 22516 15994 22528
rect 16025 22525 16037 22528
rect 16071 22525 16083 22559
rect 16025 22519 16083 22525
rect 16393 22559 16451 22565
rect 16393 22525 16405 22559
rect 16439 22556 16451 22559
rect 16666 22556 16672 22568
rect 16439 22528 16672 22556
rect 16439 22525 16451 22528
rect 16393 22519 16451 22525
rect 16666 22516 16672 22528
rect 16724 22556 16730 22568
rect 17126 22556 17132 22568
rect 16724 22528 17132 22556
rect 16724 22516 16730 22528
rect 17126 22516 17132 22528
rect 17184 22516 17190 22568
rect 18230 22556 18236 22568
rect 18191 22528 18236 22556
rect 18230 22516 18236 22528
rect 18288 22516 18294 22568
rect 19444 22565 19472 22596
rect 19429 22559 19487 22565
rect 19429 22525 19441 22559
rect 19475 22525 19487 22559
rect 19429 22519 19487 22525
rect 16574 22488 16580 22500
rect 15856 22460 16580 22488
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 18049 22491 18107 22497
rect 18049 22457 18061 22491
rect 18095 22488 18107 22491
rect 19150 22488 19156 22500
rect 18095 22460 19156 22488
rect 18095 22457 18107 22460
rect 18049 22451 18107 22457
rect 19150 22448 19156 22460
rect 19208 22448 19214 22500
rect 7098 22420 7104 22432
rect 5552 22392 6960 22420
rect 7059 22392 7104 22420
rect 3421 22383 3479 22389
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 9398 22380 9404 22432
rect 9456 22420 9462 22432
rect 9582 22420 9588 22432
rect 9456 22392 9588 22420
rect 9456 22380 9462 22392
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22420 9830 22432
rect 10134 22420 10140 22432
rect 9824 22392 10140 22420
rect 9824 22380 9830 22392
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 11146 22420 11152 22432
rect 11107 22392 11152 22420
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 14366 22420 14372 22432
rect 14327 22392 14372 22420
rect 14366 22380 14372 22392
rect 14424 22380 14430 22432
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 19518 22420 19524 22432
rect 14608 22392 19524 22420
rect 14608 22380 14614 22392
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 1104 22330 24840 22352
rect 1104 22278 8912 22330
rect 8964 22278 8976 22330
rect 9028 22278 9040 22330
rect 9092 22278 9104 22330
rect 9156 22278 16843 22330
rect 16895 22278 16907 22330
rect 16959 22278 16971 22330
rect 17023 22278 17035 22330
rect 17087 22278 24840 22330
rect 1104 22256 24840 22278
rect 8478 22216 8484 22228
rect 6840 22188 8484 22216
rect 6840 22157 6868 22188
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13725 22219 13783 22225
rect 13725 22216 13737 22219
rect 13596 22188 13737 22216
rect 13596 22176 13602 22188
rect 13725 22185 13737 22188
rect 13771 22216 13783 22219
rect 14550 22216 14556 22228
rect 13771 22188 14556 22216
rect 13771 22185 13783 22188
rect 13725 22179 13783 22185
rect 14550 22176 14556 22188
rect 14608 22176 14614 22228
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 17678 22216 17684 22228
rect 15620 22188 17684 22216
rect 15620 22176 15626 22188
rect 17678 22176 17684 22188
rect 17736 22176 17742 22228
rect 6825 22151 6883 22157
rect 6825 22117 6837 22151
rect 6871 22117 6883 22151
rect 6825 22111 6883 22117
rect 7190 22108 7196 22160
rect 7248 22148 7254 22160
rect 10781 22151 10839 22157
rect 7248 22120 8340 22148
rect 7248 22108 7254 22120
rect 1765 22083 1823 22089
rect 1765 22049 1777 22083
rect 1811 22080 1823 22083
rect 2314 22080 2320 22092
rect 1811 22052 2320 22080
rect 1811 22049 1823 22052
rect 1765 22043 1823 22049
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2869 22083 2927 22089
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 4893 22083 4951 22089
rect 2915 22052 4568 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 4062 21972 4068 22024
rect 4120 22012 4126 22024
rect 4433 22015 4491 22021
rect 4433 22012 4445 22015
rect 4120 21984 4445 22012
rect 4120 21972 4126 21984
rect 4433 21981 4445 21984
rect 4479 21981 4491 22015
rect 4433 21975 4491 21981
rect 1949 21947 2007 21953
rect 1949 21913 1961 21947
rect 1995 21944 2007 21947
rect 3418 21944 3424 21956
rect 1995 21916 3424 21944
rect 1995 21913 2007 21916
rect 1949 21907 2007 21913
rect 3418 21904 3424 21916
rect 3476 21904 3482 21956
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2280 21848 3065 21876
rect 2280 21836 2286 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 4540 21876 4568 22052
rect 4893 22049 4905 22083
rect 4939 22080 4951 22083
rect 4982 22080 4988 22092
rect 4939 22052 4988 22080
rect 4939 22049 4951 22052
rect 4893 22043 4951 22049
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 5258 22080 5264 22092
rect 5219 22052 5264 22080
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 7009 22083 7067 22089
rect 7009 22049 7021 22083
rect 7055 22080 7067 22083
rect 8018 22080 8024 22092
rect 7055 22052 8024 22080
rect 7055 22049 7067 22052
rect 7009 22043 7067 22049
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8205 22083 8263 22089
rect 8205 22049 8217 22083
rect 8251 22049 8263 22083
rect 8312 22080 8340 22120
rect 10781 22117 10793 22151
rect 10827 22148 10839 22151
rect 11238 22148 11244 22160
rect 10827 22120 11244 22148
rect 10827 22117 10839 22120
rect 10781 22111 10839 22117
rect 11238 22108 11244 22120
rect 11296 22108 11302 22160
rect 8389 22083 8447 22089
rect 8389 22080 8401 22083
rect 8312 22052 8401 22080
rect 8205 22043 8263 22049
rect 8389 22049 8401 22052
rect 8435 22049 8447 22083
rect 9674 22080 9680 22092
rect 8389 22043 8447 22049
rect 8680 22052 9680 22080
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5442 22012 5448 22024
rect 5132 21984 5448 22012
rect 5132 21972 5138 21984
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 7282 22012 7288 22024
rect 7243 21984 7288 22012
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 8220 22012 8248 22043
rect 8680 22012 8708 22052
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 10597 22083 10655 22089
rect 10597 22080 10609 22083
rect 10192 22052 10609 22080
rect 10192 22040 10198 22052
rect 10597 22049 10609 22052
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 10873 22083 10931 22089
rect 10873 22049 10885 22083
rect 10919 22080 10931 22083
rect 11146 22080 11152 22092
rect 10919 22052 11152 22080
rect 10919 22049 10931 22052
rect 10873 22043 10931 22049
rect 11146 22040 11152 22052
rect 11204 22040 11210 22092
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 12250 22080 12256 22092
rect 11379 22052 12256 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22080 12495 22083
rect 14366 22080 14372 22092
rect 12483 22052 14372 22080
rect 12483 22049 12495 22052
rect 12437 22043 12495 22049
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 17865 22083 17923 22089
rect 17865 22049 17877 22083
rect 17911 22080 17923 22083
rect 18230 22080 18236 22092
rect 17911 22052 18236 22080
rect 17911 22049 17923 22052
rect 17865 22043 17923 22049
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 18690 22080 18696 22092
rect 18651 22052 18696 22080
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19789 22083 19847 22089
rect 19789 22080 19801 22083
rect 19576 22052 19801 22080
rect 19576 22040 19582 22052
rect 19789 22049 19801 22052
rect 19835 22049 19847 22083
rect 19789 22043 19847 22049
rect 8220 21984 8708 22012
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 9858 22012 9864 22024
rect 8803 21984 9864 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 11422 21972 11428 22024
rect 11480 22012 11486 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11480 21984 12173 22012
rect 11480 21972 11486 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 16172 21984 16221 22012
rect 16172 21972 16178 21984
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16482 22012 16488 22024
rect 16443 21984 16488 22012
rect 16209 21975 16267 21981
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 19889 22015 19947 22021
rect 19889 22012 19901 22015
rect 16632 21984 19901 22012
rect 16632 21972 16638 21984
rect 19889 21981 19901 21984
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 4614 21904 4620 21956
rect 4672 21944 4678 21956
rect 5169 21947 5227 21953
rect 5169 21944 5181 21947
rect 4672 21916 5181 21944
rect 4672 21904 4678 21916
rect 5169 21913 5181 21916
rect 5215 21913 5227 21947
rect 5169 21907 5227 21913
rect 6822 21904 6828 21956
rect 6880 21944 6886 21956
rect 9766 21944 9772 21956
rect 6880 21916 9772 21944
rect 6880 21904 6886 21916
rect 9766 21904 9772 21916
rect 9824 21904 9830 21956
rect 4706 21876 4712 21888
rect 4540 21848 4712 21876
rect 3053 21839 3111 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 11330 21876 11336 21888
rect 7616 21848 11336 21876
rect 7616 21836 7622 21848
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 14182 21876 14188 21888
rect 12032 21848 14188 21876
rect 12032 21836 12038 21848
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15746 21876 15752 21888
rect 15344 21848 15752 21876
rect 15344 21836 15350 21848
rect 15746 21836 15752 21848
rect 15804 21876 15810 21888
rect 18877 21879 18935 21885
rect 18877 21876 18889 21879
rect 15804 21848 18889 21876
rect 15804 21836 15810 21848
rect 18877 21845 18889 21848
rect 18923 21845 18935 21879
rect 18877 21839 18935 21845
rect 1104 21786 24840 21808
rect 1104 21734 4947 21786
rect 4999 21734 5011 21786
rect 5063 21734 5075 21786
rect 5127 21734 5139 21786
rect 5191 21734 12878 21786
rect 12930 21734 12942 21786
rect 12994 21734 13006 21786
rect 13058 21734 13070 21786
rect 13122 21734 20808 21786
rect 20860 21734 20872 21786
rect 20924 21734 20936 21786
rect 20988 21734 21000 21786
rect 21052 21734 24840 21786
rect 1104 21712 24840 21734
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 8389 21675 8447 21681
rect 8389 21672 8401 21675
rect 4028 21644 8401 21672
rect 4028 21632 4034 21644
rect 8389 21641 8401 21644
rect 8435 21641 8447 21675
rect 8389 21635 8447 21641
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 11425 21675 11483 21681
rect 11425 21672 11437 21675
rect 11388 21644 11437 21672
rect 11388 21632 11394 21644
rect 11425 21641 11437 21644
rect 11471 21641 11483 21675
rect 11425 21635 11483 21641
rect 11606 21632 11612 21684
rect 11664 21672 11670 21684
rect 14182 21672 14188 21684
rect 11664 21644 14044 21672
rect 14143 21644 14188 21672
rect 11664 21632 11670 21644
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 8110 21604 8116 21616
rect 7616 21576 8116 21604
rect 7616 21564 7622 21576
rect 8110 21564 8116 21576
rect 8168 21564 8174 21616
rect 8478 21564 8484 21616
rect 8536 21604 8542 21616
rect 9214 21604 9220 21616
rect 8536 21576 9220 21604
rect 8536 21564 8542 21576
rect 9214 21564 9220 21576
rect 9272 21604 9278 21616
rect 11146 21604 11152 21616
rect 9272 21576 11152 21604
rect 9272 21564 9278 21576
rect 11146 21564 11152 21576
rect 11204 21564 11210 21616
rect 11882 21564 11888 21616
rect 11940 21604 11946 21616
rect 12437 21607 12495 21613
rect 12437 21604 12449 21607
rect 11940 21576 12449 21604
rect 11940 21564 11946 21576
rect 12437 21573 12449 21576
rect 12483 21573 12495 21607
rect 12437 21567 12495 21573
rect 5353 21539 5411 21545
rect 2056 21508 3372 21536
rect 2056 21477 2084 21508
rect 3344 21480 3372 21508
rect 5353 21505 5365 21539
rect 5399 21536 5411 21539
rect 5810 21536 5816 21548
rect 5399 21508 5816 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 7800 21508 7880 21536
rect 7800 21496 7806 21508
rect 2041 21471 2099 21477
rect 2041 21437 2053 21471
rect 2087 21437 2099 21471
rect 3142 21468 3148 21480
rect 3103 21440 3148 21468
rect 2041 21431 2099 21437
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 3326 21468 3332 21480
rect 3287 21440 3332 21468
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3878 21428 3884 21480
rect 3936 21468 3942 21480
rect 4062 21468 4068 21480
rect 3936 21440 3981 21468
rect 4023 21440 4068 21468
rect 3936 21428 3942 21440
rect 4062 21428 4068 21440
rect 4120 21428 4126 21480
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 6546 21468 6552 21480
rect 5491 21440 6552 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 6546 21428 6552 21440
rect 6604 21428 6610 21480
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21468 6883 21471
rect 6914 21468 6920 21480
rect 6871 21440 6920 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 7852 21468 7880 21508
rect 8220 21508 9965 21536
rect 8220 21477 8248 21508
rect 9953 21505 9965 21508
rect 9999 21505 10011 21539
rect 13170 21536 13176 21548
rect 13131 21508 13176 21536
rect 9953 21499 10011 21505
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7852 21440 7941 21468
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 8205 21471 8263 21477
rect 8205 21437 8217 21471
rect 8251 21437 8263 21471
rect 8205 21431 8263 21437
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21437 9551 21471
rect 9493 21431 9551 21437
rect 3896 21400 3924 21428
rect 2240 21372 3924 21400
rect 2240 21341 2268 21372
rect 5718 21360 5724 21412
rect 5776 21400 5782 21412
rect 5905 21403 5963 21409
rect 5905 21400 5917 21403
rect 5776 21372 5917 21400
rect 5776 21360 5782 21372
rect 5905 21369 5917 21372
rect 5951 21369 5963 21403
rect 8110 21400 8116 21412
rect 5905 21363 5963 21369
rect 6932 21372 7972 21400
rect 8071 21372 8116 21400
rect 2225 21335 2283 21341
rect 2225 21301 2237 21335
rect 2271 21301 2283 21335
rect 4338 21332 4344 21344
rect 4299 21304 4344 21332
rect 2225 21295 2283 21301
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 4706 21292 4712 21344
rect 4764 21332 4770 21344
rect 6932 21332 6960 21372
rect 4764 21304 6960 21332
rect 7009 21335 7067 21341
rect 4764 21292 4770 21304
rect 7009 21301 7021 21335
rect 7055 21332 7067 21335
rect 7650 21332 7656 21344
rect 7055 21304 7656 21332
rect 7055 21301 7067 21304
rect 7009 21295 7067 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 7944 21332 7972 21372
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 9508 21400 9536 21431
rect 9582 21428 9588 21480
rect 9640 21468 9646 21480
rect 9766 21468 9772 21480
rect 9640 21440 9685 21468
rect 9727 21440 9772 21468
rect 9640 21428 9646 21440
rect 9766 21428 9772 21440
rect 9824 21468 9830 21480
rect 10962 21468 10968 21480
rect 9824 21440 10968 21468
rect 9824 21428 9830 21440
rect 10962 21428 10968 21440
rect 11020 21428 11026 21480
rect 11146 21428 11152 21480
rect 11204 21468 11210 21480
rect 11247 21471 11305 21477
rect 11247 21468 11259 21471
rect 11204 21440 11259 21468
rect 11204 21428 11210 21440
rect 11247 21437 11259 21440
rect 11293 21437 11305 21471
rect 12710 21468 12716 21480
rect 12671 21440 12716 21468
rect 11247 21431 11305 21437
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 14016 21477 14044 21644
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 16301 21675 16359 21681
rect 16301 21641 16313 21675
rect 16347 21672 16359 21675
rect 16482 21672 16488 21684
rect 16347 21644 16488 21672
rect 16347 21641 16359 21644
rect 16301 21635 16359 21641
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 15105 21539 15163 21545
rect 15105 21536 15117 21539
rect 14792 21508 15117 21536
rect 14792 21496 14798 21508
rect 15105 21505 15117 21508
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 17586 21496 17592 21548
rect 17644 21536 17650 21548
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 17644 21508 18613 21536
rect 17644 21496 17650 21508
rect 18601 21505 18613 21508
rect 18647 21505 18659 21539
rect 19242 21536 19248 21548
rect 18601 21499 18659 21505
rect 18708 21508 19248 21536
rect 14001 21471 14059 21477
rect 14001 21437 14013 21471
rect 14047 21437 14059 21471
rect 14001 21431 14059 21437
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21468 15347 21471
rect 15838 21468 15844 21480
rect 15335 21440 15844 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 16025 21471 16083 21477
rect 16025 21437 16037 21471
rect 16071 21468 16083 21471
rect 16298 21468 16304 21480
rect 16071 21440 16304 21468
rect 16071 21437 16083 21440
rect 16025 21431 16083 21437
rect 16298 21428 16304 21440
rect 16356 21428 16362 21480
rect 18708 21477 18736 21508
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 19058 21468 19064 21480
rect 19019 21440 19064 21468
rect 18693 21431 18751 21437
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 19150 21428 19156 21480
rect 19208 21468 19214 21480
rect 20073 21471 20131 21477
rect 19208 21440 19253 21468
rect 19208 21428 19214 21440
rect 20073 21437 20085 21471
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 10410 21400 10416 21412
rect 9508 21372 10416 21400
rect 10410 21360 10416 21372
rect 10468 21360 10474 21412
rect 12621 21403 12679 21409
rect 12621 21369 12633 21403
rect 12667 21400 12679 21403
rect 13170 21400 13176 21412
rect 12667 21372 13176 21400
rect 12667 21369 12679 21372
rect 12621 21363 12679 21369
rect 13170 21360 13176 21372
rect 13228 21360 13234 21412
rect 18046 21400 18052 21412
rect 18007 21372 18052 21400
rect 18046 21360 18052 21372
rect 18104 21360 18110 21412
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 20088 21400 20116 21431
rect 18380 21372 20116 21400
rect 18380 21360 18386 21372
rect 11146 21332 11152 21344
rect 7944 21304 11152 21332
rect 11146 21292 11152 21304
rect 11204 21332 11210 21344
rect 11974 21332 11980 21344
rect 11204 21304 11980 21332
rect 11204 21292 11210 21304
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 20162 21332 20168 21344
rect 20123 21304 20168 21332
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 1104 21242 24840 21264
rect 1104 21190 8912 21242
rect 8964 21190 8976 21242
rect 9028 21190 9040 21242
rect 9092 21190 9104 21242
rect 9156 21190 16843 21242
rect 16895 21190 16907 21242
rect 16959 21190 16971 21242
rect 17023 21190 17035 21242
rect 17087 21190 24840 21242
rect 1104 21168 24840 21190
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 20162 21128 20168 21140
rect 4120 21100 20168 21128
rect 4120 21088 4126 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 3050 21060 3056 21072
rect 2963 21032 3056 21060
rect 3050 21020 3056 21032
rect 3108 21060 3114 21072
rect 3694 21060 3700 21072
rect 3108 21032 3700 21060
rect 3108 21020 3114 21032
rect 3694 21020 3700 21032
rect 3752 21020 3758 21072
rect 6546 21060 6552 21072
rect 6507 21032 6552 21060
rect 6546 21020 6552 21032
rect 6604 21020 6610 21072
rect 8478 21060 8484 21072
rect 6932 21032 8484 21060
rect 1412 20964 2084 20992
rect 1412 20936 1440 20964
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 1670 20924 1676 20936
rect 1631 20896 1676 20924
rect 1670 20884 1676 20896
rect 1728 20884 1734 20936
rect 2056 20924 2084 20964
rect 2314 20952 2320 21004
rect 2372 20992 2378 21004
rect 4338 20992 4344 21004
rect 2372 20964 4200 20992
rect 4299 20964 4344 20992
rect 2372 20952 2378 20964
rect 2498 20924 2504 20936
rect 2056 20896 2504 20924
rect 2498 20884 2504 20896
rect 2556 20924 2562 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 2556 20896 4077 20924
rect 2556 20884 2562 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 4172 20924 4200 20964
rect 4338 20952 4344 20964
rect 4396 20952 4402 21004
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20992 5779 20995
rect 6932 20992 6960 21032
rect 8478 21020 8484 21032
rect 8536 21020 8542 21072
rect 9858 21060 9864 21072
rect 9819 21032 9864 21060
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 10410 21060 10416 21072
rect 10371 21032 10416 21060
rect 10410 21020 10416 21032
rect 10468 21020 10474 21072
rect 12710 21020 12716 21072
rect 12768 21060 12774 21072
rect 15841 21063 15899 21069
rect 15841 21060 15853 21063
rect 12768 21032 15853 21060
rect 12768 21020 12774 21032
rect 15841 21029 15853 21032
rect 15887 21029 15899 21063
rect 15841 21023 15899 21029
rect 7098 20992 7104 21004
rect 5767 20964 6960 20992
rect 7059 20964 7104 20992
rect 5767 20961 5779 20964
rect 5721 20955 5779 20961
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 7282 20992 7288 21004
rect 7243 20964 7288 20992
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20961 7435 20995
rect 7926 20992 7932 21004
rect 7887 20964 7932 20992
rect 7377 20955 7435 20961
rect 6822 20924 6828 20936
rect 4172 20896 6828 20924
rect 4065 20887 4123 20893
rect 6822 20884 6828 20896
rect 6880 20924 6886 20936
rect 7392 20924 7420 20955
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 9122 20952 9128 21004
rect 9180 20992 9186 21004
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9180 20964 9689 20992
rect 9180 20952 9186 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 9953 20995 10011 21001
rect 9953 20961 9965 20995
rect 9999 20992 10011 20995
rect 10594 20992 10600 21004
rect 9999 20964 10600 20992
rect 9999 20961 10011 20964
rect 9953 20955 10011 20961
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 12802 20992 12808 21004
rect 12483 20964 12808 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 7650 20924 7656 20936
rect 6880 20896 7420 20924
rect 7563 20896 7656 20924
rect 6880 20884 6886 20896
rect 7116 20868 7144 20896
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 11256 20924 11284 20955
rect 12802 20952 12808 20964
rect 12860 20992 12866 21004
rect 12989 20995 13047 21001
rect 12989 20992 13001 20995
rect 12860 20964 13001 20992
rect 12860 20952 12866 20964
rect 12989 20961 13001 20964
rect 13035 20961 13047 20995
rect 12989 20955 13047 20961
rect 13173 20995 13231 21001
rect 13173 20961 13185 20995
rect 13219 20992 13231 20995
rect 13354 20992 13360 21004
rect 13219 20964 13360 20992
rect 13219 20961 13231 20964
rect 13173 20955 13231 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15286 20992 15292 21004
rect 15247 20964 15292 20992
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20992 15531 20995
rect 15562 20992 15568 21004
rect 15519 20964 15568 20992
rect 15519 20961 15531 20964
rect 15473 20955 15531 20961
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20992 17095 20995
rect 18046 20992 18052 21004
rect 17083 20964 18052 20992
rect 17083 20961 17095 20964
rect 17037 20955 17095 20961
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 19058 20992 19064 21004
rect 18248 20964 19064 20992
rect 18248 20936 18276 20964
rect 19058 20952 19064 20964
rect 19116 20992 19122 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 19116 20964 19257 20992
rect 19116 20952 19122 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 7800 20896 11284 20924
rect 12345 20927 12403 20933
rect 7800 20884 7806 20896
rect 12345 20893 12357 20927
rect 12391 20893 12403 20927
rect 16114 20924 16120 20936
rect 12345 20887 12403 20893
rect 15580 20896 16120 20924
rect 7098 20816 7104 20868
rect 7156 20816 7162 20868
rect 7668 20856 7696 20884
rect 9122 20856 9128 20868
rect 7668 20828 9128 20856
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 11606 20856 11612 20868
rect 11164 20828 11612 20856
rect 6822 20748 6828 20800
rect 6880 20788 6886 20800
rect 11164 20788 11192 20828
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 12360 20856 12388 20887
rect 15580 20868 15608 20896
rect 16114 20884 16120 20896
rect 16172 20924 16178 20936
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16172 20896 16773 20924
rect 16172 20884 16178 20896
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 18230 20924 18236 20936
rect 18191 20896 18236 20924
rect 16761 20887 16819 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 12526 20856 12532 20868
rect 12360 20828 12532 20856
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 13357 20859 13415 20865
rect 13357 20856 13369 20859
rect 12676 20828 13369 20856
rect 12676 20816 12682 20828
rect 13357 20825 13369 20828
rect 13403 20825 13415 20859
rect 13357 20819 13415 20825
rect 15562 20816 15568 20868
rect 15620 20816 15626 20868
rect 11330 20788 11336 20800
rect 6880 20760 11192 20788
rect 11291 20760 11336 20788
rect 6880 20748 6886 20760
rect 11330 20748 11336 20760
rect 11388 20788 11394 20800
rect 11882 20788 11888 20800
rect 11388 20760 11888 20788
rect 11388 20748 11394 20760
rect 11882 20748 11888 20760
rect 11940 20748 11946 20800
rect 16298 20748 16304 20800
rect 16356 20788 16362 20800
rect 18230 20788 18236 20800
rect 16356 20760 18236 20788
rect 16356 20748 16362 20760
rect 18230 20748 18236 20760
rect 18288 20788 18294 20800
rect 19337 20791 19395 20797
rect 19337 20788 19349 20791
rect 18288 20760 19349 20788
rect 18288 20748 18294 20760
rect 19337 20757 19349 20760
rect 19383 20757 19395 20791
rect 19337 20751 19395 20757
rect 1104 20698 24840 20720
rect 1104 20646 4947 20698
rect 4999 20646 5011 20698
rect 5063 20646 5075 20698
rect 5127 20646 5139 20698
rect 5191 20646 12878 20698
rect 12930 20646 12942 20698
rect 12994 20646 13006 20698
rect 13058 20646 13070 20698
rect 13122 20646 20808 20698
rect 20860 20646 20872 20698
rect 20924 20646 20936 20698
rect 20988 20646 21000 20698
rect 21052 20646 24840 20698
rect 1104 20624 24840 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 7024 20556 9536 20584
rect 2038 20476 2044 20528
rect 2096 20516 2102 20528
rect 5353 20519 5411 20525
rect 5353 20516 5365 20519
rect 2096 20488 5365 20516
rect 2096 20476 2102 20488
rect 5353 20485 5365 20488
rect 5399 20485 5411 20519
rect 7024 20516 7052 20556
rect 5353 20479 5411 20485
rect 5460 20488 7052 20516
rect 3050 20448 3056 20460
rect 2608 20420 3056 20448
rect 2222 20380 2228 20392
rect 2183 20352 2228 20380
rect 2222 20340 2228 20352
rect 2280 20340 2286 20392
rect 2314 20340 2320 20392
rect 2372 20380 2378 20392
rect 2608 20389 2636 20420
rect 3050 20408 3056 20420
rect 3108 20408 3114 20460
rect 2593 20383 2651 20389
rect 2372 20352 2417 20380
rect 2372 20340 2378 20352
rect 2593 20349 2605 20383
rect 2639 20349 2651 20383
rect 2593 20343 2651 20349
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20349 2743 20383
rect 4706 20380 4712 20392
rect 4667 20352 4712 20380
rect 2685 20343 2743 20349
rect 2498 20272 2504 20324
rect 2556 20312 2562 20324
rect 2700 20312 2728 20343
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 4798 20340 4804 20392
rect 4856 20380 4862 20392
rect 5460 20389 5488 20488
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 7156 20488 7328 20516
rect 7156 20476 7162 20488
rect 7190 20448 7196 20460
rect 7024 20420 7196 20448
rect 7024 20389 7052 20420
rect 7190 20408 7196 20420
rect 7248 20408 7254 20460
rect 4893 20383 4951 20389
rect 4893 20380 4905 20383
rect 4856 20352 4905 20380
rect 4856 20340 4862 20352
rect 4893 20349 4905 20352
rect 4939 20349 4951 20383
rect 4893 20343 4951 20349
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20349 5503 20383
rect 5445 20343 5503 20349
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20380 7159 20383
rect 7300 20380 7328 20488
rect 8202 20476 8208 20528
rect 8260 20516 8266 20528
rect 8757 20519 8815 20525
rect 8757 20516 8769 20519
rect 8260 20488 8769 20516
rect 8260 20476 8266 20488
rect 8757 20485 8769 20488
rect 8803 20516 8815 20519
rect 8803 20488 9444 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 7147 20352 7328 20380
rect 8573 20383 8631 20389
rect 7147 20349 7159 20352
rect 7101 20343 7159 20349
rect 8573 20349 8585 20383
rect 8619 20380 8631 20383
rect 8846 20380 8852 20392
rect 8619 20352 8852 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 9416 20380 9444 20488
rect 9508 20448 9536 20556
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 10137 20587 10195 20593
rect 10137 20584 10149 20587
rect 9640 20556 10149 20584
rect 9640 20544 9646 20556
rect 10137 20553 10149 20556
rect 10183 20553 10195 20587
rect 10137 20547 10195 20553
rect 11425 20587 11483 20593
rect 11425 20553 11437 20587
rect 11471 20584 11483 20587
rect 15102 20584 15108 20596
rect 11471 20556 15108 20584
rect 11471 20553 11483 20556
rect 11425 20547 11483 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 18322 20584 18328 20596
rect 18283 20556 18328 20584
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 9677 20519 9735 20525
rect 9677 20485 9689 20519
rect 9723 20516 9735 20519
rect 11330 20516 11336 20528
rect 9723 20488 11336 20516
rect 9723 20485 9735 20488
rect 9677 20479 9735 20485
rect 11330 20476 11336 20488
rect 11388 20476 11394 20528
rect 11698 20448 11704 20460
rect 9508 20420 11704 20448
rect 11698 20408 11704 20420
rect 11756 20448 11762 20460
rect 11974 20448 11980 20460
rect 11756 20420 11980 20448
rect 11756 20408 11762 20420
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 15654 20448 15660 20460
rect 13412 20420 14504 20448
rect 15615 20420 15660 20448
rect 13412 20408 13418 20420
rect 9582 20380 9588 20392
rect 9416 20352 9588 20380
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 9950 20380 9956 20392
rect 9911 20352 9956 20380
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 11241 20383 11299 20389
rect 11241 20380 11253 20383
rect 11204 20352 11253 20380
rect 11204 20340 11210 20352
rect 11241 20349 11253 20352
rect 11287 20380 11299 20383
rect 11330 20380 11336 20392
rect 11287 20352 11336 20380
rect 11287 20349 11299 20352
rect 11241 20343 11299 20349
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20349 13231 20383
rect 13173 20343 13231 20349
rect 13449 20383 13507 20389
rect 13449 20349 13461 20383
rect 13495 20380 13507 20383
rect 14366 20380 14372 20392
rect 13495 20352 14372 20380
rect 13495 20349 13507 20352
rect 13449 20343 13507 20349
rect 2556 20284 2728 20312
rect 6825 20315 6883 20321
rect 2556 20272 2562 20284
rect 6825 20281 6837 20315
rect 6871 20312 6883 20315
rect 6914 20312 6920 20324
rect 6871 20284 6920 20312
rect 6871 20281 6883 20284
rect 6825 20275 6883 20281
rect 6914 20272 6920 20284
rect 6972 20272 6978 20324
rect 7193 20315 7251 20321
rect 7193 20312 7205 20315
rect 7024 20284 7205 20312
rect 7024 20256 7052 20284
rect 7193 20281 7205 20284
rect 7239 20281 7251 20315
rect 7558 20312 7564 20324
rect 7519 20284 7564 20312
rect 7193 20275 7251 20281
rect 7558 20272 7564 20284
rect 7616 20272 7622 20324
rect 9861 20315 9919 20321
rect 9861 20281 9873 20315
rect 9907 20312 9919 20315
rect 10962 20312 10968 20324
rect 9907 20284 10968 20312
rect 9907 20281 9919 20284
rect 9861 20275 9919 20281
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 7006 20204 7012 20256
rect 7064 20204 7070 20256
rect 13188 20244 13216 20343
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 14476 20380 14504 20420
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16574 20448 16580 20460
rect 16080 20420 16344 20448
rect 16535 20420 16580 20448
rect 16080 20408 16086 20420
rect 16316 20389 16344 20420
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 17126 20448 17132 20460
rect 16684 20420 17132 20448
rect 16684 20389 16712 20420
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17770 20408 17776 20460
rect 17828 20448 17834 20460
rect 18196 20451 18254 20457
rect 18196 20448 18208 20451
rect 17828 20420 18208 20448
rect 17828 20408 17834 20420
rect 18196 20417 18208 20420
rect 18242 20417 18254 20451
rect 18414 20448 18420 20460
rect 18375 20420 18420 20448
rect 18196 20411 18254 20417
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 14476 20352 16129 20380
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20349 16359 20383
rect 16301 20343 16359 20349
rect 16669 20383 16727 20389
rect 16669 20349 16681 20383
rect 16715 20349 16727 20383
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 16669 20343 16727 20349
rect 16776 20352 19625 20380
rect 14829 20315 14887 20321
rect 14829 20281 14841 20315
rect 14875 20312 14887 20315
rect 15286 20312 15292 20324
rect 14875 20284 15292 20312
rect 14875 20281 14887 20284
rect 14829 20275 14887 20281
rect 15286 20272 15292 20284
rect 15344 20312 15350 20324
rect 16776 20312 16804 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 15344 20284 16804 20312
rect 15344 20272 15350 20284
rect 17218 20272 17224 20324
rect 17276 20312 17282 20324
rect 18049 20315 18107 20321
rect 18049 20312 18061 20315
rect 17276 20284 18061 20312
rect 17276 20272 17282 20284
rect 18049 20281 18061 20284
rect 18095 20281 18107 20315
rect 19705 20315 19763 20321
rect 19705 20312 19717 20315
rect 18049 20275 18107 20281
rect 18156 20284 19717 20312
rect 15562 20244 15568 20256
rect 13188 20216 15568 20244
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 18156 20244 18184 20284
rect 19705 20281 19717 20284
rect 19751 20281 19763 20315
rect 19705 20275 19763 20281
rect 18690 20244 18696 20256
rect 16172 20216 18184 20244
rect 18651 20216 18696 20244
rect 16172 20204 16178 20216
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 1104 20154 24840 20176
rect 1104 20102 8912 20154
rect 8964 20102 8976 20154
rect 9028 20102 9040 20154
rect 9092 20102 9104 20154
rect 9156 20102 16843 20154
rect 16895 20102 16907 20154
rect 16959 20102 16971 20154
rect 17023 20102 17035 20154
rect 17087 20102 24840 20154
rect 1104 20080 24840 20102
rect 1489 20043 1547 20049
rect 1489 20009 1501 20043
rect 1535 20040 1547 20043
rect 3602 20040 3608 20052
rect 1535 20012 3608 20040
rect 1535 20009 1547 20012
rect 1489 20003 1547 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 4356 20012 6837 20040
rect 2130 19932 2136 19984
rect 2188 19972 2194 19984
rect 2590 19972 2596 19984
rect 2188 19944 2596 19972
rect 2188 19932 2194 19944
rect 2590 19932 2596 19944
rect 2648 19932 2654 19984
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1486 19904 1492 19916
rect 1443 19876 1492 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 4356 19913 4384 20012
rect 6825 20009 6837 20012
rect 6871 20040 6883 20043
rect 6914 20040 6920 20052
rect 6871 20012 6920 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 6914 20000 6920 20012
rect 6972 20040 6978 20052
rect 7742 20040 7748 20052
rect 6972 20012 7748 20040
rect 6972 20000 6978 20012
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 8110 20000 8116 20052
rect 8168 20040 8174 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8168 20012 8493 20040
rect 8168 20000 8174 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 8588 20012 13124 20040
rect 8386 19932 8392 19984
rect 8444 19972 8450 19984
rect 8588 19972 8616 20012
rect 8444 19944 8616 19972
rect 8444 19932 8450 19944
rect 9582 19932 9588 19984
rect 9640 19972 9646 19984
rect 13096 19972 13124 20012
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13228 20012 14105 20040
rect 13228 20000 13234 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 14700 20012 15485 20040
rect 14700 20000 14706 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 13538 19972 13544 19984
rect 9640 19944 9904 19972
rect 13096 19944 13544 19972
rect 9640 19932 9646 19944
rect 2409 19907 2467 19913
rect 2409 19904 2421 19907
rect 2096 19876 2421 19904
rect 2096 19864 2102 19876
rect 2409 19873 2421 19876
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 4341 19907 4399 19913
rect 4341 19873 4353 19907
rect 4387 19873 4399 19907
rect 5718 19904 5724 19916
rect 5679 19876 5724 19904
rect 4341 19867 4399 19873
rect 5718 19864 5724 19876
rect 5776 19864 5782 19916
rect 8018 19904 8024 19916
rect 7979 19876 8024 19904
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8297 19907 8355 19913
rect 8297 19904 8309 19907
rect 8260 19876 8309 19904
rect 8260 19864 8266 19876
rect 8297 19873 8309 19876
rect 8343 19873 8355 19907
rect 8297 19867 8355 19873
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 9766 19904 9772 19916
rect 9723 19876 9772 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 9876 19913 9904 19944
rect 13538 19932 13544 19944
rect 13596 19932 13602 19984
rect 13630 19932 13636 19984
rect 13688 19972 13694 19984
rect 18877 19975 18935 19981
rect 18877 19972 18889 19975
rect 13688 19944 14044 19972
rect 13688 19932 13694 19944
rect 9861 19907 9919 19913
rect 9861 19873 9873 19907
rect 9907 19904 9919 19907
rect 11054 19904 11060 19916
rect 9907 19876 11060 19904
rect 9907 19873 9919 19876
rect 9861 19867 9919 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 11422 19904 11428 19916
rect 11379 19876 11428 19904
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 12618 19904 12624 19916
rect 11655 19876 12624 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 14016 19913 14044 19944
rect 17420 19944 18889 19972
rect 17420 19913 17448 19944
rect 18877 19941 18889 19944
rect 18923 19941 18935 19975
rect 18877 19935 18935 19941
rect 13817 19907 13875 19913
rect 13817 19904 13829 19907
rect 12728 19876 13829 19904
rect 2556 19839 2614 19845
rect 2556 19805 2568 19839
rect 2602 19836 2614 19839
rect 2682 19836 2688 19848
rect 2602 19808 2688 19836
rect 2602 19805 2614 19808
rect 2556 19799 2614 19805
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 3050 19836 3056 19848
rect 2823 19808 3056 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 5902 19836 5908 19848
rect 5491 19808 5908 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 2130 19728 2136 19780
rect 2188 19768 2194 19780
rect 2869 19771 2927 19777
rect 2869 19768 2881 19771
rect 2188 19740 2881 19768
rect 2188 19728 2194 19740
rect 2869 19737 2881 19740
rect 2915 19737 2927 19771
rect 8110 19768 8116 19780
rect 8071 19740 8116 19768
rect 2869 19731 2927 19737
rect 8110 19728 8116 19740
rect 8168 19728 8174 19780
rect 9582 19728 9588 19780
rect 9640 19768 9646 19780
rect 9858 19768 9864 19780
rect 9640 19740 9864 19768
rect 9640 19728 9646 19740
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 2590 19660 2596 19712
rect 2648 19700 2654 19712
rect 2685 19703 2743 19709
rect 2685 19700 2697 19703
rect 2648 19672 2697 19700
rect 2648 19660 2654 19672
rect 2685 19669 2697 19672
rect 2731 19669 2743 19703
rect 2685 19663 2743 19669
rect 2774 19660 2780 19712
rect 2832 19700 2838 19712
rect 2958 19700 2964 19712
rect 2832 19672 2964 19700
rect 2832 19660 2838 19672
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 7742 19700 7748 19712
rect 4571 19672 7748 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 9953 19703 10011 19709
rect 9953 19700 9965 19703
rect 8352 19672 9965 19700
rect 8352 19660 8358 19672
rect 9953 19669 9965 19672
rect 9999 19669 10011 19703
rect 9953 19663 10011 19669
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 12728 19709 12756 19876
rect 13817 19873 13829 19876
rect 13863 19873 13875 19907
rect 13817 19867 13875 19873
rect 14001 19907 14059 19913
rect 14001 19873 14013 19907
rect 14047 19873 14059 19907
rect 14001 19867 14059 19873
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19904 17555 19907
rect 17586 19904 17592 19916
rect 17543 19876 17592 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 10468 19672 12725 19700
rect 10468 19660 10474 19672
rect 12713 19669 12725 19672
rect 12759 19669 12771 19703
rect 12713 19663 12771 19669
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 14642 19700 14648 19712
rect 13596 19672 14648 19700
rect 13596 19660 13602 19672
rect 14642 19660 14648 19672
rect 14700 19700 14706 19712
rect 15304 19700 15332 19867
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 17770 19904 17776 19916
rect 17731 19876 17776 19904
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 17954 19904 17960 19916
rect 17915 19876 17960 19904
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 18785 19907 18843 19913
rect 18785 19904 18797 19907
rect 18656 19876 18797 19904
rect 18656 19864 18662 19876
rect 18785 19873 18797 19876
rect 18831 19904 18843 19907
rect 19150 19904 19156 19916
rect 18831 19876 19156 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 14700 19672 15332 19700
rect 14700 19660 14706 19672
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 16853 19703 16911 19709
rect 16853 19700 16865 19703
rect 16724 19672 16865 19700
rect 16724 19660 16730 19672
rect 16853 19669 16865 19672
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 1104 19610 24840 19632
rect 1104 19558 4947 19610
rect 4999 19558 5011 19610
rect 5063 19558 5075 19610
rect 5127 19558 5139 19610
rect 5191 19558 12878 19610
rect 12930 19558 12942 19610
rect 12994 19558 13006 19610
rect 13058 19558 13070 19610
rect 13122 19558 20808 19610
rect 20860 19558 20872 19610
rect 20924 19558 20936 19610
rect 20988 19558 21000 19610
rect 21052 19558 24840 19610
rect 1104 19536 24840 19558
rect 2590 19456 2596 19508
rect 2648 19496 2654 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2648 19468 2973 19496
rect 2648 19456 2654 19468
rect 2961 19465 2973 19468
rect 3007 19465 3019 19499
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 2961 19459 3019 19465
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 5902 19456 5908 19508
rect 5960 19496 5966 19508
rect 6457 19499 6515 19505
rect 6457 19496 6469 19499
rect 5960 19468 6469 19496
rect 5960 19456 5966 19468
rect 6457 19465 6469 19468
rect 6503 19465 6515 19499
rect 6457 19459 6515 19465
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 7929 19499 7987 19505
rect 7929 19496 7941 19499
rect 7800 19468 7941 19496
rect 7800 19456 7806 19468
rect 7929 19465 7941 19468
rect 7975 19465 7987 19499
rect 7929 19459 7987 19465
rect 2682 19388 2688 19440
rect 2740 19428 2746 19440
rect 2823 19431 2881 19437
rect 2823 19428 2835 19431
rect 2740 19400 2835 19428
rect 2740 19388 2746 19400
rect 2823 19397 2835 19400
rect 2869 19397 2881 19431
rect 2823 19391 2881 19397
rect 4525 19431 4583 19437
rect 4525 19397 4537 19431
rect 4571 19428 4583 19431
rect 5442 19428 5448 19440
rect 4571 19400 5448 19428
rect 4571 19397 4583 19400
rect 4525 19391 4583 19397
rect 3050 19360 3056 19372
rect 3011 19332 3056 19360
rect 3050 19320 3056 19332
rect 3108 19320 3114 19372
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 4617 19363 4675 19369
rect 4617 19360 4629 19363
rect 3660 19332 4629 19360
rect 3660 19320 3666 19332
rect 4617 19329 4629 19332
rect 4663 19329 4675 19363
rect 4617 19323 4675 19329
rect 4724 19304 4752 19400
rect 5442 19388 5448 19400
rect 5500 19388 5506 19440
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 6546 19428 6552 19440
rect 6236 19400 6552 19428
rect 6236 19388 6242 19400
rect 6546 19388 6552 19400
rect 6604 19388 6610 19440
rect 7944 19428 7972 19459
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 8168 19468 8401 19496
rect 8168 19456 8174 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 8389 19459 8447 19465
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 13354 19496 13360 19508
rect 9631 19468 13360 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 14366 19496 14372 19508
rect 14327 19468 14372 19496
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18288 19468 18337 19496
rect 18288 19456 18294 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18325 19459 18383 19465
rect 10505 19431 10563 19437
rect 10505 19428 10517 19431
rect 7944 19400 10517 19428
rect 10505 19397 10517 19400
rect 10551 19428 10563 19431
rect 10870 19428 10876 19440
rect 10551 19400 10876 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 10962 19388 10968 19440
rect 11020 19388 11026 19440
rect 10980 19360 11008 19388
rect 16114 19360 16120 19372
rect 10980 19332 11100 19360
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19261 1731 19295
rect 1673 19255 1731 19261
rect 1688 19224 1716 19255
rect 1762 19252 1768 19304
rect 1820 19292 1826 19304
rect 2685 19295 2743 19301
rect 1820 19264 1865 19292
rect 1820 19252 1826 19264
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 2958 19292 2964 19304
rect 2731 19264 2964 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 4338 19252 4344 19304
rect 4396 19301 4402 19304
rect 4396 19295 4454 19301
rect 4396 19261 4408 19295
rect 4442 19292 4454 19295
rect 4442 19264 4660 19292
rect 4442 19261 4454 19264
rect 4396 19255 4454 19261
rect 4396 19252 4402 19255
rect 4632 19236 4660 19264
rect 4706 19252 4712 19304
rect 4764 19252 4770 19304
rect 6178 19252 6184 19304
rect 6236 19292 6242 19304
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 6236 19264 6653 19292
rect 6236 19252 6242 19264
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7006 19292 7012 19304
rect 6871 19264 7012 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19292 8263 19295
rect 8294 19292 8300 19304
rect 8251 19264 8300 19292
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 9485 19295 9543 19301
rect 9485 19261 9497 19295
rect 9531 19292 9543 19295
rect 10410 19292 10416 19304
rect 9531 19264 10416 19292
rect 9531 19261 9543 19264
rect 9485 19255 9543 19261
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 10962 19292 10968 19304
rect 10827 19264 10968 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 2406 19224 2412 19236
rect 1688 19196 2412 19224
rect 2406 19184 2412 19196
rect 2464 19184 2470 19236
rect 3418 19224 3424 19236
rect 3379 19196 3424 19224
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 4249 19227 4307 19233
rect 4249 19193 4261 19227
rect 4295 19193 4307 19227
rect 4249 19187 4307 19193
rect 4264 19156 4292 19187
rect 4614 19184 4620 19236
rect 4672 19184 4678 19236
rect 7742 19184 7748 19236
rect 7800 19224 7806 19236
rect 8113 19227 8171 19233
rect 8113 19224 8125 19227
rect 7800 19196 8125 19224
rect 7800 19184 7806 19196
rect 8113 19193 8125 19196
rect 8159 19193 8171 19227
rect 10686 19224 10692 19236
rect 10647 19196 10692 19224
rect 8113 19187 8171 19193
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 11072 19224 11100 19332
rect 15304 19332 16120 19360
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 10928 19196 11100 19224
rect 10928 19184 10934 19196
rect 11146 19184 11152 19236
rect 11204 19224 11210 19236
rect 11241 19227 11299 19233
rect 11241 19224 11253 19227
rect 11204 19196 11253 19224
rect 11204 19184 11210 19196
rect 11241 19193 11253 19196
rect 11287 19193 11299 19227
rect 11241 19187 11299 19193
rect 13170 19184 13176 19236
rect 13228 19224 13234 19236
rect 13464 19224 13492 19255
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 13909 19295 13967 19301
rect 13909 19292 13921 19295
rect 13780 19264 13921 19292
rect 13780 19252 13786 19264
rect 13909 19261 13921 19264
rect 13955 19261 13967 19295
rect 13909 19255 13967 19261
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 15304 19292 15332 19332
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 17126 19360 17132 19372
rect 16408 19332 17132 19360
rect 14139 19264 15332 19292
rect 15381 19295 15439 19301
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 15470 19292 15476 19304
rect 15427 19264 15476 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 16022 19292 16028 19304
rect 15983 19264 16028 19292
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16408 19301 16436 19332
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 18230 19369 18236 19372
rect 18196 19363 18236 19369
rect 18196 19360 18208 19363
rect 17788 19332 18208 19360
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19261 16451 19295
rect 16393 19255 16451 19261
rect 13228 19196 13492 19224
rect 13228 19184 13234 19196
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 16408 19224 16436 19255
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 17788 19292 17816 19332
rect 18196 19329 18208 19332
rect 18288 19360 18294 19372
rect 18417 19363 18475 19369
rect 18288 19332 18344 19360
rect 18196 19323 18236 19329
rect 18230 19320 18236 19323
rect 18288 19320 18294 19332
rect 18417 19329 18429 19363
rect 18463 19360 18475 19363
rect 18463 19332 18497 19360
rect 18463 19329 18475 19332
rect 18417 19323 18475 19329
rect 16540 19264 17816 19292
rect 16540 19252 16546 19264
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18432 19292 18460 19323
rect 17920 19264 18460 19292
rect 17920 19252 17926 19264
rect 14240 19196 16436 19224
rect 14240 19184 14246 19196
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 17126 19224 17132 19236
rect 16632 19196 17132 19224
rect 16632 19184 16638 19196
rect 17126 19184 17132 19196
rect 17184 19224 17190 19236
rect 18049 19227 18107 19233
rect 18049 19224 18061 19227
rect 17184 19196 18061 19224
rect 17184 19184 17190 19196
rect 18049 19193 18061 19196
rect 18095 19193 18107 19227
rect 18049 19187 18107 19193
rect 4338 19156 4344 19168
rect 4264 19128 4344 19156
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 7009 19159 7067 19165
rect 7009 19125 7021 19159
rect 7055 19156 7067 19159
rect 7374 19156 7380 19168
rect 7055 19128 7380 19156
rect 7055 19125 7067 19128
rect 7009 19119 7067 19125
rect 7374 19116 7380 19128
rect 7432 19156 7438 19168
rect 8202 19156 8208 19168
rect 7432 19128 8208 19156
rect 7432 19116 7438 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10042 19156 10048 19168
rect 9732 19128 10048 19156
rect 9732 19116 9738 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 16298 19156 16304 19168
rect 15804 19128 16304 19156
rect 15804 19116 15810 19128
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 18693 19159 18751 19165
rect 18693 19156 18705 19159
rect 18380 19128 18705 19156
rect 18380 19116 18386 19128
rect 18693 19125 18705 19128
rect 18739 19125 18751 19159
rect 18693 19119 18751 19125
rect 1104 19066 24840 19088
rect 1104 19014 8912 19066
rect 8964 19014 8976 19066
rect 9028 19014 9040 19066
rect 9092 19014 9104 19066
rect 9156 19014 16843 19066
rect 16895 19014 16907 19066
rect 16959 19014 16971 19066
rect 17023 19014 17035 19066
rect 17087 19014 24840 19066
rect 1104 18992 24840 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 2406 18952 2412 18964
rect 1544 18924 2412 18952
rect 1544 18912 1550 18924
rect 2406 18912 2412 18924
rect 2464 18952 2470 18964
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 2464 18924 2789 18952
rect 2464 18912 2470 18924
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 6512 18924 7420 18952
rect 6512 18912 6518 18924
rect 4522 18884 4528 18896
rect 4264 18856 4528 18884
rect 4264 18825 4292 18856
rect 4522 18844 4528 18856
rect 4580 18884 4586 18896
rect 4580 18856 4844 18884
rect 4580 18844 4586 18856
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 4614 18776 4620 18828
rect 4672 18816 4678 18828
rect 4816 18825 4844 18856
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4672 18788 4721 18816
rect 4672 18776 4678 18788
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 4801 18819 4859 18825
rect 4801 18785 4813 18819
rect 4847 18785 4859 18819
rect 4801 18779 4859 18785
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 7282 18816 7288 18828
rect 6963 18788 7144 18816
rect 7243 18788 7288 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4154 18748 4160 18760
rect 3936 18720 4160 18748
rect 3936 18708 3942 18720
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 5684 18720 6285 18748
rect 5684 18708 5690 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 3568 18584 5273 18612
rect 3568 18572 3574 18584
rect 5261 18581 5273 18584
rect 5307 18581 5319 18615
rect 7024 18612 7052 18711
rect 7116 18680 7144 18788
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 7392 18816 7420 18924
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7708 18924 8493 18952
rect 7708 18912 7714 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 10134 18952 10140 18964
rect 9999 18924 10140 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 8496 18884 8524 18915
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 11977 18955 12035 18961
rect 11977 18952 11989 18955
rect 10928 18924 11989 18952
rect 10928 18912 10934 18924
rect 11977 18921 11989 18924
rect 12023 18921 12035 18955
rect 11977 18915 12035 18921
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 15473 18955 15531 18961
rect 15473 18952 15485 18955
rect 13780 18924 15485 18952
rect 13780 18912 13786 18924
rect 15473 18921 15485 18924
rect 15519 18921 15531 18955
rect 15473 18915 15531 18921
rect 18230 18912 18236 18964
rect 18288 18952 18294 18964
rect 19153 18955 19211 18961
rect 19153 18952 19165 18955
rect 18288 18924 19165 18952
rect 18288 18912 18294 18924
rect 19153 18921 19165 18924
rect 19199 18921 19211 18955
rect 19153 18915 19211 18921
rect 10410 18884 10416 18896
rect 8496 18856 10416 18884
rect 10410 18844 10416 18856
rect 10468 18884 10474 18896
rect 16022 18884 16028 18896
rect 10468 18856 10732 18884
rect 10468 18844 10474 18856
rect 10704 18825 10732 18856
rect 13832 18856 16028 18884
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 7392 18788 8309 18816
rect 8297 18785 8309 18788
rect 8343 18785 8355 18819
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 8297 18779 8355 18785
rect 9508 18788 10333 18816
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7374 18748 7380 18760
rect 7239 18720 7380 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 9508 18748 9536 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11701 18819 11759 18825
rect 10836 18788 10881 18816
rect 10836 18776 10842 18788
rect 11701 18785 11713 18819
rect 11747 18816 11759 18819
rect 11790 18816 11796 18828
rect 11747 18788 11796 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18816 11943 18819
rect 12618 18816 12624 18828
rect 11931 18788 12624 18816
rect 11931 18785 11943 18788
rect 11885 18779 11943 18785
rect 12618 18776 12624 18788
rect 12676 18816 12682 18828
rect 13630 18816 13636 18828
rect 12676 18788 13636 18816
rect 12676 18776 12682 18788
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 13832 18825 13860 18856
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18785 13875 18819
rect 14182 18816 14188 18828
rect 14143 18788 14188 18816
rect 13817 18779 13875 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18816 14427 18819
rect 15194 18816 15200 18828
rect 14415 18788 15200 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15344 18788 15389 18816
rect 15344 18776 15350 18788
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 16853 18819 16911 18825
rect 16853 18816 16865 18819
rect 16724 18788 16865 18816
rect 16724 18776 16730 18788
rect 16853 18785 16865 18788
rect 16899 18785 16911 18819
rect 16853 18779 16911 18785
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 17920 18788 19073 18816
rect 17920 18776 17926 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 7524 18720 9536 18748
rect 7524 18708 7530 18720
rect 7650 18680 7656 18692
rect 7116 18652 7656 18680
rect 7650 18640 7656 18652
rect 7708 18640 7714 18692
rect 9508 18680 9536 18720
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9640 18720 10425 18748
rect 9640 18708 9646 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 13906 18748 13912 18760
rect 13867 18720 13912 18748
rect 10413 18711 10471 18717
rect 10042 18680 10048 18692
rect 9508 18652 10048 18680
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10428 18680 10456 18711
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 15528 18720 16589 18748
rect 15528 18708 15534 18720
rect 16577 18717 16589 18720
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 19518 18680 19524 18692
rect 10428 18652 15884 18680
rect 9674 18612 9680 18624
rect 7024 18584 9680 18612
rect 5261 18575 5319 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 13449 18615 13507 18621
rect 13449 18581 13461 18615
rect 13495 18612 13507 18615
rect 15746 18612 15752 18624
rect 13495 18584 15752 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 15856 18612 15884 18652
rect 17512 18652 19524 18680
rect 17512 18612 17540 18652
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 15856 18584 17540 18612
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 17957 18615 18015 18621
rect 17957 18612 17969 18615
rect 17920 18584 17969 18612
rect 17920 18572 17926 18584
rect 17957 18581 17969 18584
rect 18003 18581 18015 18615
rect 17957 18575 18015 18581
rect 1104 18522 24840 18544
rect 1104 18470 4947 18522
rect 4999 18470 5011 18522
rect 5063 18470 5075 18522
rect 5127 18470 5139 18522
rect 5191 18470 12878 18522
rect 12930 18470 12942 18522
rect 12994 18470 13006 18522
rect 13058 18470 13070 18522
rect 13122 18470 20808 18522
rect 20860 18470 20872 18522
rect 20924 18470 20936 18522
rect 20988 18470 21000 18522
rect 21052 18470 24840 18522
rect 1104 18448 24840 18470
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8570 18408 8576 18420
rect 8352 18380 8576 18408
rect 8352 18368 8358 18380
rect 8570 18368 8576 18380
rect 8628 18368 8634 18420
rect 9861 18411 9919 18417
rect 9861 18377 9873 18411
rect 9907 18408 9919 18411
rect 10134 18408 10140 18420
rect 9907 18380 10140 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 10134 18368 10140 18380
rect 10192 18408 10198 18420
rect 10192 18380 19472 18408
rect 10192 18368 10198 18380
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 11146 18340 11152 18352
rect 10919 18312 11152 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 13354 18340 13360 18352
rect 13004 18312 13360 18340
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 2498 18272 2504 18284
rect 2455 18244 2504 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 2498 18232 2504 18244
rect 2556 18272 2562 18284
rect 3510 18272 3516 18284
rect 2556 18244 3372 18272
rect 3471 18244 3516 18272
rect 2556 18232 2562 18244
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18204 2099 18207
rect 2682 18204 2688 18216
rect 2087 18176 2688 18204
rect 2087 18173 2099 18176
rect 2041 18167 2099 18173
rect 2682 18164 2688 18176
rect 2740 18204 2746 18216
rect 3050 18204 3056 18216
rect 2740 18176 3056 18204
rect 2740 18164 2746 18176
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3237 18207 3295 18213
rect 3237 18173 3249 18207
rect 3283 18173 3295 18207
rect 3344 18204 3372 18244
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4338 18272 4344 18284
rect 4212 18244 4344 18272
rect 4212 18232 4218 18244
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 6822 18232 6828 18284
rect 6880 18232 6886 18284
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 11238 18272 11244 18284
rect 8260 18244 11100 18272
rect 11199 18244 11244 18272
rect 8260 18232 8266 18244
rect 5721 18207 5779 18213
rect 5721 18204 5733 18207
rect 3344 18176 5733 18204
rect 3237 18167 3295 18173
rect 5721 18173 5733 18176
rect 5767 18173 5779 18207
rect 6840 18204 6868 18232
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 6840 18176 7021 18204
rect 5721 18167 5779 18173
rect 7009 18173 7021 18176
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 7377 18207 7435 18213
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 7466 18204 7472 18216
rect 7423 18176 7472 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 1762 18096 1768 18148
rect 1820 18136 1826 18148
rect 1857 18139 1915 18145
rect 1857 18136 1869 18139
rect 1820 18108 1869 18136
rect 1820 18096 1826 18108
rect 1857 18105 1869 18108
rect 1903 18105 1915 18139
rect 3252 18136 3280 18167
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18173 8355 18207
rect 8570 18204 8576 18216
rect 8531 18176 8576 18204
rect 8297 18167 8355 18173
rect 1857 18099 1915 18105
rect 2056 18108 3280 18136
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 2056 18068 2084 18108
rect 1452 18040 2084 18068
rect 3252 18068 3280 18108
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 6362 18136 6368 18148
rect 4948 18108 6368 18136
rect 4948 18096 4954 18108
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 6825 18139 6883 18145
rect 6825 18105 6837 18139
rect 6871 18136 6883 18139
rect 7558 18136 7564 18148
rect 6871 18108 7564 18136
rect 6871 18105 6883 18108
rect 6825 18099 6883 18105
rect 7558 18096 7564 18108
rect 7616 18096 7622 18148
rect 3602 18068 3608 18080
rect 3252 18040 3608 18068
rect 1452 18028 1458 18040
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4617 18071 4675 18077
rect 4617 18068 4629 18071
rect 4396 18040 4629 18068
rect 4396 18028 4402 18040
rect 4617 18037 4629 18040
rect 4663 18037 4675 18071
rect 4617 18031 4675 18037
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5813 18071 5871 18077
rect 5813 18068 5825 18071
rect 5592 18040 5825 18068
rect 5592 18028 5598 18040
rect 5813 18037 5825 18040
rect 5859 18037 5871 18071
rect 5813 18031 5871 18037
rect 5902 18028 5908 18080
rect 5960 18068 5966 18080
rect 8312 18068 8340 18167
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 10778 18204 10784 18216
rect 10739 18176 10784 18204
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 11072 18213 11100 18244
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 13004 18272 13032 18312
rect 13354 18300 13360 18312
rect 13412 18340 13418 18352
rect 13722 18340 13728 18352
rect 13412 18312 13728 18340
rect 13412 18300 13418 18312
rect 13722 18300 13728 18312
rect 13780 18300 13786 18352
rect 18598 18272 18604 18284
rect 12768 18244 13032 18272
rect 18559 18244 18604 18272
rect 12768 18232 12774 18244
rect 12820 18213 12848 18244
rect 11057 18207 11115 18213
rect 11057 18173 11069 18207
rect 11103 18173 11115 18207
rect 11057 18167 11115 18173
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18173 12863 18207
rect 12805 18167 12863 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18173 12955 18207
rect 13004 18204 13032 18244
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 13004 18176 13369 18204
rect 12897 18167 12955 18173
rect 13357 18173 13369 18176
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 13906 18204 13912 18216
rect 13587 18176 13912 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 12912 18136 12940 18167
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 15470 18204 15476 18216
rect 15431 18176 15476 18204
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15746 18204 15752 18216
rect 15707 18176 15752 18204
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 19444 18213 19472 18380
rect 19518 18368 19524 18420
rect 19576 18408 19582 18420
rect 19576 18380 19621 18408
rect 19576 18368 19582 18380
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 18012 18176 18061 18204
rect 18012 18164 18018 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18233 18207 18291 18213
rect 18233 18173 18245 18207
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 13630 18136 13636 18148
rect 12912 18108 13636 18136
rect 13630 18096 13636 18108
rect 13688 18096 13694 18148
rect 17129 18139 17187 18145
rect 17129 18105 17141 18139
rect 17175 18136 17187 18139
rect 17862 18136 17868 18148
rect 17175 18108 17868 18136
rect 17175 18105 17187 18108
rect 17129 18099 17187 18105
rect 17862 18096 17868 18108
rect 17920 18136 17926 18148
rect 18248 18136 18276 18167
rect 17920 18108 18276 18136
rect 17920 18096 17926 18108
rect 13814 18068 13820 18080
rect 5960 18040 8340 18068
rect 13775 18040 13820 18068
rect 5960 18028 5966 18040
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 16390 18068 16396 18080
rect 15344 18040 16396 18068
rect 15344 18028 15350 18040
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 1104 17978 24840 18000
rect 1104 17926 8912 17978
rect 8964 17926 8976 17978
rect 9028 17926 9040 17978
rect 9092 17926 9104 17978
rect 9156 17926 16843 17978
rect 16895 17926 16907 17978
rect 16959 17926 16971 17978
rect 17023 17926 17035 17978
rect 17087 17926 24840 17978
rect 1104 17904 24840 17926
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 4614 17864 4620 17876
rect 4479 17836 4620 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 7006 17864 7012 17876
rect 6967 17836 7012 17864
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 14366 17864 14372 17876
rect 12492 17836 14372 17864
rect 12492 17824 12498 17836
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16485 17867 16543 17873
rect 16485 17864 16497 17867
rect 15804 17836 16497 17864
rect 15804 17824 15810 17836
rect 16485 17833 16497 17836
rect 16531 17833 16543 17867
rect 16485 17827 16543 17833
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 1670 17796 1676 17808
rect 1627 17768 1676 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 1670 17756 1676 17768
rect 1728 17756 1734 17808
rect 5534 17796 5540 17808
rect 2240 17768 5540 17796
rect 2240 17737 2268 17768
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 13906 17756 13912 17808
rect 13964 17796 13970 17808
rect 18693 17799 18751 17805
rect 18693 17796 18705 17799
rect 13964 17768 18705 17796
rect 13964 17756 13970 17768
rect 18693 17765 18705 17768
rect 18739 17765 18751 17799
rect 18693 17759 18751 17765
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17697 2283 17731
rect 2225 17691 2283 17697
rect 2314 17688 2320 17740
rect 2372 17728 2378 17740
rect 2372 17700 2417 17728
rect 2372 17688 2378 17700
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 2556 17700 2605 17728
rect 2556 17688 2562 17700
rect 2593 17697 2605 17700
rect 2639 17728 2651 17731
rect 2682 17728 2688 17740
rect 2639 17700 2688 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 2958 17728 2964 17740
rect 2823 17700 2964 17728
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 3881 17731 3939 17737
rect 3881 17697 3893 17731
rect 3927 17697 3939 17731
rect 4338 17728 4344 17740
rect 4299 17700 4344 17728
rect 3881 17691 3939 17697
rect 3896 17660 3924 17691
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 6178 17728 6184 17740
rect 4448 17700 6184 17728
rect 4448 17660 4476 17700
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 8113 17731 8171 17737
rect 8113 17728 8125 17731
rect 7432 17700 8125 17728
rect 7432 17688 7438 17700
rect 8113 17697 8125 17700
rect 8159 17697 8171 17731
rect 8113 17691 8171 17697
rect 8202 17688 8208 17740
rect 8260 17728 8266 17740
rect 10781 17731 10839 17737
rect 8260 17700 8305 17728
rect 8260 17688 8266 17700
rect 10781 17697 10793 17731
rect 10827 17697 10839 17731
rect 10781 17691 10839 17697
rect 10873 17731 10931 17737
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 12437 17731 12495 17737
rect 10919 17700 12296 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 3896 17632 4476 17660
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 5718 17660 5724 17672
rect 5679 17632 5724 17660
rect 5445 17623 5503 17629
rect 4614 17552 4620 17604
rect 4672 17592 4678 17604
rect 4890 17592 4896 17604
rect 4672 17564 4896 17592
rect 4672 17552 4678 17564
rect 4890 17552 4896 17564
rect 4948 17552 4954 17604
rect 3326 17484 3332 17536
rect 3384 17524 3390 17536
rect 3510 17524 3516 17536
rect 3384 17496 3516 17524
rect 3384 17484 3390 17496
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 3694 17524 3700 17536
rect 3655 17496 3700 17524
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 5460 17524 5488 17623
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 7926 17660 7932 17672
rect 7839 17632 7932 17660
rect 7926 17620 7932 17632
rect 7984 17660 7990 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 7984 17632 10609 17660
rect 7984 17620 7990 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10796 17660 10824 17691
rect 11606 17660 11612 17672
rect 10796 17632 11612 17660
rect 10597 17623 10655 17629
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 12158 17660 12164 17672
rect 12216 17669 12222 17672
rect 11716 17632 12164 17660
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 8662 17592 8668 17604
rect 7064 17564 8668 17592
rect 7064 17552 7070 17564
rect 8662 17552 8668 17564
rect 8720 17552 8726 17604
rect 11422 17552 11428 17604
rect 11480 17592 11486 17604
rect 11716 17592 11744 17632
rect 12158 17620 12164 17632
rect 12216 17623 12226 17669
rect 12268 17660 12296 17700
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 13814 17728 13820 17740
rect 12483 17700 13820 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 15838 17728 15844 17740
rect 15519 17700 15844 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 16022 17728 16028 17740
rect 15983 17700 16028 17728
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16209 17731 16267 17737
rect 16209 17697 16221 17731
rect 16255 17728 16267 17731
rect 16482 17728 16488 17740
rect 16255 17700 16488 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17497 17731 17555 17737
rect 17497 17728 17509 17731
rect 16632 17700 17509 17728
rect 16632 17688 16638 17700
rect 17497 17697 17509 17700
rect 17543 17697 17555 17731
rect 17497 17691 17555 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 13354 17660 13360 17672
rect 12268 17632 13360 17660
rect 12216 17620 12222 17623
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 13648 17632 15301 17660
rect 11480 17564 11744 17592
rect 11480 17552 11486 17564
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 13648 17592 13676 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 13228 17564 13676 17592
rect 13725 17595 13783 17601
rect 13228 17552 13234 17564
rect 13725 17561 13737 17595
rect 13771 17592 13783 17595
rect 18616 17592 18644 17691
rect 13771 17564 18644 17592
rect 13771 17561 13783 17564
rect 13725 17555 13783 17561
rect 5902 17524 5908 17536
rect 5460 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8389 17527 8447 17533
rect 8389 17524 8401 17527
rect 8076 17496 8401 17524
rect 8076 17484 8082 17496
rect 8389 17493 8401 17496
rect 8435 17493 8447 17527
rect 8389 17487 8447 17493
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10836 17496 11069 17524
rect 10836 17484 10842 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 13740 17524 13768 17555
rect 11756 17496 13768 17524
rect 11756 17484 11762 17496
rect 13814 17484 13820 17536
rect 13872 17524 13878 17536
rect 17681 17527 17739 17533
rect 17681 17524 17693 17527
rect 13872 17496 17693 17524
rect 13872 17484 13878 17496
rect 17681 17493 17693 17496
rect 17727 17493 17739 17527
rect 17681 17487 17739 17493
rect 1104 17434 24840 17456
rect 1104 17382 4947 17434
rect 4999 17382 5011 17434
rect 5063 17382 5075 17434
rect 5127 17382 5139 17434
rect 5191 17382 12878 17434
rect 12930 17382 12942 17434
rect 12994 17382 13006 17434
rect 13058 17382 13070 17434
rect 13122 17382 20808 17434
rect 20860 17382 20872 17434
rect 20924 17382 20936 17434
rect 20988 17382 21000 17434
rect 21052 17382 24840 17434
rect 1104 17360 24840 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 2222 17320 2228 17332
rect 1719 17292 2228 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 4338 17320 4344 17332
rect 4172 17292 4344 17320
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 2648 17224 2697 17252
rect 2648 17212 2654 17224
rect 2685 17221 2697 17224
rect 2731 17252 2743 17255
rect 4172 17252 4200 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 10686 17280 10692 17332
rect 10744 17320 10750 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 10744 17292 11069 17320
rect 10744 17280 10750 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 11664 17292 12725 17320
rect 11664 17280 11670 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 12713 17283 12771 17289
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 17037 17323 17095 17329
rect 17037 17320 17049 17323
rect 16080 17292 17049 17320
rect 16080 17280 16086 17292
rect 17037 17289 17049 17292
rect 17083 17289 17095 17323
rect 17037 17283 17095 17289
rect 2731 17224 4200 17252
rect 4249 17255 4307 17261
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 4706 17252 4712 17264
rect 4295 17224 4712 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 4706 17212 4712 17224
rect 4764 17212 4770 17264
rect 7466 17252 7472 17264
rect 5460 17224 7472 17252
rect 3050 17184 3056 17196
rect 3011 17156 3056 17184
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 2130 17116 2136 17128
rect 1627 17088 2136 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 2682 17116 2688 17128
rect 2639 17088 2688 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 4154 17116 4160 17128
rect 2915 17088 4160 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 5460 17125 5488 17224
rect 7466 17212 7472 17224
rect 7524 17252 7530 17264
rect 7524 17224 19196 17252
rect 7524 17212 7530 17224
rect 5718 17184 5724 17196
rect 5679 17156 5724 17184
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 7742 17184 7748 17196
rect 7703 17156 7748 17184
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 8662 17184 8668 17196
rect 8623 17156 8668 17184
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 12434 17184 12440 17196
rect 10796 17156 12440 17184
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17085 5503 17119
rect 5626 17116 5632 17128
rect 5587 17088 5632 17116
rect 5445 17079 5503 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 7116 17088 7389 17116
rect 7116 16980 7144 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 7524 17088 8769 17116
rect 7524 17076 7530 17088
rect 8757 17085 8769 17088
rect 8803 17116 8815 17119
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 8803 17088 9321 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17116 9551 17119
rect 10134 17116 10140 17128
rect 9539 17088 10140 17116
rect 9539 17085 9551 17088
rect 9493 17079 9551 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10594 17116 10600 17128
rect 10376 17088 10600 17116
rect 10376 17076 10382 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10796 17125 10824 17156
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 12584 17156 14657 17184
rect 12584 17144 12590 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 19058 17184 19064 17196
rect 17552 17156 19064 17184
rect 17552 17144 17558 17156
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 12618 17116 12624 17128
rect 12579 17088 12624 17116
rect 10965 17079 11023 17085
rect 7193 17051 7251 17057
rect 7193 17017 7205 17051
rect 7239 17048 7251 17051
rect 8018 17048 8024 17060
rect 7239 17020 8024 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 9858 17048 9864 17060
rect 9819 17020 9864 17048
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 8294 16980 8300 16992
rect 7116 16952 8300 16980
rect 8294 16940 8300 16952
rect 8352 16980 8358 16992
rect 10980 16980 11008 17079
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13780 17088 14013 17116
rect 13780 17076 13786 17088
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14826 17116 14832 17128
rect 14739 17088 14832 17116
rect 14001 17079 14059 17085
rect 14826 17076 14832 17088
rect 14884 17116 14890 17128
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 14884 17088 15393 17116
rect 14884 17076 14890 17088
rect 15381 17085 15393 17088
rect 15427 17085 15439 17119
rect 15562 17116 15568 17128
rect 15523 17088 15568 17116
rect 15381 17079 15439 17085
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 15396 17048 15424 17079
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 15838 17116 15844 17128
rect 15672 17088 15844 17116
rect 15672 17048 15700 17088
rect 15838 17076 15844 17088
rect 15896 17116 15902 17128
rect 16853 17119 16911 17125
rect 15896 17088 16160 17116
rect 15896 17076 15902 17088
rect 12492 17020 12537 17048
rect 15396 17020 15700 17048
rect 15933 17051 15991 17057
rect 12492 17008 12498 17020
rect 15933 17017 15945 17051
rect 15979 17048 15991 17051
rect 16022 17048 16028 17060
rect 15979 17020 16028 17048
rect 15979 17017 15991 17020
rect 15933 17011 15991 17017
rect 16022 17008 16028 17020
rect 16080 17008 16086 17060
rect 16132 17048 16160 17088
rect 16853 17085 16865 17119
rect 16899 17116 16911 17119
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 16899 17088 18061 17116
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 18049 17085 18061 17088
rect 18095 17116 18107 17119
rect 18230 17116 18236 17128
rect 18095 17088 18236 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 19168 17125 19196 17224
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 16132 17020 18276 17048
rect 8352 16952 11008 16980
rect 8352 16940 8358 16952
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 12216 16952 13829 16980
rect 12216 16940 12222 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 17126 16980 17132 16992
rect 15620 16952 17132 16980
rect 15620 16940 15626 16952
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 18248 16989 18276 17020
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16949 18291 16983
rect 18233 16943 18291 16949
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 19245 16983 19303 16989
rect 19245 16980 19257 16983
rect 18564 16952 19257 16980
rect 18564 16940 18570 16952
rect 19245 16949 19257 16952
rect 19291 16949 19303 16983
rect 19245 16943 19303 16949
rect 1104 16890 24840 16912
rect 1104 16838 8912 16890
rect 8964 16838 8976 16890
rect 9028 16838 9040 16890
rect 9092 16838 9104 16890
rect 9156 16838 16843 16890
rect 16895 16838 16907 16890
rect 16959 16838 16971 16890
rect 17023 16838 17035 16890
rect 17087 16838 24840 16890
rect 1104 16816 24840 16838
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6454 16776 6460 16788
rect 5592 16748 6460 16776
rect 5592 16736 5598 16748
rect 6454 16736 6460 16748
rect 6512 16736 6518 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 19058 16736 19064 16788
rect 19116 16776 19122 16788
rect 19337 16779 19395 16785
rect 19337 16776 19349 16779
rect 19116 16748 19349 16776
rect 19116 16736 19122 16748
rect 19337 16745 19349 16748
rect 19383 16745 19395 16779
rect 19337 16739 19395 16745
rect 3786 16668 3792 16720
rect 3844 16708 3850 16720
rect 4522 16708 4528 16720
rect 3844 16680 4384 16708
rect 4435 16680 4528 16708
rect 3844 16668 3850 16680
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 4356 16649 4384 16680
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 1670 16572 1676 16584
rect 1631 16544 1676 16572
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 3050 16572 3056 16584
rect 2963 16544 3056 16572
rect 3050 16532 3056 16544
rect 3108 16572 3114 16584
rect 4154 16572 4160 16584
rect 3108 16544 4160 16572
rect 3108 16532 3114 16544
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4264 16572 4292 16603
rect 4448 16572 4476 16680
rect 4522 16668 4528 16680
rect 4580 16708 4586 16720
rect 4580 16680 4844 16708
rect 4580 16668 4586 16680
rect 4706 16640 4712 16652
rect 4667 16612 4712 16640
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 4816 16649 4844 16680
rect 11054 16668 11060 16720
rect 11112 16708 11118 16720
rect 11698 16708 11704 16720
rect 11112 16680 11284 16708
rect 11659 16680 11704 16708
rect 11112 16668 11118 16680
rect 4801 16643 4859 16649
rect 4801 16609 4813 16643
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16640 6331 16643
rect 6454 16640 6460 16652
rect 6319 16612 6460 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 7524 16612 7573 16640
rect 7524 16600 7530 16612
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7561 16603 7619 16609
rect 7760 16612 8125 16640
rect 4264 16544 4476 16572
rect 7377 16575 7435 16581
rect 4356 16516 4384 16544
rect 7377 16541 7389 16575
rect 7423 16541 7435 16575
rect 7576 16572 7604 16603
rect 7760 16572 7788 16612
rect 8113 16609 8125 16612
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16640 8355 16643
rect 9582 16640 9588 16652
rect 8343 16612 9588 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 8570 16572 8576 16584
rect 7576 16544 7788 16572
rect 8531 16544 8576 16572
rect 7377 16535 7435 16541
rect 4338 16464 4344 16516
rect 4396 16464 4402 16516
rect 7392 16504 7420 16535
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 10336 16572 10364 16603
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10468 16612 10701 16640
rect 10468 16600 10474 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11146 16640 11152 16652
rect 10919 16612 11152 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 11256 16640 11284 16680
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11256 16612 11897 16640
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 13081 16643 13139 16649
rect 13081 16609 13093 16643
rect 13127 16609 13139 16643
rect 13262 16640 13268 16652
rect 13223 16612 13268 16640
rect 13081 16603 13139 16609
rect 10100 16544 10364 16572
rect 13096 16572 13124 16603
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13722 16600 13728 16652
rect 13780 16640 13786 16652
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 13780 16612 14657 16640
rect 13780 16600 13786 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 15470 16640 15476 16652
rect 14645 16603 14703 16609
rect 14752 16612 15476 16640
rect 13446 16572 13452 16584
rect 13096 16544 13452 16572
rect 10100 16532 10106 16544
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 14752 16572 14780 16612
rect 15470 16600 15476 16612
rect 15528 16640 15534 16652
rect 15746 16640 15752 16652
rect 15528 16612 15752 16640
rect 15528 16600 15534 16612
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 16022 16640 16028 16652
rect 15983 16612 16028 16640
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 16172 16612 18245 16640
rect 16172 16600 16178 16612
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 19242 16640 19248 16652
rect 19203 16612 19248 16640
rect 18233 16603 18291 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 14476 16544 14780 16572
rect 8294 16504 8300 16516
rect 7392 16476 8300 16504
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 14476 16513 14504 16544
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 15620 16544 18337 16572
rect 15620 16532 15626 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16473 14519 16507
rect 14461 16467 14519 16473
rect 14642 16464 14648 16516
rect 14700 16504 14706 16516
rect 15102 16504 15108 16516
rect 14700 16476 15108 16504
rect 14700 16464 14706 16476
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 4028 16408 5273 16436
rect 4028 16396 4034 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 8570 16436 8576 16448
rect 8444 16408 8576 16436
rect 8444 16396 8450 16408
rect 8570 16396 8576 16408
rect 8628 16396 8634 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11977 16439 12035 16445
rect 11977 16436 11989 16439
rect 11020 16408 11989 16436
rect 11020 16396 11026 16408
rect 11977 16405 11989 16408
rect 12023 16405 12035 16439
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 11977 16399 12035 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14550 16436 14556 16448
rect 14332 16408 14556 16436
rect 14332 16396 14338 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 17313 16439 17371 16445
rect 17313 16436 17325 16439
rect 17000 16408 17325 16436
rect 17000 16396 17006 16408
rect 17313 16405 17325 16408
rect 17359 16436 17371 16439
rect 18414 16436 18420 16448
rect 17359 16408 18420 16436
rect 17359 16405 17371 16408
rect 17313 16399 17371 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 1104 16346 24840 16368
rect 1104 16294 4947 16346
rect 4999 16294 5011 16346
rect 5063 16294 5075 16346
rect 5127 16294 5139 16346
rect 5191 16294 12878 16346
rect 12930 16294 12942 16346
rect 12994 16294 13006 16346
rect 13058 16294 13070 16346
rect 13122 16294 20808 16346
rect 20860 16294 20872 16346
rect 20924 16294 20936 16346
rect 20988 16294 21000 16346
rect 21052 16294 24840 16346
rect 1104 16272 24840 16294
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 8260 16204 8493 16232
rect 8260 16192 8266 16204
rect 8481 16201 8493 16204
rect 8527 16201 8539 16235
rect 8481 16195 8539 16201
rect 11241 16235 11299 16241
rect 11241 16201 11253 16235
rect 11287 16232 11299 16235
rect 12250 16232 12256 16244
rect 11287 16204 12256 16232
rect 11287 16201 11299 16204
rect 11241 16195 11299 16201
rect 12250 16192 12256 16204
rect 12308 16232 12314 16244
rect 16114 16232 16120 16244
rect 12308 16204 16120 16232
rect 12308 16192 12314 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17126 16232 17132 16244
rect 17083 16204 17132 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 17586 16192 17592 16244
rect 17644 16232 17650 16244
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 17644 16204 18337 16232
rect 17644 16192 17650 16204
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18325 16195 18383 16201
rect 18693 16235 18751 16241
rect 18693 16201 18705 16235
rect 18739 16232 18751 16235
rect 19242 16232 19248 16244
rect 18739 16204 19248 16232
rect 18739 16201 18751 16204
rect 18693 16195 18751 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 2409 16167 2467 16173
rect 2409 16133 2421 16167
rect 2455 16164 2467 16167
rect 2590 16164 2596 16176
rect 2455 16136 2596 16164
rect 2455 16133 2467 16136
rect 2409 16127 2467 16133
rect 2590 16124 2596 16136
rect 2648 16124 2654 16176
rect 3970 16096 3976 16108
rect 3931 16068 3976 16096
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4154 16056 4160 16108
rect 4212 16096 4218 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 4212 16068 5089 16096
rect 4212 16056 4218 16068
rect 5077 16065 5089 16068
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 6822 16096 6828 16108
rect 6236 16068 6828 16096
rect 6236 16056 6242 16068
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9916 16068 9965 16096
rect 9916 16056 9922 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 12158 16056 12164 16108
rect 12216 16096 12222 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12216 16068 12449 16096
rect 12216 16056 12222 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 15010 16096 15016 16108
rect 12437 16059 12495 16065
rect 12636 16068 14872 16096
rect 14971 16068 15016 16096
rect 2314 16037 2320 16040
rect 2280 16031 2320 16037
rect 2280 15997 2292 16031
rect 2280 15991 2320 15997
rect 2314 15988 2320 15991
rect 2372 15988 2378 16040
rect 2498 16037 2504 16040
rect 2472 16031 2504 16037
rect 2472 16028 2484 16031
rect 2411 16000 2484 16028
rect 2472 15997 2484 16000
rect 2556 16028 2562 16040
rect 3050 16028 3056 16040
rect 2556 16000 3056 16028
rect 2472 15991 2504 15997
rect 2498 15988 2504 15991
rect 2556 15988 2562 16000
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3694 16028 3700 16040
rect 3655 16000 3700 16028
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 6362 16028 6368 16040
rect 6323 16000 6368 16028
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 7156 16000 8217 16028
rect 7156 15988 7162 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 9766 16028 9772 16040
rect 9723 16000 9772 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 2038 15920 2044 15972
rect 2096 15960 2102 15972
rect 2133 15963 2191 15969
rect 2133 15960 2145 15963
rect 2096 15932 2145 15960
rect 2096 15920 2102 15932
rect 2133 15929 2145 15932
rect 2179 15929 2191 15963
rect 2133 15923 2191 15929
rect 2869 15963 2927 15969
rect 2869 15929 2881 15963
rect 2915 15960 2927 15963
rect 2958 15960 2964 15972
rect 2915 15932 2964 15960
rect 2915 15929 2927 15932
rect 2869 15923 2927 15929
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 6825 15963 6883 15969
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7374 15960 7380 15972
rect 6871 15932 7380 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 8404 15892 8432 15991
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 12636 16028 12664 16068
rect 12308 16000 12664 16028
rect 12713 16031 12771 16037
rect 12308 15988 12314 16000
rect 12713 15997 12725 16031
rect 12759 16028 12771 16031
rect 13538 16028 13544 16040
rect 12759 16000 13544 16028
rect 12759 15997 12771 16000
rect 12713 15991 12771 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 14844 16028 14872 16068
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 16206 16096 16212 16108
rect 15948 16068 16212 16096
rect 15378 16028 15384 16040
rect 14844 16000 15384 16028
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 15565 16031 15623 16037
rect 15565 15997 15577 16031
rect 15611 16028 15623 16031
rect 15654 16028 15660 16040
rect 15611 16000 15660 16028
rect 15611 15997 15623 16000
rect 15565 15991 15623 15997
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 15948 16037 15976 16068
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 17494 16056 17500 16108
rect 17552 16096 17558 16108
rect 18196 16099 18254 16105
rect 18196 16096 18208 16099
rect 17552 16068 18208 16096
rect 17552 16056 17558 16068
rect 18196 16065 18208 16068
rect 18242 16065 18254 16099
rect 18414 16096 18420 16108
rect 18375 16068 18420 16096
rect 18196 16059 18254 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 16114 16028 16120 16040
rect 16075 16000 16120 16028
rect 15933 15991 15991 15997
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18690 16028 18696 16040
rect 18095 16000 18696 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 14093 15963 14151 15969
rect 14093 15960 14105 15963
rect 13504 15932 14105 15960
rect 13504 15920 13510 15932
rect 14093 15929 14105 15932
rect 14139 15960 14151 15963
rect 16574 15960 16580 15972
rect 14139 15932 16580 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 13170 15892 13176 15904
rect 8404 15864 13176 15892
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 1104 15802 24840 15824
rect 1104 15750 8912 15802
rect 8964 15750 8976 15802
rect 9028 15750 9040 15802
rect 9092 15750 9104 15802
rect 9156 15750 16843 15802
rect 16895 15750 16907 15802
rect 16959 15750 16971 15802
rect 17023 15750 17035 15802
rect 17087 15750 24840 15802
rect 1104 15728 24840 15750
rect 9769 15691 9827 15697
rect 9769 15688 9781 15691
rect 2240 15660 9781 15688
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 1670 15620 1676 15632
rect 1627 15592 1676 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 1670 15580 1676 15592
rect 1728 15580 1734 15632
rect 2240 15561 2268 15660
rect 9769 15657 9781 15660
rect 9815 15657 9827 15691
rect 9769 15651 9827 15657
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 14458 15688 14464 15700
rect 13495 15660 14464 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 15470 15688 15476 15700
rect 14700 15660 15476 15688
rect 14700 15648 14706 15660
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 17954 15688 17960 15700
rect 17915 15660 17960 15688
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 4709 15623 4767 15629
rect 4709 15589 4721 15623
rect 4755 15620 4767 15623
rect 5258 15620 5264 15632
rect 4755 15592 5264 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 6733 15623 6791 15629
rect 6733 15620 6745 15623
rect 6696 15592 6745 15620
rect 6696 15580 6702 15592
rect 6733 15589 6745 15592
rect 6779 15589 6791 15623
rect 6733 15583 6791 15589
rect 13832 15592 14320 15620
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2498 15512 2504 15564
rect 2556 15552 2562 15564
rect 2593 15555 2651 15561
rect 2593 15552 2605 15555
rect 2556 15524 2605 15552
rect 2556 15512 2562 15524
rect 2593 15521 2605 15524
rect 2639 15521 2651 15555
rect 2593 15515 2651 15521
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2740 15524 2789 15552
rect 2740 15512 2746 15524
rect 2777 15521 2789 15524
rect 2823 15552 2835 15555
rect 3602 15552 3608 15564
rect 2823 15524 3608 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3602 15512 3608 15524
rect 3660 15512 3666 15564
rect 4062 15512 4068 15564
rect 4120 15552 4126 15564
rect 4120 15524 5488 15552
rect 4120 15512 4126 15524
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 2406 15484 2412 15496
rect 2363 15456 2412 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4212 15456 5273 15484
rect 4212 15444 4218 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5460 15484 5488 15524
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 7190 15552 7196 15564
rect 5592 15524 5637 15552
rect 6656 15524 7196 15552
rect 5592 15512 5598 15524
rect 6656 15496 6684 15524
rect 7190 15512 7196 15524
rect 7248 15552 7254 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7248 15524 7389 15552
rect 7248 15512 7254 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 7834 15552 7840 15564
rect 7791 15524 7840 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 8386 15552 8392 15564
rect 7975 15524 8392 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 9214 15552 9220 15564
rect 9171 15524 9220 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5460 15456 5733 15484
rect 5261 15447 5319 15453
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8202 15484 8208 15496
rect 7515 15456 8208 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 2958 15376 2964 15428
rect 3016 15416 3022 15428
rect 9692 15416 9720 15515
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 10689 15555 10747 15561
rect 10689 15552 10701 15555
rect 9824 15524 10701 15552
rect 9824 15512 9830 15524
rect 10689 15521 10701 15524
rect 10735 15552 10747 15555
rect 12158 15552 12164 15564
rect 10735 15524 12164 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 13832 15561 13860 15592
rect 13817 15555 13875 15561
rect 13817 15521 13829 15555
rect 13863 15521 13875 15555
rect 13817 15515 13875 15521
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 12526 15484 12532 15496
rect 11011 15456 12532 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13906 15484 13912 15496
rect 13867 15456 13912 15484
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 3016 15388 9720 15416
rect 14200 15416 14228 15515
rect 14292 15484 14320 15592
rect 14550 15580 14556 15632
rect 14608 15620 14614 15632
rect 15289 15623 15347 15629
rect 15289 15620 15301 15623
rect 14608 15592 15301 15620
rect 14608 15580 14614 15592
rect 15289 15589 15301 15592
rect 15335 15589 15347 15623
rect 15289 15583 15347 15589
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 18969 15623 19027 15629
rect 18969 15620 18981 15623
rect 15436 15592 18981 15620
rect 15436 15580 15442 15592
rect 18969 15589 18981 15592
rect 19015 15589 19027 15623
rect 18969 15583 19027 15589
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15552 14427 15555
rect 15470 15552 15476 15564
rect 14415 15524 15476 15552
rect 14415 15521 14427 15524
rect 14369 15515 14427 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15654 15552 15660 15564
rect 15580 15524 15660 15552
rect 15580 15484 15608 15524
rect 15654 15512 15660 15524
rect 15712 15552 15718 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15712 15524 15945 15552
rect 15712 15512 15718 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 16298 15552 16304 15564
rect 16259 15524 16304 15552
rect 15933 15515 15991 15521
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 17313 15555 17371 15561
rect 17313 15552 17325 15555
rect 16724 15524 17325 15552
rect 16724 15512 16730 15524
rect 17313 15521 17325 15524
rect 17359 15521 17371 15555
rect 18877 15555 18935 15561
rect 18877 15552 18889 15555
rect 17313 15515 17371 15521
rect 17420 15524 18889 15552
rect 15746 15484 15752 15496
rect 14292 15456 15608 15484
rect 15707 15456 15752 15484
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 16206 15484 16212 15496
rect 16167 15456 16212 15484
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 16316 15416 16344 15512
rect 14200 15388 16344 15416
rect 3016 15376 3022 15388
rect 8941 15351 8999 15357
rect 8941 15317 8953 15351
rect 8987 15348 8999 15351
rect 9214 15348 9220 15360
rect 8987 15320 9220 15348
rect 8987 15317 8999 15320
rect 8941 15311 8999 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12434 15348 12440 15360
rect 12299 15320 12440 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12434 15308 12440 15320
rect 12492 15348 12498 15360
rect 17420 15348 17448 15524
rect 18877 15521 18889 15524
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 18138 15484 18144 15496
rect 17727 15456 18144 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 18138 15444 18144 15456
rect 18196 15484 18202 15496
rect 18414 15484 18420 15496
rect 18196 15456 18420 15484
rect 18196 15444 18202 15456
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 17494 15425 17500 15428
rect 17478 15419 17500 15425
rect 17478 15385 17490 15419
rect 17478 15379 17500 15385
rect 17494 15376 17500 15379
rect 17552 15376 17558 15428
rect 17586 15348 17592 15360
rect 12492 15320 17448 15348
rect 17547 15320 17592 15348
rect 12492 15308 12498 15320
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 1104 15258 24840 15280
rect 1104 15206 4947 15258
rect 4999 15206 5011 15258
rect 5063 15206 5075 15258
rect 5127 15206 5139 15258
rect 5191 15206 12878 15258
rect 12930 15206 12942 15258
rect 12994 15206 13006 15258
rect 13058 15206 13070 15258
rect 13122 15206 20808 15258
rect 20860 15206 20872 15258
rect 20924 15206 20936 15258
rect 20988 15206 21000 15258
rect 21052 15206 24840 15258
rect 1104 15184 24840 15206
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 5442 15144 5448 15156
rect 5316 15116 5448 15144
rect 5316 15104 5322 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 19153 15147 19211 15153
rect 19153 15144 19165 15147
rect 8260 15116 19165 15144
rect 8260 15104 8266 15116
rect 19153 15113 19165 15116
rect 19199 15113 19211 15147
rect 19153 15107 19211 15113
rect 3602 15036 3608 15088
rect 3660 15076 3666 15088
rect 3660 15048 4200 15076
rect 3660 15036 3666 15048
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 15008 2283 15011
rect 2682 15008 2688 15020
rect 2271 14980 2688 15008
rect 2271 14977 2283 14980
rect 2225 14971 2283 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3142 15008 3148 15020
rect 3103 14980 3148 15008
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 4172 15008 4200 15048
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 9585 15079 9643 15085
rect 9585 15076 9597 15079
rect 8628 15048 9597 15076
rect 8628 15036 8634 15048
rect 9585 15045 9597 15048
rect 9631 15045 9643 15079
rect 13538 15076 13544 15088
rect 13499 15048 13544 15076
rect 9585 15039 9643 15045
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 15746 15076 15752 15088
rect 14752 15048 15752 15076
rect 4172 14980 11376 15008
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2498 14940 2504 14952
rect 1903 14912 2504 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2498 14900 2504 14912
rect 2556 14900 2562 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 3237 14943 3295 14949
rect 3237 14940 3249 14943
rect 2832 14912 3249 14940
rect 2832 14900 2838 14912
rect 3237 14909 3249 14912
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14909 3755 14943
rect 3697 14903 3755 14909
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 3970 14940 3976 14952
rect 3835 14912 3976 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 1762 14872 1768 14884
rect 1719 14844 1768 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 1762 14832 1768 14844
rect 1820 14872 1826 14884
rect 2590 14872 2596 14884
rect 1820 14844 2596 14872
rect 1820 14832 1826 14844
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 3712 14872 3740 14903
rect 3970 14900 3976 14912
rect 4028 14940 4034 14952
rect 4338 14940 4344 14952
rect 4028 14912 4344 14940
rect 4028 14900 4034 14912
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 5258 14940 5264 14952
rect 4672 14912 5264 14940
rect 4672 14900 4678 14912
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 5960 14912 6837 14940
rect 5960 14900 5966 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 8570 14940 8576 14952
rect 7147 14912 8576 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 9766 14940 9772 14952
rect 9727 14912 9772 14940
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10042 14940 10048 14952
rect 9999 14912 10048 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10410 14940 10416 14952
rect 10367 14912 10416 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10870 14940 10876 14952
rect 10551 14912 10876 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11348 14949 11376 14980
rect 12590 14980 12848 15008
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 12590 14949 12618 14980
rect 12575 14943 12633 14949
rect 12575 14940 12587 14943
rect 12216 14912 12587 14940
rect 12216 14900 12222 14912
rect 12575 14909 12587 14912
rect 12621 14909 12633 14943
rect 12710 14940 12716 14952
rect 12671 14912 12716 14940
rect 12575 14903 12633 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 12820 14940 12848 14980
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 13688 14980 14657 15008
rect 13688 14968 13694 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 12820 14912 13185 14940
rect 13173 14909 13185 14912
rect 13219 14940 13231 14943
rect 13262 14940 13268 14952
rect 13219 14912 13268 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14940 13415 14943
rect 14752 14940 14780 15048
rect 15746 15036 15752 15048
rect 15804 15076 15810 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 15804 15048 16957 15076
rect 15804 15036 15810 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 13403 14912 14780 14940
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 14884 14912 15393 14940
rect 14884 14900 14890 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 15746 14940 15752 14952
rect 15611 14912 15752 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16632 14912 16865 14940
rect 16632 14900 16638 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 18012 14912 18061 14940
rect 18012 14900 18018 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 4062 14872 4068 14884
rect 3712 14844 4068 14872
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14872 8539 14875
rect 9674 14872 9680 14884
rect 8527 14844 9680 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 9674 14832 9680 14844
rect 9732 14872 9738 14884
rect 19076 14872 19104 14903
rect 9732 14844 19104 14872
rect 9732 14832 9738 14844
rect 3234 14764 3240 14816
rect 3292 14804 3298 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3292 14776 4261 14804
rect 3292 14764 3298 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 4249 14767 4307 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 11422 14804 11428 14816
rect 11383 14776 11428 14804
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 14642 14804 14648 14816
rect 11756 14776 14648 14804
rect 11756 14764 11762 14776
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15620 14776 15853 14804
rect 15620 14764 15626 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 18104 14776 18153 14804
rect 18104 14764 18110 14776
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18141 14767 18199 14773
rect 1104 14714 24840 14736
rect 1104 14662 8912 14714
rect 8964 14662 8976 14714
rect 9028 14662 9040 14714
rect 9092 14662 9104 14714
rect 9156 14662 16843 14714
rect 16895 14662 16907 14714
rect 16959 14662 16971 14714
rect 17023 14662 17035 14714
rect 17087 14662 24840 14714
rect 1104 14640 24840 14662
rect 11422 14600 11428 14612
rect 2148 14572 11428 14600
rect 2148 14473 2176 14572
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 11940 14572 15148 14600
rect 11940 14560 11946 14572
rect 2222 14492 2228 14544
rect 2280 14532 2286 14544
rect 4062 14532 4068 14544
rect 2280 14504 4068 14532
rect 2280 14492 2286 14504
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 8570 14532 8576 14544
rect 8531 14504 8576 14532
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8846 14492 8852 14544
rect 8904 14532 8910 14544
rect 12158 14532 12164 14544
rect 8904 14504 11376 14532
rect 8904 14492 8910 14504
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14433 2191 14467
rect 2498 14464 2504 14476
rect 2459 14436 2504 14464
rect 2133 14427 2191 14433
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14464 7527 14467
rect 7926 14464 7932 14476
rect 7515 14436 7932 14464
rect 7515 14433 7527 14436
rect 7469 14427 7527 14433
rect 7926 14424 7932 14436
rect 7984 14464 7990 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7984 14436 8033 14464
rect 7984 14424 7990 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8021 14427 8079 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 11238 14464 11244 14476
rect 11199 14436 11244 14464
rect 9677 14427 9735 14433
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2406 14396 2412 14408
rect 2271 14368 2412 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2590 14396 2596 14408
rect 2551 14368 2596 14396
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 3694 14396 3700 14408
rect 3016 14368 3700 14396
rect 3016 14356 3022 14368
rect 3694 14356 3700 14368
rect 3752 14396 3758 14408
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 3752 14368 4813 14396
rect 3752 14356 3758 14368
rect 4801 14365 4813 14368
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5258 14396 5264 14408
rect 5123 14368 5264 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 5902 14288 5908 14340
rect 5960 14328 5966 14340
rect 9692 14328 9720 14427
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 11348 14464 11376 14504
rect 12084 14504 12164 14532
rect 11422 14464 11428 14476
rect 11335 14436 11428 14464
rect 11422 14424 11428 14436
rect 11480 14473 11486 14476
rect 11480 14467 11529 14473
rect 11480 14433 11483 14467
rect 11517 14433 11529 14467
rect 11606 14464 11612 14476
rect 11567 14436 11612 14464
rect 11480 14427 11529 14433
rect 11480 14424 11486 14427
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12084 14473 12112 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 13722 14532 13728 14544
rect 12952 14504 13728 14532
rect 12952 14492 12958 14504
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 15120 14532 15148 14572
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15746 14600 15752 14612
rect 15252 14572 15752 14600
rect 15252 14560 15258 14572
rect 15746 14560 15752 14572
rect 15804 14600 15810 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 15804 14572 15853 14600
rect 15804 14560 15810 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 15654 14532 15660 14544
rect 15120 14504 15660 14532
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 12069 14467 12127 14473
rect 12069 14433 12081 14467
rect 12115 14433 12127 14467
rect 12250 14464 12256 14476
rect 12211 14436 12256 14464
rect 12069 14427 12127 14433
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16850 14464 16856 14476
rect 15795 14436 16856 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 5960 14300 9720 14328
rect 11057 14331 11115 14337
rect 5960 14288 5966 14300
rect 11057 14297 11069 14331
rect 11103 14328 11115 14331
rect 12894 14328 12900 14340
rect 11103 14300 12900 14328
rect 11103 14297 11115 14300
rect 11057 14291 11115 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13556 14328 13584 14427
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 15286 14356 15292 14408
rect 15344 14396 15350 14408
rect 15838 14396 15844 14408
rect 15344 14368 15844 14396
rect 15344 14356 15350 14368
rect 15838 14356 15844 14368
rect 15896 14396 15902 14408
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 15896 14368 16773 14396
rect 15896 14356 15902 14368
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17126 14396 17132 14408
rect 17083 14368 17132 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 13004 14300 13584 14328
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 1670 14260 1676 14272
rect 1627 14232 1676 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 5442 14260 5448 14272
rect 2740 14232 5448 14260
rect 2740 14220 2746 14232
rect 5442 14220 5448 14232
rect 5500 14260 5506 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5500 14232 6193 14260
rect 5500 14220 5506 14232
rect 6181 14229 6193 14232
rect 6227 14260 6239 14263
rect 6822 14260 6828 14272
rect 6227 14232 6828 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 7984 14232 9873 14260
rect 7984 14220 7990 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 9861 14223 9919 14229
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 13004 14260 13032 14300
rect 13630 14260 13636 14272
rect 10008 14232 13032 14260
rect 13591 14232 13636 14260
rect 10008 14220 10014 14232
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 17862 14260 17868 14272
rect 13964 14232 17868 14260
rect 13964 14220 13970 14232
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18138 14260 18144 14272
rect 18012 14232 18144 14260
rect 18012 14220 18018 14232
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 1104 14170 24840 14192
rect 1104 14118 4947 14170
rect 4999 14118 5011 14170
rect 5063 14118 5075 14170
rect 5127 14118 5139 14170
rect 5191 14118 12878 14170
rect 12930 14118 12942 14170
rect 12994 14118 13006 14170
rect 13058 14118 13070 14170
rect 13122 14118 20808 14170
rect 20860 14118 20872 14170
rect 20924 14118 20936 14170
rect 20988 14118 21000 14170
rect 21052 14118 24840 14170
rect 1104 14096 24840 14118
rect 2041 14059 2099 14065
rect 2041 14025 2053 14059
rect 2087 14056 2099 14059
rect 3970 14056 3976 14068
rect 2087 14028 3976 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 7064 14028 7113 14056
rect 7064 14016 7070 14028
rect 7101 14025 7113 14028
rect 7147 14056 7159 14059
rect 9950 14056 9956 14068
rect 7147 14028 9956 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 11238 14056 11244 14068
rect 10643 14028 11244 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11425 14059 11483 14065
rect 11425 14025 11437 14059
rect 11471 14056 11483 14059
rect 11698 14056 11704 14068
rect 11471 14028 11704 14056
rect 11471 14025 11483 14028
rect 11425 14019 11483 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12342 14056 12348 14068
rect 12032 14028 12348 14056
rect 12032 14016 12038 14028
rect 12342 14016 12348 14028
rect 12400 14056 12406 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12400 14028 12725 14056
rect 12400 14016 12406 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 19153 14059 19211 14065
rect 19153 14056 19165 14059
rect 12713 14019 12771 14025
rect 15304 14028 19165 14056
rect 5813 13991 5871 13997
rect 5813 13957 5825 13991
rect 5859 13988 5871 13991
rect 7466 13988 7472 14000
rect 5859 13960 7472 13988
rect 5859 13957 5871 13960
rect 5813 13951 5871 13957
rect 7466 13948 7472 13960
rect 7524 13988 7530 14000
rect 7524 13960 8616 13988
rect 7524 13948 7530 13960
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3234 13920 3240 13932
rect 3195 13892 3240 13920
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4120 13892 4353 13920
rect 4120 13880 4126 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 5902 13920 5908 13932
rect 4341 13883 4399 13889
rect 5644 13892 5908 13920
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13852 1915 13855
rect 2774 13852 2780 13864
rect 1903 13824 2780 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 2774 13812 2780 13824
rect 2832 13852 2838 13864
rect 3970 13852 3976 13864
rect 2832 13824 3976 13852
rect 2832 13812 2838 13824
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 5644 13861 5672 13892
rect 5902 13880 5908 13892
rect 5960 13880 5966 13932
rect 6822 13920 6828 13932
rect 6783 13892 6828 13920
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 7926 13880 7932 13932
rect 7984 13920 7990 13932
rect 7984 13892 8524 13920
rect 7984 13880 7990 13892
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6604 13824 6929 13852
rect 6604 13812 6610 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7742 13812 7748 13864
rect 7800 13852 7806 13864
rect 8496 13861 8524 13892
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7800 13824 8309 13852
rect 7800 13812 7806 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8481 13855 8539 13861
rect 8481 13821 8493 13855
rect 8527 13821 8539 13855
rect 8588 13852 8616 13960
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 9272 13960 10517 13988
rect 9272 13948 9278 13960
rect 10505 13957 10517 13960
rect 10551 13957 10563 13991
rect 11256 13988 11284 14016
rect 12526 13988 12532 14000
rect 11256 13960 12532 13988
rect 10505 13951 10563 13957
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 13354 13948 13360 14000
rect 13412 13988 13418 14000
rect 13817 13991 13875 13997
rect 13817 13988 13829 13991
rect 13412 13960 13829 13988
rect 13412 13948 13418 13960
rect 13817 13957 13829 13960
rect 13863 13957 13875 13991
rect 13817 13951 13875 13957
rect 15304 13920 15332 14028
rect 19153 14025 19165 14028
rect 19199 14025 19211 14059
rect 19153 14019 19211 14025
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18141 13991 18199 13997
rect 18141 13988 18153 13991
rect 17920 13960 18153 13988
rect 17920 13948 17926 13960
rect 18141 13957 18153 13960
rect 18187 13957 18199 13991
rect 18141 13951 18199 13957
rect 15562 13920 15568 13932
rect 10336 13892 15332 13920
rect 15523 13892 15568 13920
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8588 13824 9045 13852
rect 8481 13815 8539 13821
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9766 13852 9772 13864
rect 9263 13824 9772 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9766 13812 9772 13824
rect 9824 13852 9830 13864
rect 10336 13852 10364 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 15712 13892 19104 13920
rect 15712 13880 15718 13892
rect 9824 13824 10364 13852
rect 10505 13855 10563 13861
rect 9824 13812 9830 13824
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10551 13824 10793 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 11241 13855 11299 13861
rect 11241 13821 11253 13855
rect 11287 13852 11299 13855
rect 11330 13852 11336 13864
rect 11287 13824 11336 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 12529 13855 12587 13861
rect 11480 13824 12480 13852
rect 11480 13812 11486 13824
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 8846 13784 8852 13796
rect 8260 13756 8852 13784
rect 8260 13744 8266 13756
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 9582 13784 9588 13796
rect 9543 13756 9588 13784
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 12452 13784 12480 13824
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 13170 13852 13176 13864
rect 12575 13824 13176 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13633 13855 13691 13861
rect 13633 13852 13645 13855
rect 13280 13824 13645 13852
rect 13280 13784 13308 13824
rect 13633 13821 13645 13824
rect 13679 13852 13691 13855
rect 13679 13824 15240 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 12452 13756 13308 13784
rect 15212 13784 15240 13824
rect 15286 13812 15292 13864
rect 15344 13852 15350 13864
rect 15344 13824 15389 13852
rect 16224 13824 16804 13852
rect 15344 13812 15350 13824
rect 15378 13784 15384 13796
rect 15212 13756 15384 13784
rect 15378 13744 15384 13756
rect 15436 13744 15442 13796
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12158 13716 12164 13728
rect 11848 13688 12164 13716
rect 11848 13676 11854 13688
rect 12158 13676 12164 13688
rect 12216 13716 12222 13728
rect 13722 13716 13728 13728
rect 12216 13688 13728 13716
rect 12216 13676 12222 13688
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 16224 13716 16252 13824
rect 16776 13784 16804 13824
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16908 13824 16957 13852
rect 16908 13812 16914 13824
rect 16945 13821 16957 13824
rect 16991 13852 17003 13855
rect 17862 13852 17868 13864
rect 16991 13824 17868 13852
rect 16991 13821 17003 13824
rect 16945 13815 17003 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 19076 13861 19104 13892
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17972 13824 18061 13852
rect 17972 13784 18000 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 16776 13756 18000 13784
rect 14424 13688 16252 13716
rect 14424 13676 14430 13688
rect 1104 13626 24840 13648
rect 1104 13574 8912 13626
rect 8964 13574 8976 13626
rect 9028 13574 9040 13626
rect 9092 13574 9104 13626
rect 9156 13574 16843 13626
rect 16895 13574 16907 13626
rect 16959 13574 16971 13626
rect 17023 13574 17035 13626
rect 17087 13574 24840 13626
rect 1104 13552 24840 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2777 13515 2835 13521
rect 2777 13512 2789 13515
rect 2556 13484 2789 13512
rect 2556 13472 2562 13484
rect 2777 13481 2789 13484
rect 2823 13481 2835 13515
rect 6086 13512 6092 13524
rect 2777 13475 2835 13481
rect 4632 13484 5396 13512
rect 6047 13484 6092 13512
rect 4632 13453 4660 13484
rect 4617 13447 4675 13453
rect 4617 13413 4629 13447
rect 4663 13413 4675 13447
rect 4617 13407 4675 13413
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 5258 13444 5264 13456
rect 5215 13416 5264 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 5368 13444 5396 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 13630 13512 13636 13524
rect 8496 13484 13636 13512
rect 8496 13444 8524 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 18506 13512 18512 13524
rect 13740 13484 18512 13512
rect 5368 13416 8524 13444
rect 11333 13447 11391 13453
rect 11333 13413 11345 13447
rect 11379 13444 11391 13447
rect 11882 13444 11888 13456
rect 11379 13416 11888 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5534 13376 5540 13388
rect 4755 13348 5540 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6638 13376 6644 13388
rect 6599 13348 6644 13376
rect 6638 13336 6644 13348
rect 6696 13336 6702 13388
rect 7006 13385 7012 13388
rect 6980 13379 7012 13385
rect 6980 13376 6992 13379
rect 6919 13348 6992 13376
rect 6980 13345 6992 13348
rect 7064 13376 7070 13388
rect 7193 13379 7251 13385
rect 7064 13348 7144 13376
rect 6980 13339 7012 13345
rect 7006 13336 7012 13339
rect 7064 13336 7070 13348
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 5810 13308 5816 13320
rect 4479 13280 5816 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 5552 13252 5580 13280
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6236 13280 6469 13308
rect 6236 13268 6242 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 7116 13308 7144 13348
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 7466 13376 7472 13388
rect 7239 13348 7472 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 7466 13336 7472 13348
rect 7524 13376 7530 13388
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7524 13348 8033 13376
rect 7524 13336 7530 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9640 13348 9965 13376
rect 9640 13336 9646 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13376 12219 13379
rect 13630 13376 13636 13388
rect 12207 13348 13636 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 7834 13308 7840 13320
rect 7116 13280 7840 13308
rect 6457 13271 6515 13277
rect 7834 13268 7840 13280
rect 7892 13308 7898 13320
rect 8110 13308 8116 13320
rect 7892 13280 8116 13308
rect 7892 13268 7898 13280
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13308 8450 13320
rect 9214 13308 9220 13320
rect 8444 13280 9220 13308
rect 8444 13268 8450 13280
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 9916 13280 12449 13308
rect 9916 13268 9922 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 13740 13308 13768 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 15286 13444 15292 13456
rect 15199 13416 15292 13444
rect 15286 13404 15292 13416
rect 15344 13444 15350 13456
rect 16114 13444 16120 13456
rect 15344 13416 16120 13444
rect 15344 13404 15350 13416
rect 16114 13404 16120 13416
rect 16172 13444 16178 13456
rect 16482 13444 16488 13456
rect 16172 13416 16488 13444
rect 16172 13404 16178 13416
rect 16482 13404 16488 13416
rect 16540 13404 16546 13456
rect 16945 13447 17003 13453
rect 16945 13413 16957 13447
rect 16991 13444 17003 13447
rect 17126 13444 17132 13456
rect 16991 13416 17132 13444
rect 16991 13413 17003 13416
rect 16945 13407 17003 13413
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 18046 13444 18052 13456
rect 17604 13416 18052 13444
rect 15436 13379 15494 13385
rect 15436 13345 15448 13379
rect 15482 13376 15494 13379
rect 16206 13376 16212 13388
rect 15482 13348 16212 13376
rect 15482 13345 15494 13348
rect 15436 13339 15494 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 17604 13385 17632 13416
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17678 13336 17684 13388
rect 17736 13376 17742 13388
rect 17954 13376 17960 13388
rect 17736 13348 17781 13376
rect 17915 13348 17960 13376
rect 17736 13336 17742 13348
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13376 18199 13379
rect 18966 13376 18972 13388
rect 18187 13348 18972 13376
rect 18187 13345 18199 13348
rect 18141 13339 18199 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 12437 13271 12495 13277
rect 13096 13280 13768 13308
rect 15657 13311 15715 13317
rect 5534 13200 5540 13252
rect 5592 13200 5598 13252
rect 5644 13212 8800 13240
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 5644 13172 5672 13212
rect 4764 13144 5672 13172
rect 4764 13132 4770 13144
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8159 13175 8217 13181
rect 8159 13172 8171 13175
rect 7892 13144 8171 13172
rect 7892 13132 7898 13144
rect 8159 13141 8171 13144
rect 8205 13141 8217 13175
rect 8159 13135 8217 13141
rect 8297 13175 8355 13181
rect 8297 13141 8309 13175
rect 8343 13172 8355 13175
rect 8386 13172 8392 13184
rect 8343 13144 8392 13172
rect 8343 13141 8355 13144
rect 8297 13135 8355 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8772 13172 8800 13212
rect 10612 13212 11192 13240
rect 10612 13172 10640 13212
rect 8772 13144 10640 13172
rect 11164 13172 11192 13212
rect 13096 13172 13124 13280
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15746 13308 15752 13320
rect 15703 13280 15752 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 13170 13200 13176 13252
rect 13228 13240 13234 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 13228 13212 13737 13240
rect 13228 13200 13234 13212
rect 13725 13209 13737 13212
rect 13771 13240 13783 13243
rect 16298 13240 16304 13252
rect 13771 13212 16304 13240
rect 13771 13209 13783 13212
rect 13725 13203 13783 13209
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 11164 13144 13124 13172
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 15378 13172 15384 13184
rect 13688 13144 15384 13172
rect 13688 13132 13694 13144
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 15565 13175 15623 13181
rect 15565 13172 15577 13175
rect 15528 13144 15577 13172
rect 15528 13132 15534 13144
rect 15565 13141 15577 13144
rect 15611 13141 15623 13175
rect 15565 13135 15623 13141
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 15749 13175 15807 13181
rect 15749 13172 15761 13175
rect 15712 13144 15761 13172
rect 15712 13132 15718 13144
rect 15749 13141 15761 13144
rect 15795 13141 15807 13175
rect 15749 13135 15807 13141
rect 1104 13082 24840 13104
rect 1104 13030 4947 13082
rect 4999 13030 5011 13082
rect 5063 13030 5075 13082
rect 5127 13030 5139 13082
rect 5191 13030 12878 13082
rect 12930 13030 12942 13082
rect 12994 13030 13006 13082
rect 13058 13030 13070 13082
rect 13122 13030 20808 13082
rect 20860 13030 20872 13082
rect 20924 13030 20936 13082
rect 20988 13030 21000 13082
rect 21052 13030 24840 13082
rect 1104 13008 24840 13030
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6420 12940 6469 12968
rect 6420 12928 6426 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 6457 12931 6515 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 11425 12971 11483 12977
rect 11425 12937 11437 12971
rect 11471 12968 11483 12971
rect 13446 12968 13452 12980
rect 11471 12940 13452 12968
rect 11471 12937 11483 12940
rect 11425 12931 11483 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 13780 12940 19288 12968
rect 13780 12928 13786 12940
rect 9858 12900 9864 12912
rect 4172 12872 9864 12900
rect 3326 12832 3332 12844
rect 1412 12804 3188 12832
rect 3287 12804 3332 12832
rect 1412 12773 1440 12804
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 1627 12736 2973 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 2961 12733 2973 12736
rect 3007 12764 3019 12767
rect 3050 12764 3056 12776
rect 3007 12736 3056 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 3160 12764 3188 12804
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 4172 12841 4200 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 14366 12900 14372 12912
rect 14327 12872 14372 12900
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 18141 12903 18199 12909
rect 18141 12900 18153 12903
rect 16540 12872 18153 12900
rect 16540 12860 16546 12872
rect 18141 12869 18153 12872
rect 18187 12869 18199 12903
rect 18141 12863 18199 12869
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4706 12832 4712 12844
rect 4304 12804 4712 12832
rect 4304 12792 4310 12804
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 5166 12832 5172 12844
rect 4816 12804 5172 12832
rect 4816 12764 4844 12804
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 8478 12832 8484 12844
rect 5684 12804 6868 12832
rect 8439 12804 8484 12832
rect 5684 12792 5690 12804
rect 6840 12773 6868 12804
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 10042 12832 10048 12844
rect 9048 12804 10048 12832
rect 3160 12736 4844 12764
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12733 5043 12767
rect 4985 12727 5043 12733
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 8938 12764 8944 12776
rect 6825 12727 6883 12733
rect 8404 12736 8944 12764
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 2498 12696 2504 12708
rect 1995 12668 2504 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 4154 12696 4160 12708
rect 2832 12668 4160 12696
rect 2832 12656 2838 12668
rect 4154 12656 4160 12668
rect 4212 12656 4218 12708
rect 5000 12696 5028 12727
rect 5258 12696 5264 12708
rect 5000 12668 5264 12696
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 6656 12696 6684 12727
rect 8404 12696 8432 12736
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9048 12773 9076 12804
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 15764 12804 19165 12832
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 10778 12764 10784 12776
rect 9631 12736 10784 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 6656 12668 8432 12696
rect 8846 12656 8852 12708
rect 8904 12656 8910 12708
rect 9416 12696 9444 12727
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11330 12764 11336 12776
rect 11287 12736 11336 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12492 12736 13001 12764
rect 12492 12724 12498 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 13262 12764 13268 12776
rect 13223 12736 13268 12764
rect 12989 12727 13047 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 10410 12696 10416 12708
rect 9416 12668 10416 12696
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 15764 12696 15792 12804
rect 19153 12801 19165 12804
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16298 12764 16304 12776
rect 16259 12736 16304 12764
rect 16025 12727 16083 12733
rect 14292 12668 15792 12696
rect 16040 12696 16068 12727
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16577 12767 16635 12773
rect 16577 12733 16589 12767
rect 16623 12764 16635 12767
rect 16666 12764 16672 12776
rect 16623 12736 16672 12764
rect 16623 12733 16635 12736
rect 16577 12727 16635 12733
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17184 12736 18061 12764
rect 17184 12724 17190 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 19061 12767 19119 12773
rect 19061 12733 19073 12767
rect 19107 12764 19119 12767
rect 19260 12764 19288 12940
rect 19107 12736 19288 12764
rect 19107 12733 19119 12736
rect 19061 12727 19119 12733
rect 18322 12696 18328 12708
rect 16040 12668 18328 12696
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 8864 12628 8892 12656
rect 14292 12628 14320 12668
rect 18322 12656 18328 12668
rect 18380 12656 18386 12708
rect 8536 12600 14320 12628
rect 8536 12588 8542 12600
rect 1104 12538 24840 12560
rect 1104 12486 8912 12538
rect 8964 12486 8976 12538
rect 9028 12486 9040 12538
rect 9092 12486 9104 12538
rect 9156 12486 16843 12538
rect 16895 12486 16907 12538
rect 16959 12486 16971 12538
rect 17023 12486 17035 12538
rect 17087 12486 24840 12538
rect 1104 12464 24840 12486
rect 1489 12427 1547 12433
rect 1489 12393 1501 12427
rect 1535 12424 1547 12427
rect 2222 12424 2228 12436
rect 1535 12396 2228 12424
rect 1535 12393 1547 12396
rect 1489 12387 1547 12393
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 2372 12396 4261 12424
rect 2372 12384 2378 12396
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2409 12359 2467 12365
rect 2409 12356 2421 12359
rect 2096 12328 2421 12356
rect 2096 12316 2102 12328
rect 2409 12325 2421 12328
rect 2455 12325 2467 12359
rect 2409 12319 2467 12325
rect 2608 12297 2636 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 4448 12396 13216 12424
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 4448 12356 4476 12396
rect 3476 12328 4476 12356
rect 3476 12316 3482 12328
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 5353 12359 5411 12365
rect 5353 12356 5365 12359
rect 4580 12328 5365 12356
rect 4580 12316 4586 12328
rect 5353 12325 5365 12328
rect 5399 12325 5411 12359
rect 6638 12356 6644 12368
rect 5353 12319 5411 12325
rect 6012 12328 6644 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12257 1455 12291
rect 1397 12251 1455 12257
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12257 2651 12291
rect 4062 12288 4068 12300
rect 3975 12260 4068 12288
rect 2593 12251 2651 12257
rect 1412 12220 1440 12251
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 6012 12297 6040 12328
rect 6638 12316 6644 12328
rect 6696 12356 6702 12368
rect 6914 12356 6920 12368
rect 6696 12328 6920 12356
rect 6696 12316 6702 12328
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 10962 12356 10968 12368
rect 10796 12328 10968 12356
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12288 6423 12291
rect 7006 12288 7012 12300
rect 6411 12260 7012 12288
rect 6411 12257 6423 12260
rect 6365 12251 6423 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 7926 12288 7932 12300
rect 7607 12260 7932 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7926 12248 7932 12260
rect 7984 12288 7990 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7984 12260 8125 12288
rect 7984 12248 7990 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12288 8355 12291
rect 8478 12288 8484 12300
rect 8343 12260 8484 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 8720 12260 10333 12288
rect 8720 12248 8726 12260
rect 10321 12257 10333 12260
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 2774 12220 2780 12232
rect 1412 12192 2780 12220
rect 2774 12180 2780 12192
rect 2832 12220 2838 12232
rect 4080 12220 4108 12248
rect 2832 12192 4108 12220
rect 2832 12180 2838 12192
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5776 12192 5825 12220
rect 5776 12180 5782 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7650 12220 7656 12232
rect 7515 12192 7656 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 6288 12152 6316 12183
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7926 12152 7932 12164
rect 6288 12124 7932 12152
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 8478 12152 8484 12164
rect 8439 12124 8484 12152
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 2590 12084 2596 12096
rect 1452 12056 2596 12084
rect 1452 12044 1458 12056
rect 2590 12044 2596 12056
rect 2648 12084 2654 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2648 12056 2697 12084
rect 2648 12044 2654 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2685 12047 2743 12053
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 9582 12084 9588 12096
rect 5500 12056 9588 12084
rect 5500 12044 5506 12056
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10796 12084 10824 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 12526 12316 12532 12368
rect 12584 12316 12590 12368
rect 13188 12356 13216 12396
rect 13262 12384 13268 12436
rect 13320 12424 13326 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13320 12396 13737 12424
rect 13320 12384 13326 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 18322 12424 18328 12436
rect 13725 12387 13783 12393
rect 13832 12396 18328 12424
rect 13832 12356 13860 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19061 12359 19119 12365
rect 19061 12356 19073 12359
rect 13188 12328 13860 12356
rect 17604 12328 19073 12356
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 11054 12288 11060 12300
rect 10919 12260 11060 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 12342 12288 12348 12300
rect 11287 12260 12348 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12544 12288 12572 12316
rect 12483 12260 12572 12288
rect 12713 12291 12771 12297
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 12759 12260 13277 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13265 12257 13277 12260
rect 13311 12288 13323 12291
rect 13354 12288 13360 12300
rect 13311 12260 13360 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 13906 12288 13912 12300
rect 13495 12260 13912 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 17126 12288 17132 12300
rect 15887 12260 17132 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17604 12297 17632 12328
rect 19061 12325 19073 12328
rect 19107 12325 19119 12359
rect 19061 12319 19119 12325
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 17862 12248 17868 12300
rect 17920 12288 17926 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17920 12260 17969 12288
rect 17920 12248 17926 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 18966 12288 18972 12300
rect 18927 12260 18972 12288
rect 17957 12251 18015 12257
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 11514 12220 11520 12232
rect 11471 12192 11520 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12636 12152 12664 12183
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 16724 12192 17509 12220
rect 16724 12180 16730 12192
rect 17497 12189 17509 12192
rect 17543 12220 17555 12223
rect 17678 12220 17684 12232
rect 17543 12192 17684 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 13722 12152 13728 12164
rect 12636 12124 13728 12152
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 17586 12152 17592 12164
rect 16071 12124 17592 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 17954 12112 17960 12164
rect 18012 12152 18018 12164
rect 18064 12152 18092 12183
rect 18012 12124 18092 12152
rect 18012 12112 18018 12124
rect 10870 12084 10876 12096
rect 10796 12056 10876 12084
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 12250 12084 12256 12096
rect 12211 12056 12256 12084
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 17037 12087 17095 12093
rect 17037 12053 17049 12087
rect 17083 12084 17095 12087
rect 18046 12084 18052 12096
rect 17083 12056 18052 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 1104 11994 24840 12016
rect 1104 11942 4947 11994
rect 4999 11942 5011 11994
rect 5063 11942 5075 11994
rect 5127 11942 5139 11994
rect 5191 11942 12878 11994
rect 12930 11942 12942 11994
rect 12994 11942 13006 11994
rect 13058 11942 13070 11994
rect 13122 11942 20808 11994
rect 20860 11942 20872 11994
rect 20924 11942 20936 11994
rect 20988 11942 21000 11994
rect 21052 11942 24840 11994
rect 1104 11920 24840 11942
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10928 11852 10977 11880
rect 10928 11840 10934 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 11112 11852 11161 11880
rect 11112 11840 11118 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 17310 11880 17316 11892
rect 11149 11843 11207 11849
rect 16500 11852 17316 11880
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 4120 11784 4353 11812
rect 4120 11772 4126 11784
rect 4341 11781 4353 11784
rect 4387 11812 4399 11815
rect 6546 11812 6552 11824
rect 4387 11784 6552 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 6546 11772 6552 11784
rect 6604 11812 6610 11824
rect 6822 11812 6828 11824
rect 6604 11784 6828 11812
rect 6604 11772 6610 11784
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 12342 11812 12348 11824
rect 9640 11784 12348 11812
rect 9640 11772 9646 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 16500 11821 16528 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19024 11852 19717 11880
rect 19024 11840 19030 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11781 16543 11815
rect 16485 11775 16543 11781
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 17218 11812 17224 11824
rect 16632 11784 17224 11812
rect 16632 11772 16638 11784
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 17644 11784 18276 11812
rect 17644 11772 17650 11784
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2096 11716 2605 11744
rect 2096 11704 2102 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 6696 11716 8217 11744
rect 6696 11704 6702 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8478 11744 8484 11756
rect 8439 11716 8484 11744
rect 8205 11707 8263 11713
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10836 11747 10894 11753
rect 10836 11744 10848 11747
rect 10468 11716 10848 11744
rect 10468 11704 10474 11716
rect 10836 11713 10848 11716
rect 10882 11744 10894 11747
rect 10962 11744 10968 11756
rect 10882 11716 10968 11744
rect 10882 11713 10894 11716
rect 10836 11707 10894 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11146 11744 11152 11756
rect 11103 11716 11152 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11146 11704 11152 11716
rect 11204 11744 11210 11756
rect 11882 11744 11888 11756
rect 11204 11716 11888 11744
rect 11204 11704 11210 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 17126 11744 17132 11756
rect 15611 11716 17132 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 2130 11676 2136 11688
rect 2091 11648 2136 11676
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 1489 11611 1547 11617
rect 1489 11577 1501 11611
rect 1535 11608 1547 11611
rect 1670 11608 1676 11620
rect 1535 11580 1676 11608
rect 1535 11577 1547 11580
rect 1489 11571 1547 11577
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 2240 11608 2268 11639
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2501 11679 2559 11685
rect 2501 11676 2513 11679
rect 2372 11648 2513 11676
rect 2372 11636 2378 11648
rect 2501 11645 2513 11648
rect 2547 11645 2559 11679
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 2501 11639 2559 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 6420 11648 6469 11676
rect 6420 11636 6426 11648
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 2406 11608 2412 11620
rect 2240 11580 2412 11608
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 4525 11611 4583 11617
rect 4525 11608 4537 11611
rect 3660 11580 4537 11608
rect 3660 11568 3666 11580
rect 4525 11577 4537 11580
rect 4571 11577 4583 11611
rect 4525 11571 4583 11577
rect 4890 11568 4896 11620
rect 4948 11608 4954 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4948 11580 5089 11608
rect 4948 11568 4954 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6840 11608 6868 11639
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7834 11676 7840 11688
rect 7064 11648 7840 11676
rect 7064 11636 7070 11648
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 12158 11676 12164 11688
rect 9907 11648 12164 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 6144 11580 6868 11608
rect 10689 11611 10747 11617
rect 6144 11568 6150 11580
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 10778 11608 10784 11620
rect 10735 11580 10784 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 12452 11552 12480 11639
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 12584 11648 13921 11676
rect 12584 11636 12590 11648
rect 13909 11645 13921 11648
rect 13955 11676 13967 11679
rect 13998 11676 14004 11688
rect 13955 11648 14004 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14458 11676 14464 11688
rect 14231 11648 14464 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16408 11608 16436 11639
rect 16574 11636 16580 11688
rect 16632 11676 16638 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16632 11648 16681 11676
rect 16632 11636 16638 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 17862 11676 17868 11688
rect 16669 11639 16727 11645
rect 16776 11648 17868 11676
rect 16776 11608 16804 11648
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 18248 11685 18276 11784
rect 18233 11679 18291 11685
rect 17972 11648 18184 11676
rect 16408 11580 16804 11608
rect 16850 11568 16856 11620
rect 16908 11568 16914 11620
rect 17129 11611 17187 11617
rect 17129 11577 17141 11611
rect 17175 11608 17187 11611
rect 17494 11608 17500 11620
rect 17175 11580 17500 11608
rect 17175 11577 17187 11580
rect 17129 11571 17187 11577
rect 17494 11568 17500 11580
rect 17552 11608 17558 11620
rect 17972 11608 18000 11648
rect 17552 11580 18000 11608
rect 18049 11611 18107 11617
rect 17552 11568 17558 11580
rect 18049 11577 18061 11611
rect 18095 11577 18107 11611
rect 18156 11608 18184 11648
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 18233 11639 18291 11645
rect 18340 11648 19625 11676
rect 18340 11608 18368 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 18156 11580 18368 11608
rect 18601 11611 18659 11617
rect 18049 11571 18107 11577
rect 18601 11577 18613 11611
rect 18647 11608 18659 11611
rect 18966 11608 18972 11620
rect 18647 11580 18972 11608
rect 18647 11577 18659 11580
rect 18601 11571 18659 11577
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6546 11540 6552 11552
rect 6319 11512 6552 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7926 11540 7932 11552
rect 7055 11512 7932 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 12434 11500 12440 11552
rect 12492 11500 12498 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12621 11543 12679 11549
rect 12621 11540 12633 11543
rect 12584 11512 12633 11540
rect 12584 11500 12590 11512
rect 12621 11509 12633 11512
rect 12667 11540 12679 11543
rect 13354 11540 13360 11552
rect 12667 11512 13360 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 16868 11540 16896 11568
rect 18064 11540 18092 11571
rect 18966 11568 18972 11580
rect 19024 11608 19030 11620
rect 19429 11611 19487 11617
rect 19429 11608 19441 11611
rect 19024 11580 19441 11608
rect 19024 11568 19030 11580
rect 19429 11577 19441 11580
rect 19475 11577 19487 11611
rect 19429 11571 19487 11577
rect 16540 11512 18092 11540
rect 16540 11500 16546 11512
rect 1104 11450 24840 11472
rect 1104 11398 8912 11450
rect 8964 11398 8976 11450
rect 9028 11398 9040 11450
rect 9092 11398 9104 11450
rect 9156 11398 16843 11450
rect 16895 11398 16907 11450
rect 16959 11398 16971 11450
rect 17023 11398 17035 11450
rect 17087 11398 24840 11450
rect 1104 11376 24840 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 6730 11336 6736 11348
rect 2832 11308 2877 11336
rect 6691 11308 6736 11336
rect 2832 11296 2838 11308
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 9769 11339 9827 11345
rect 9769 11336 9781 11339
rect 6880 11308 9781 11336
rect 6880 11296 6886 11308
rect 9769 11305 9781 11308
rect 9815 11305 9827 11339
rect 15562 11336 15568 11348
rect 9769 11299 9827 11305
rect 15396 11308 15568 11336
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 5500 11240 9720 11268
rect 5500 11228 5506 11240
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 4304 11172 4629 11200
rect 4304 11160 4310 11172
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 4890 11200 4896 11212
rect 4851 11172 4896 11200
rect 4617 11163 4675 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6972 11172 7297 11200
rect 6972 11160 6978 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8478 11200 8484 11212
rect 7883 11172 8484 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1578 11132 1584 11144
rect 1443 11104 1584 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1578 11092 1584 11104
rect 1636 11132 1642 11144
rect 1854 11132 1860 11144
rect 1636 11104 1860 11132
rect 1636 11092 1642 11104
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4154 11132 4160 11144
rect 4111 11104 4160 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 4856 11104 5089 11132
rect 4856 11092 4862 11104
rect 5077 11101 5089 11104
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7668 11132 7696 11163
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 9692 11209 9720 11240
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 11572 11172 13277 11200
rect 11572 11160 11578 11172
rect 12728 11144 12756 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 13449 11203 13507 11209
rect 13449 11200 13461 11203
rect 13412 11172 13461 11200
rect 13412 11160 13418 11172
rect 13449 11169 13461 11172
rect 13495 11169 13507 11203
rect 15396 11200 15424 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 17862 11296 17868 11348
rect 17920 11336 17926 11348
rect 19153 11339 19211 11345
rect 19153 11336 19165 11339
rect 17920 11308 19165 11336
rect 17920 11296 17926 11308
rect 19153 11305 19165 11308
rect 19199 11305 19211 11339
rect 19153 11299 19211 11305
rect 16945 11271 17003 11277
rect 16945 11237 16957 11271
rect 16991 11268 17003 11271
rect 17126 11268 17132 11280
rect 16991 11240 17132 11268
rect 16991 11237 17003 11240
rect 16945 11231 17003 11237
rect 17126 11228 17132 11240
rect 17184 11228 17190 11280
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15396 11172 15577 11200
rect 13449 11163 13507 11169
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 18046 11200 18052 11212
rect 18007 11172 18052 11200
rect 15565 11163 15623 11169
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 8110 11132 8116 11144
rect 7668 11104 8116 11132
rect 7377 11095 7435 11101
rect 7392 11064 7420 11095
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 9824 11104 10793 11132
rect 9824 11092 9830 11104
rect 10781 11101 10793 11104
rect 10827 11101 10839 11135
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 10781 11095 10839 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 12710 11092 12716 11144
rect 12768 11092 12774 11144
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 13688 11104 13737 11132
rect 13688 11092 13694 11104
rect 13725 11101 13737 11104
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14056 11104 15301 11132
rect 14056 11092 14062 11104
rect 15289 11101 15301 11104
rect 15335 11132 15347 11135
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 15335 11104 17785 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 7834 11064 7840 11076
rect 7392 11036 7840 11064
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 12158 11064 12164 11076
rect 12119 11036 12164 11064
rect 12158 11024 12164 11036
rect 12216 11064 12222 11076
rect 12434 11064 12440 11076
rect 12216 11036 12440 11064
rect 12216 11024 12222 11036
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 13464 11036 13676 11064
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 11238 10996 11244 11008
rect 6236 10968 11244 10996
rect 6236 10956 6242 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 11974 10956 11980 11008
rect 12032 10996 12038 11008
rect 13464 10996 13492 11036
rect 12032 10968 13492 10996
rect 13648 10996 13676 11036
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14734 11064 14740 11076
rect 14148 11036 14740 11064
rect 14148 11024 14154 11036
rect 14734 11024 14740 11036
rect 14792 11024 14798 11076
rect 16022 10996 16028 11008
rect 13648 10968 16028 10996
rect 12032 10956 12038 10968
rect 16022 10956 16028 10968
rect 16080 10956 16086 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 18414 10996 18420 11008
rect 16356 10968 18420 10996
rect 16356 10956 16362 10968
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 1104 10906 24840 10928
rect 1104 10854 4947 10906
rect 4999 10854 5011 10906
rect 5063 10854 5075 10906
rect 5127 10854 5139 10906
rect 5191 10854 12878 10906
rect 12930 10854 12942 10906
rect 12994 10854 13006 10906
rect 13058 10854 13070 10906
rect 13122 10854 20808 10906
rect 20860 10854 20872 10906
rect 20924 10854 20936 10906
rect 20988 10854 21000 10906
rect 21052 10854 24840 10906
rect 1104 10832 24840 10854
rect 3694 10752 3700 10804
rect 3752 10792 3758 10804
rect 5442 10792 5448 10804
rect 3752 10764 4844 10792
rect 5403 10764 5448 10792
rect 3752 10752 3758 10764
rect 4816 10724 4844 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6917 10795 6975 10801
rect 6917 10792 6929 10795
rect 5592 10764 6929 10792
rect 5592 10752 5598 10764
rect 6917 10761 6929 10764
rect 6963 10761 6975 10795
rect 6917 10755 6975 10761
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10792 10471 10795
rect 11054 10792 11060 10804
rect 10459 10764 11060 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 15473 10795 15531 10801
rect 11164 10764 15424 10792
rect 4816 10696 6868 10724
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 4154 10656 4160 10668
rect 1912 10628 3924 10656
rect 4115 10628 4160 10656
rect 1912 10616 1918 10628
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10588 2927 10591
rect 3142 10588 3148 10600
rect 2915 10560 3148 10588
rect 2915 10557 2927 10560
rect 2869 10551 2927 10557
rect 2608 10520 2636 10551
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 3896 10597 3924 10628
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 6546 10588 6552 10600
rect 3927 10560 6408 10588
rect 6507 10560 6552 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 3234 10520 3240 10532
rect 2608 10492 3240 10520
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 2590 10452 2596 10464
rect 2551 10424 2596 10452
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 6380 10461 6408 10560
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6840 10597 6868 10696
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 11164 10724 11192 10764
rect 7432 10696 11192 10724
rect 7432 10684 7438 10696
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 14369 10727 14427 10733
rect 11296 10696 14320 10724
rect 11296 10684 11302 10696
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10656 11115 10659
rect 11698 10656 11704 10668
rect 11103 10628 11704 10656
rect 11103 10625 11115 10628
rect 11057 10619 11115 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 11848 10628 13185 10656
rect 11848 10616 11854 10628
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 14292 10656 14320 10696
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 14458 10724 14464 10736
rect 14415 10696 14464 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 15396 10724 15424 10764
rect 15473 10761 15485 10795
rect 15519 10792 15531 10795
rect 15562 10792 15568 10804
rect 15519 10764 15568 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 16666 10792 16672 10804
rect 16448 10764 16672 10792
rect 16448 10752 16454 10764
rect 16666 10752 16672 10764
rect 16724 10792 16730 10804
rect 17586 10792 17592 10804
rect 16724 10764 17592 10792
rect 16724 10752 16730 10764
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 15396 10696 20208 10724
rect 14292 10628 19380 10656
rect 13173 10619 13231 10625
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6840 10520 6868 10551
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7708 10560 7849 10588
rect 7708 10548 7714 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 8018 10588 8024 10600
rect 7979 10560 8024 10588
rect 7837 10551 7895 10557
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 10778 10588 10784 10600
rect 8803 10560 10784 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 7926 10520 7932 10532
rect 6840 10492 7932 10520
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 8036 10520 8064 10548
rect 8588 10520 8616 10551
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10557 11391 10591
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11333 10551 11391 10557
rect 8036 10492 8616 10520
rect 6365 10455 6423 10461
rect 6365 10421 6377 10455
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7374 10452 7380 10464
rect 7064 10424 7380 10452
rect 7064 10412 7070 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9033 10455 9091 10461
rect 9033 10421 9045 10455
rect 9079 10452 9091 10455
rect 9950 10452 9956 10464
rect 9079 10424 9956 10452
rect 9079 10421 9091 10424
rect 9033 10415 9091 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10980 10452 11008 10551
rect 11348 10520 11376 10551
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 12526 10588 12532 10600
rect 11624 10560 12532 10588
rect 11624 10520 11652 10560
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 13262 10548 13268 10600
rect 13320 10588 13326 10600
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 13320 10560 13369 10588
rect 13320 10548 13326 10560
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13357 10551 13415 10557
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 15286 10588 15292 10600
rect 14139 10560 15292 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 16022 10588 16028 10600
rect 15983 10560 16028 10588
rect 16022 10548 16028 10560
rect 16080 10548 16086 10600
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16390 10588 16396 10600
rect 16172 10560 16217 10588
rect 16351 10560 16396 10588
rect 16172 10548 16178 10560
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 18049 10591 18107 10597
rect 16540 10560 16585 10588
rect 16540 10548 16546 10560
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18230 10588 18236 10600
rect 18095 10560 18236 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 19153 10591 19211 10597
rect 19153 10588 19165 10591
rect 18472 10560 19165 10588
rect 18472 10548 18478 10560
rect 19153 10557 19165 10560
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 11348 10492 11652 10520
rect 11992 10492 19257 10520
rect 11992 10452 12020 10492
rect 19245 10489 19257 10492
rect 19291 10489 19303 10523
rect 19352 10520 19380 10628
rect 20180 10597 20208 10696
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 20257 10523 20315 10529
rect 20257 10520 20269 10523
rect 19352 10492 20269 10520
rect 19245 10483 19303 10489
rect 20257 10489 20269 10492
rect 20303 10489 20315 10523
rect 20257 10483 20315 10489
rect 10980 10424 12020 10452
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13906 10452 13912 10464
rect 13780 10424 13912 10452
rect 13780 10412 13786 10424
rect 13906 10412 13912 10424
rect 13964 10452 13970 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 13964 10424 18245 10452
rect 13964 10412 13970 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18233 10415 18291 10421
rect 1104 10362 24840 10384
rect 1104 10310 8912 10362
rect 8964 10310 8976 10362
rect 9028 10310 9040 10362
rect 9092 10310 9104 10362
rect 9156 10310 16843 10362
rect 16895 10310 16907 10362
rect 16959 10310 16971 10362
rect 17023 10310 17035 10362
rect 17087 10310 24840 10362
rect 1104 10288 24840 10310
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 11330 10248 11336 10260
rect 2464 10220 4016 10248
rect 2464 10208 2470 10220
rect 2590 10112 2596 10124
rect 2551 10084 2596 10112
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3142 10112 3148 10124
rect 3103 10084 3148 10112
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 3694 10044 3700 10056
rect 2731 10016 3700 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 2038 9976 2044 9988
rect 1999 9948 2044 9976
rect 2038 9936 2044 9948
rect 2096 9936 2102 9988
rect 3988 9976 4016 10220
rect 4080 10220 11336 10248
rect 4080 10121 4108 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13906 10248 13912 10260
rect 13688 10220 13912 10248
rect 13688 10208 13694 10220
rect 13906 10208 13912 10220
rect 13964 10248 13970 10260
rect 13964 10220 15516 10248
rect 13964 10208 13970 10220
rect 7006 10180 7012 10192
rect 6967 10152 7012 10180
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7466 10180 7472 10192
rect 7156 10152 7472 10180
rect 7156 10140 7162 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 15488 10180 15516 10220
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 16080 10220 19165 10248
rect 16080 10208 16086 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 16298 10180 16304 10192
rect 15488 10152 16304 10180
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 16482 10180 16488 10192
rect 16443 10152 16488 10180
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 17221 10183 17279 10189
rect 17221 10149 17233 10183
rect 17267 10180 17279 10183
rect 17954 10180 17960 10192
rect 17267 10152 17960 10180
rect 17267 10149 17279 10152
rect 17221 10143 17279 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 6638 10112 6644 10124
rect 5399 10084 6644 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7024 10084 7849 10112
rect 7024 10056 7052 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 7837 10075 7895 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9950 10112 9956 10124
rect 9911 10084 9956 10112
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 12250 10112 12256 10124
rect 11112 10084 12256 10112
rect 11112 10072 11118 10084
rect 12250 10072 12256 10084
rect 12308 10112 12314 10124
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12308 10084 12725 10112
rect 12308 10072 12314 10084
rect 12713 10081 12725 10084
rect 12759 10081 12771 10115
rect 12713 10075 12771 10081
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10112 13231 10115
rect 13722 10112 13728 10124
rect 13219 10084 13728 10112
rect 13219 10081 13231 10084
rect 13173 10075 13231 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 13955 10084 15148 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 11974 10044 11980 10056
rect 7984 10016 11980 10044
rect 7984 10004 7990 10016
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12492 10016 13001 10044
rect 12492 10004 12498 10016
rect 12989 10013 13001 10016
rect 13035 10013 13047 10047
rect 15120 10044 15148 10084
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 16666 10121 16672 10124
rect 15295 10115 15353 10121
rect 15295 10112 15307 10115
rect 15252 10084 15307 10112
rect 15252 10072 15258 10084
rect 15295 10081 15307 10084
rect 15341 10081 15353 10115
rect 15295 10075 15353 10081
rect 16632 10115 16672 10121
rect 16632 10081 16644 10115
rect 16632 10075 16672 10081
rect 16666 10072 16672 10075
rect 16724 10072 16730 10124
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 16776 10084 18061 10112
rect 16206 10044 16212 10056
rect 15120 10016 16212 10044
rect 12989 10007 13047 10013
rect 16206 10004 16212 10016
rect 16264 10044 16270 10056
rect 16390 10044 16396 10056
rect 16264 10016 16396 10044
rect 16264 10004 16270 10016
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 16776 10044 16804 10084
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 18966 10072 18972 10124
rect 19024 10112 19030 10124
rect 19061 10115 19119 10121
rect 19061 10112 19073 10115
rect 19024 10084 19073 10112
rect 19024 10072 19030 10084
rect 19061 10081 19073 10084
rect 19107 10081 19119 10115
rect 20898 10112 20904 10124
rect 20859 10084 20904 10112
rect 19061 10075 19119 10081
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 16540 10016 16804 10044
rect 16853 10047 16911 10053
rect 16540 10004 16546 10016
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 17218 10044 17224 10056
rect 16899 10016 17224 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 4249 9979 4307 9985
rect 4249 9976 4261 9979
rect 3988 9948 4261 9976
rect 4249 9945 4261 9948
rect 4295 9945 4307 9979
rect 4249 9939 4307 9945
rect 7484 9948 9720 9976
rect 4264 9908 4292 9939
rect 7484 9908 7512 9948
rect 4264 9880 7512 9908
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 8018 9908 8024 9920
rect 7616 9880 8024 9908
rect 7616 9868 7622 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 9692 9908 9720 9948
rect 13262 9936 13268 9988
rect 13320 9976 13326 9988
rect 16761 9979 16819 9985
rect 13320 9948 15516 9976
rect 13320 9936 13326 9948
rect 10134 9908 10140 9920
rect 9692 9880 10140 9908
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 11241 9911 11299 9917
rect 11241 9877 11253 9911
rect 11287 9908 11299 9911
rect 11514 9908 11520 9920
rect 11287 9880 11520 9908
rect 11287 9877 11299 9880
rect 11241 9871 11299 9877
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12400 9880 12541 9908
rect 12400 9868 12406 9880
rect 12529 9877 12541 9880
rect 12575 9908 12587 9911
rect 13998 9908 14004 9920
rect 12575 9880 14004 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 13998 9868 14004 9880
rect 14056 9868 14062 9920
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15488 9917 15516 9948
rect 16761 9945 16773 9979
rect 16807 9976 16819 9979
rect 17310 9976 17316 9988
rect 16807 9948 17316 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 18230 9976 18236 9988
rect 17420 9948 18236 9976
rect 15473 9911 15531 9917
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 17420 9908 17448 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 18138 9908 18144 9920
rect 15519 9880 17448 9908
rect 18099 9880 18144 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 20993 9911 21051 9917
rect 20993 9877 21005 9911
rect 21039 9908 21051 9911
rect 21174 9908 21180 9920
rect 21039 9880 21180 9908
rect 21039 9877 21051 9880
rect 20993 9871 21051 9877
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 1104 9818 24840 9840
rect 1104 9766 4947 9818
rect 4999 9766 5011 9818
rect 5063 9766 5075 9818
rect 5127 9766 5139 9818
rect 5191 9766 12878 9818
rect 12930 9766 12942 9818
rect 12994 9766 13006 9818
rect 13058 9766 13070 9818
rect 13122 9766 20808 9818
rect 20860 9766 20872 9818
rect 20924 9766 20936 9818
rect 20988 9766 21000 9818
rect 21052 9766 24840 9818
rect 1104 9744 24840 9766
rect 4540 9676 5488 9704
rect 3050 9596 3056 9648
rect 3108 9636 3114 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 3108 9608 3433 9636
rect 3108 9596 3114 9608
rect 3421 9605 3433 9608
rect 3467 9636 3479 9639
rect 4540 9636 4568 9676
rect 5166 9636 5172 9648
rect 3467 9608 4568 9636
rect 4632 9608 5172 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 4632 9577 4660 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5460 9636 5488 9676
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 5776 9676 5821 9704
rect 9692 9676 10640 9704
rect 5776 9664 5782 9676
rect 9692 9636 9720 9676
rect 5460 9608 9720 9636
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6270 9568 6276 9580
rect 5868 9540 6276 9568
rect 5868 9528 5874 9540
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 8803 9540 9965 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 10612 9568 10640 9676
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 18138 9704 18144 9716
rect 10836 9676 18144 9704
rect 10836 9664 10842 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 11020 9608 16160 9636
rect 11020 9596 11026 9608
rect 10612 9540 11376 9568
rect 9953 9531 10011 9537
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1964 9472 2145 9500
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 1964 9432 1992 9472
rect 2133 9469 2145 9472
rect 2179 9500 2191 9503
rect 4709 9503 4767 9509
rect 2179 9472 4660 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 1811 9404 1992 9432
rect 4632 9432 4660 9472
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4890 9500 4896 9512
rect 4755 9472 4896 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5132 9472 5273 9500
rect 5132 9460 5138 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9500 5503 9503
rect 6178 9500 6184 9512
rect 5491 9472 6184 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 7558 9460 7564 9512
rect 7616 9509 7622 9512
rect 7616 9503 7665 9509
rect 7616 9469 7619 9503
rect 7653 9469 7665 9503
rect 7742 9500 7748 9512
rect 7703 9472 7748 9500
rect 7616 9463 7665 9469
rect 7616 9460 7622 9463
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8570 9500 8576 9512
rect 8251 9472 8576 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 7466 9432 7472 9444
rect 4632 9404 7472 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 8128 9432 8156 9463
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9674 9500 9680 9512
rect 9635 9472 9680 9500
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10410 9500 10416 9512
rect 9784 9472 10416 9500
rect 9784 9432 9812 9472
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 8128 9404 9812 9432
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3878 9364 3884 9376
rect 3476 9336 3884 9364
rect 3476 9324 3482 9336
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 7834 9364 7840 9376
rect 5500 9336 7840 9364
rect 5500 9324 5506 9336
rect 7834 9324 7840 9336
rect 7892 9364 7898 9376
rect 10962 9364 10968 9376
rect 7892 9336 10968 9364
rect 7892 9324 7898 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11238 9364 11244 9376
rect 11199 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11348 9364 11376 9540
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 11940 9540 12541 9568
rect 11940 9528 11946 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13722 9568 13728 9580
rect 13587 9540 13728 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 11974 9460 11980 9512
rect 12032 9500 12038 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12032 9472 12449 9500
rect 12032 9460 12038 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13688 9472 14197 9500
rect 13688 9460 13694 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 16132 9500 16160 9608
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 16356 9540 20116 9568
rect 16356 9528 16362 9540
rect 16197 9503 16255 9509
rect 16197 9500 16209 9503
rect 16132 9472 16209 9500
rect 14369 9463 14427 9469
rect 16197 9469 16209 9472
rect 16243 9469 16255 9503
rect 16197 9463 16255 9469
rect 14384 9432 14412 9463
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17276 9472 18061 9500
rect 17276 9460 17282 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 20088 9509 20116 9540
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 18196 9472 19073 9500
rect 18196 9460 18202 9472
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 15470 9432 15476 9444
rect 14384 9404 15476 9432
rect 15470 9392 15476 9404
rect 15528 9432 15534 9444
rect 15528 9404 18184 9432
rect 15528 9392 15534 9404
rect 16298 9364 16304 9376
rect 11348 9336 16304 9364
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16574 9364 16580 9376
rect 16439 9336 16580 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 18156 9373 18184 9404
rect 18230 9392 18236 9444
rect 18288 9432 18294 9444
rect 19153 9435 19211 9441
rect 19153 9432 19165 9435
rect 18288 9404 19165 9432
rect 18288 9392 18294 9404
rect 19153 9401 19165 9404
rect 19199 9401 19211 9435
rect 19153 9395 19211 9401
rect 18141 9367 18199 9373
rect 18141 9333 18153 9367
rect 18187 9333 18199 9367
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 18141 9327 18199 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 1104 9274 24840 9296
rect 1104 9222 8912 9274
rect 8964 9222 8976 9274
rect 9028 9222 9040 9274
rect 9092 9222 9104 9274
rect 9156 9222 16843 9274
rect 16895 9222 16907 9274
rect 16959 9222 16971 9274
rect 17023 9222 17035 9274
rect 17087 9222 24840 9274
rect 1104 9200 24840 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 2130 9160 2136 9172
rect 1535 9132 2136 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 2700 9132 19625 9160
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2700 9033 2728 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 19613 9123 19671 9129
rect 3142 9092 3148 9104
rect 3103 9064 3148 9092
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 5350 9092 5356 9104
rect 3936 9064 5356 9092
rect 3936 9052 3942 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 5629 9095 5687 9101
rect 5629 9061 5641 9095
rect 5675 9061 5687 9095
rect 5629 9055 5687 9061
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 2424 8956 2452 8987
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4212 8996 4537 9024
rect 4212 8984 4218 8996
rect 4525 8993 4537 8996
rect 4571 9024 4583 9027
rect 5074 9024 5080 9036
rect 4571 8996 5080 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 9024 5319 9027
rect 5442 9024 5448 9036
rect 5307 8996 5448 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5644 9024 5672 9055
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 8205 9095 8263 9101
rect 8205 9092 8217 9095
rect 8168 9064 8217 9092
rect 8168 9052 8174 9064
rect 8205 9061 8217 9064
rect 8251 9092 8263 9095
rect 8294 9092 8300 9104
rect 8251 9064 8300 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 9214 9052 9220 9104
rect 9272 9092 9278 9104
rect 9769 9095 9827 9101
rect 9769 9092 9781 9095
rect 9272 9064 9781 9092
rect 9272 9052 9278 9064
rect 9769 9061 9781 9064
rect 9815 9061 9827 9095
rect 9769 9055 9827 9061
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 14277 9095 14335 9101
rect 12492 9064 14044 9092
rect 12492 9052 12498 9064
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 5644 8996 6837 9024
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 8018 9024 8024 9036
rect 6972 8996 8024 9024
rect 6972 8984 6978 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 9685 9027 9743 9033
rect 9685 8993 9697 9027
rect 9731 8993 9743 9027
rect 9685 8987 9743 8993
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11054 9024 11060 9036
rect 10919 8996 11060 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 2866 8956 2872 8968
rect 2424 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6730 8956 6736 8968
rect 6595 8928 6736 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 4062 8888 4068 8900
rect 2547 8860 4068 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 4448 8888 4476 8919
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 9692 8956 9720 8987
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11241 9027 11299 9033
rect 11241 8993 11253 9027
rect 11287 9024 11299 9027
rect 12342 9024 12348 9036
rect 11287 8996 12348 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12894 9024 12900 9036
rect 12855 8996 12900 9024
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 13814 9024 13820 9036
rect 13771 8996 13820 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 14016 9024 14044 9064
rect 14277 9061 14289 9095
rect 14323 9092 14335 9095
rect 14550 9092 14556 9104
rect 14323 9064 14556 9092
rect 14323 9061 14335 9064
rect 14277 9055 14335 9061
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 17368 9064 18552 9092
rect 17368 9052 17374 9064
rect 18138 9024 18144 9036
rect 14016 8996 18144 9024
rect 13909 8987 13967 8993
rect 11146 8956 11152 8968
rect 9692 8928 11152 8956
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11514 8956 11520 8968
rect 11475 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13924 8956 13952 8987
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18524 9033 18552 9064
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 8993 18567 9027
rect 18509 8987 18567 8993
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 12584 8928 13952 8956
rect 12584 8916 12590 8928
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 16025 8959 16083 8965
rect 16025 8956 16037 8959
rect 14056 8928 16037 8956
rect 14056 8916 14062 8928
rect 16025 8925 16037 8928
rect 16071 8925 16083 8959
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16025 8919 16083 8925
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17276 8928 17417 8956
rect 17276 8916 17282 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 6454 8888 6460 8900
rect 4448 8860 6460 8888
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 10778 8888 10784 8900
rect 9600 8860 10784 8888
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 9600 8820 9628 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 19536 8888 19564 8987
rect 17552 8860 19564 8888
rect 17552 8848 17558 8860
rect 3016 8792 9628 8820
rect 3016 8780 3022 8792
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 9732 8792 10701 8820
rect 9732 8780 9738 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13262 8820 13268 8832
rect 12492 8792 13268 8820
rect 12492 8780 12498 8792
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 18601 8823 18659 8829
rect 18601 8820 18613 8823
rect 16448 8792 18613 8820
rect 16448 8780 16454 8792
rect 18601 8789 18613 8792
rect 18647 8789 18659 8823
rect 18601 8783 18659 8789
rect 1104 8730 24840 8752
rect 1104 8678 4947 8730
rect 4999 8678 5011 8730
rect 5063 8678 5075 8730
rect 5127 8678 5139 8730
rect 5191 8678 12878 8730
rect 12930 8678 12942 8730
rect 12994 8678 13006 8730
rect 13058 8678 13070 8730
rect 13122 8678 20808 8730
rect 20860 8678 20872 8730
rect 20924 8678 20936 8730
rect 20988 8678 21000 8730
rect 21052 8678 24840 8730
rect 1104 8656 24840 8678
rect 4338 8616 4344 8628
rect 4299 8588 4344 8616
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7524 8588 12848 8616
rect 7524 8576 7530 8588
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 2682 8548 2688 8560
rect 2372 8520 2688 8548
rect 2372 8508 2378 8520
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 5350 8548 5356 8560
rect 3804 8520 5356 8548
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 2682 8412 2688 8424
rect 2547 8384 2688 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 2958 8412 2964 8424
rect 2919 8384 2964 8412
rect 2777 8375 2835 8381
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 1949 8347 2007 8353
rect 1949 8344 1961 8347
rect 1728 8316 1961 8344
rect 1728 8304 1734 8316
rect 1949 8313 1961 8316
rect 1995 8313 2007 8347
rect 2792 8344 2820 8375
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3804 8412 3832 8520
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 5629 8551 5687 8557
rect 5629 8548 5641 8551
rect 5408 8520 5641 8548
rect 5408 8508 5414 8520
rect 5629 8517 5641 8520
rect 5675 8517 5687 8551
rect 5629 8511 5687 8517
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 7190 8548 7196 8560
rect 6972 8520 7196 8548
rect 6972 8508 6978 8520
rect 7190 8508 7196 8520
rect 7248 8548 7254 8560
rect 10962 8548 10968 8560
rect 7248 8520 10732 8548
rect 10923 8520 10968 8548
rect 7248 8508 7254 8520
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 4430 8480 4436 8492
rect 3927 8452 4436 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3804 8384 4077 8412
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4246 8412 4252 8424
rect 4203 8384 4252 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5534 8412 5540 8424
rect 5491 8384 5540 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6420 8384 6837 8412
rect 6420 8372 6426 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 8386 8412 8392 8424
rect 8347 8384 8392 8412
rect 6825 8375 6883 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 10704 8421 10732 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 11330 8480 11336 8492
rect 11103 8452 11336 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11330 8440 11336 8452
rect 11388 8480 11394 8492
rect 11974 8480 11980 8492
rect 11388 8452 11980 8480
rect 11388 8440 11394 8452
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 10689 8415 10747 8421
rect 9355 8384 10640 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 4522 8344 4528 8356
rect 2792 8316 4528 8344
rect 1949 8307 2007 8313
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 8588 8344 8616 8372
rect 9140 8344 9168 8375
rect 9766 8344 9772 8356
rect 8588 8316 9772 8344
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 10612 8344 10640 8384
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10836 8415 10894 8421
rect 10836 8381 10848 8415
rect 10882 8412 10894 8415
rect 11238 8412 11244 8424
rect 10882 8384 11244 8412
rect 10882 8381 10894 8384
rect 10836 8375 10894 8381
rect 11238 8372 11244 8384
rect 11296 8412 11302 8424
rect 12342 8412 12348 8424
rect 11296 8384 12348 8412
rect 11296 8372 11302 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12710 8344 12716 8356
rect 10612 8316 11468 8344
rect 12671 8316 12716 8344
rect 10888 8288 10916 8316
rect 382 8236 388 8288
rect 440 8276 446 8288
rect 6086 8276 6092 8288
rect 440 8248 6092 8276
rect 440 8236 446 8248
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 7006 8276 7012 8288
rect 6967 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 9582 8276 9588 8288
rect 9543 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10870 8236 10876 8288
rect 10928 8236 10934 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11333 8279 11391 8285
rect 11333 8276 11345 8279
rect 11112 8248 11345 8276
rect 11112 8236 11118 8248
rect 11333 8245 11345 8248
rect 11379 8245 11391 8279
rect 11440 8276 11468 8316
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 12820 8344 12848 8588
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 13320 8588 16957 8616
rect 13320 8576 13326 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 19150 8616 19156 8628
rect 19111 8588 19156 8616
rect 16945 8579 17003 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 12878 8551 12936 8557
rect 12878 8517 12890 8551
rect 12924 8517 12936 8551
rect 12878 8511 12936 8517
rect 12989 8551 13047 8557
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 13814 8548 13820 8560
rect 13035 8520 13820 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 12893 8480 12921 8511
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 15933 8551 15991 8557
rect 14056 8520 14320 8548
rect 14056 8508 14062 8520
rect 13262 8480 13268 8492
rect 12893 8452 13268 8480
rect 13262 8440 13268 8452
rect 13320 8480 13326 8492
rect 13722 8480 13728 8492
rect 13320 8452 13728 8480
rect 13320 8440 13326 8452
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14292 8424 14320 8520
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 17218 8548 17224 8560
rect 15979 8520 17224 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 20162 8480 20168 8492
rect 14792 8452 20168 8480
rect 14792 8440 14798 8452
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 13052 8415 13110 8421
rect 13052 8381 13064 8415
rect 13098 8412 13110 8415
rect 13354 8412 13360 8424
rect 13098 8384 13360 8412
rect 13098 8381 13110 8384
rect 13052 8375 13110 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13998 8412 14004 8424
rect 13495 8384 14004 8412
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14332 8384 14381 8412
rect 14332 8372 14338 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 14976 8384 16865 8412
rect 14976 8372 14982 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 18012 8384 18061 8412
rect 18012 8372 18018 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 19058 8412 19064 8424
rect 19019 8384 19064 8412
rect 18049 8375 18107 8381
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 21174 8344 21180 8356
rect 12820 8316 13400 8344
rect 13262 8276 13268 8288
rect 11440 8248 13268 8276
rect 11333 8239 11391 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 13372 8276 13400 8316
rect 15304 8316 21180 8344
rect 15304 8276 15332 8316
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 18138 8276 18144 8288
rect 13372 8248 15332 8276
rect 18099 8248 18144 8276
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 1104 8186 24840 8208
rect 1104 8134 8912 8186
rect 8964 8134 8976 8186
rect 9028 8134 9040 8186
rect 9092 8134 9104 8186
rect 9156 8134 16843 8186
rect 16895 8134 16907 8186
rect 16959 8134 16971 8186
rect 17023 8134 17035 8186
rect 17087 8134 24840 8186
rect 1104 8112 24840 8134
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4028 8044 4261 8072
rect 4028 8032 4034 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 7374 8072 7380 8084
rect 4249 8035 4307 8041
rect 6104 8044 7380 8072
rect 6104 8013 6132 8044
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 10962 8072 10968 8084
rect 9784 8044 10968 8072
rect 6089 8007 6147 8013
rect 6089 7973 6101 8007
rect 6135 7973 6147 8007
rect 6914 8004 6920 8016
rect 6089 7967 6147 7973
rect 6472 7976 6920 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4338 7936 4344 7948
rect 4111 7908 4344 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5537 7939 5595 7945
rect 5537 7936 5549 7939
rect 5316 7908 5549 7936
rect 5316 7896 5322 7908
rect 5537 7905 5549 7908
rect 5583 7905 5595 7939
rect 5537 7899 5595 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6472 7936 6500 7976
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 9784 8004 9812 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 12250 8072 12256 8084
rect 11296 8044 12256 8072
rect 11296 8032 11302 8044
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12710 8072 12716 8084
rect 12492 8044 12716 8072
rect 12492 8032 12498 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 15381 8075 15439 8081
rect 15381 8072 15393 8075
rect 13320 8044 15393 8072
rect 13320 8032 13326 8044
rect 15381 8041 15393 8044
rect 15427 8041 15439 8075
rect 15381 8035 15439 8041
rect 7300 7976 9812 8004
rect 5675 7908 6500 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6604 7908 7113 7936
rect 6604 7896 6610 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7868 1458 7880
rect 1854 7868 1860 7880
rect 1452 7840 1860 7868
rect 1452 7828 1458 7840
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 5350 7868 5356 7880
rect 5311 7840 5356 7868
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4120 7772 7052 7800
rect 4120 7760 4126 7772
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6788 7704 6929 7732
rect 6788 7692 6794 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 7024 7732 7052 7772
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7300 7800 7328 7976
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 12161 8007 12219 8013
rect 12161 8004 12173 8007
rect 11572 7976 12173 8004
rect 11572 7964 11578 7976
rect 12161 7973 12173 7976
rect 12207 7973 12219 8007
rect 13630 8004 13636 8016
rect 12161 7967 12219 7973
rect 12728 7976 13636 8004
rect 12728 7948 12756 7976
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 14550 8004 14556 8016
rect 14108 7976 14556 8004
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 7558 7936 7564 7948
rect 7423 7908 7564 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 7558 7896 7564 7908
rect 7616 7936 7622 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7616 7908 7941 7936
rect 7616 7896 7622 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 9214 7936 9220 7948
rect 8159 7908 9220 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9953 7939 10011 7945
rect 9953 7936 9965 7939
rect 9640 7908 9965 7936
rect 9640 7896 9646 7908
rect 9953 7905 9965 7908
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 12710 7896 12716 7948
rect 12768 7896 12774 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 12860 7908 12905 7936
rect 12860 7896 12866 7908
rect 13078 7896 13084 7948
rect 13136 7936 13142 7948
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 13136 7908 13185 7936
rect 13136 7896 13142 7908
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13265 7871 13323 7877
rect 12952 7840 12997 7868
rect 12952 7828 12958 7840
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 14108 7868 14136 7976
rect 14550 7964 14556 7976
rect 14608 7964 14614 8016
rect 16298 8004 16304 8016
rect 16259 7976 16304 8004
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 18138 8004 18144 8016
rect 16960 7976 18144 8004
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7936 14335 7939
rect 14366 7936 14372 7948
rect 14323 7908 14372 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 13311 7840 14136 7868
rect 14200 7868 14228 7899
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 16960 7945 16988 7976
rect 18138 7964 18144 7976
rect 18196 7964 18202 8016
rect 16945 7939 17003 7945
rect 16945 7905 16957 7939
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 17276 7908 17325 7936
rect 17276 7896 17282 7908
rect 17313 7905 17325 7908
rect 17359 7905 17371 7939
rect 17494 7936 17500 7948
rect 17455 7908 17500 7936
rect 17313 7899 17371 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 14458 7868 14464 7880
rect 14200 7840 14464 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16632 7840 17049 7868
rect 16632 7828 16638 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 8294 7800 8300 7812
rect 7156 7772 7328 7800
rect 8255 7772 8300 7800
rect 7156 7760 7162 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 11698 7800 11704 7812
rect 10612 7772 11704 7800
rect 10612 7732 10640 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 12342 7800 12348 7812
rect 12032 7772 12348 7800
rect 12032 7760 12038 7772
rect 12342 7760 12348 7772
rect 12400 7800 12406 7812
rect 12400 7772 12480 7800
rect 12400 7760 12406 7772
rect 7024 7704 10640 7732
rect 12452 7732 12480 7772
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 16850 7800 16856 7812
rect 12860 7772 16856 7800
rect 12860 7760 12866 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 14918 7732 14924 7744
rect 12452 7704 14924 7732
rect 6917 7695 6975 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 1104 7642 24840 7664
rect 1104 7590 4947 7642
rect 4999 7590 5011 7642
rect 5063 7590 5075 7642
rect 5127 7590 5139 7642
rect 5191 7590 12878 7642
rect 12930 7590 12942 7642
rect 12994 7590 13006 7642
rect 13058 7590 13070 7642
rect 13122 7590 20808 7642
rect 20860 7590 20872 7642
rect 20924 7590 20936 7642
rect 20988 7590 21000 7642
rect 21052 7590 24840 7642
rect 1104 7568 24840 7590
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 3970 7528 3976 7540
rect 3844 7500 3976 7528
rect 3844 7488 3850 7500
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 4580 7500 7021 7528
rect 4580 7488 4586 7500
rect 7009 7497 7021 7500
rect 7055 7528 7067 7531
rect 9490 7528 9496 7540
rect 7055 7500 9496 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10686 7528 10692 7540
rect 10100 7500 10692 7528
rect 10100 7488 10106 7500
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 18414 7528 18420 7540
rect 11756 7500 18420 7528
rect 11756 7488 11762 7500
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10502 7460 10508 7472
rect 9732 7432 10508 7460
rect 9732 7420 9738 7432
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11103 7432 12480 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 5442 7392 5448 7404
rect 2240 7364 3832 7392
rect 2240 7333 2268 7364
rect 2231 7327 2289 7333
rect 2231 7293 2243 7327
rect 2277 7293 2289 7327
rect 2231 7287 2289 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3694 7324 3700 7336
rect 3651 7296 3700 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 2406 7188 2412 7200
rect 2367 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2682 7148 2688 7200
rect 2740 7188 2746 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 2740 7160 3433 7188
rect 2740 7148 2746 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3804 7188 3832 7364
rect 3896 7364 5448 7392
rect 3896 7333 3924 7364
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 6788 7364 8033 7392
rect 6788 7352 6794 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8294 7392 8300 7404
rect 8255 7364 8300 7392
rect 8021 7355 8079 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 10928 7395 10986 7401
rect 10928 7361 10940 7395
rect 10974 7392 10986 7395
rect 11606 7392 11612 7404
rect 10974 7364 11612 7392
rect 10974 7361 10986 7364
rect 10928 7355 10986 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 12452 7392 12480 7432
rect 12526 7420 12532 7472
rect 12584 7469 12590 7472
rect 12584 7463 12633 7469
rect 12584 7429 12587 7463
rect 12621 7429 12633 7463
rect 12584 7423 12633 7429
rect 12713 7463 12771 7469
rect 12713 7429 12725 7463
rect 12759 7460 12771 7463
rect 13722 7460 13728 7472
rect 12759 7432 13728 7460
rect 12759 7429 12771 7432
rect 12713 7423 12771 7429
rect 12584 7420 12590 7423
rect 12728 7392 12756 7423
rect 13722 7420 13728 7432
rect 13780 7420 13786 7472
rect 16850 7460 16856 7472
rect 16811 7432 16856 7460
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 12452 7364 12756 7392
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 13170 7392 13176 7404
rect 12860 7364 13176 7392
rect 12860 7352 12866 7364
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14240 7364 14565 7392
rect 14240 7352 14246 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 19058 7392 19064 7404
rect 14553 7355 14611 7361
rect 15764 7364 19064 7392
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4580 7296 4905 7324
rect 4580 7284 4586 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 5258 7324 5264 7336
rect 5215 7296 5264 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 5675 7296 6837 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 11120 7327 11178 7333
rect 11120 7293 11132 7327
rect 11166 7324 11178 7327
rect 11517 7327 11575 7333
rect 11166 7296 11468 7324
rect 11166 7293 11178 7296
rect 11120 7287 11178 7293
rect 5074 7256 5080 7268
rect 5035 7228 5080 7256
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 10781 7259 10839 7265
rect 10781 7225 10793 7259
rect 10827 7256 10839 7259
rect 10962 7256 10968 7268
rect 10827 7228 10968 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 6914 7188 6920 7200
rect 3804 7160 6920 7188
rect 3421 7151 3479 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7188 9643 7191
rect 11054 7188 11060 7200
rect 9631 7160 11060 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11440 7188 11468 7296
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 14274 7324 14280 7336
rect 11563 7296 12756 7324
rect 14235 7296 14280 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 12434 7216 12440 7268
rect 12492 7256 12498 7268
rect 12728 7256 12756 7296
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 15764 7324 15792 7364
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 14384 7296 15792 7324
rect 16761 7327 16819 7333
rect 14384 7256 14412 7296
rect 16761 7293 16773 7327
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 16776 7256 16804 7287
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17552 7296 18061 7324
rect 17552 7284 17558 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 17310 7256 17316 7268
rect 12492 7228 12537 7256
rect 12728 7228 14412 7256
rect 15212 7228 16804 7256
rect 16868 7228 17316 7256
rect 12492 7216 12498 7228
rect 12802 7188 12808 7200
rect 11440 7160 12808 7188
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13081 7191 13139 7197
rect 13081 7157 13093 7191
rect 13127 7188 13139 7191
rect 13722 7188 13728 7200
rect 13127 7160 13728 7188
rect 13127 7157 13139 7160
rect 13081 7151 13139 7157
rect 13722 7148 13728 7160
rect 13780 7188 13786 7200
rect 15212 7188 15240 7228
rect 13780 7160 15240 7188
rect 15841 7191 15899 7197
rect 13780 7148 13786 7160
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16574 7188 16580 7200
rect 15887 7160 16580 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 16574 7148 16580 7160
rect 16632 7188 16638 7200
rect 16868 7188 16896 7228
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 16632 7160 16896 7188
rect 16632 7148 16638 7160
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 18141 7191 18199 7197
rect 18141 7188 18153 7191
rect 17184 7160 18153 7188
rect 17184 7148 17190 7160
rect 18141 7157 18153 7160
rect 18187 7157 18199 7191
rect 18141 7151 18199 7157
rect 1104 7098 24840 7120
rect 1104 7046 8912 7098
rect 8964 7046 8976 7098
rect 9028 7046 9040 7098
rect 9092 7046 9104 7098
rect 9156 7046 16843 7098
rect 16895 7046 16907 7098
rect 16959 7046 16971 7098
rect 17023 7046 17035 7098
rect 17087 7046 24840 7098
rect 1104 7024 24840 7046
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 12158 6984 12164 6996
rect 4304 6956 4568 6984
rect 4304 6944 4310 6956
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 4154 6916 4160 6928
rect 3752 6888 4160 6916
rect 3752 6876 3758 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 4430 6916 4436 6928
rect 4391 6888 4436 6916
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2731 6820 2820 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1728 6752 1869 6780
rect 1728 6740 1734 6752
rect 1857 6749 1869 6752
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2424 6712 2452 6743
rect 2682 6712 2688 6724
rect 2424 6684 2688 6712
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 2792 6644 2820 6820
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 4246 6848 4252 6860
rect 3016 6820 4252 6848
rect 3016 6808 3022 6820
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 2869 6743 2927 6749
rect 2884 6712 2912 6743
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4356 6780 4384 6811
rect 4212 6752 4384 6780
rect 4540 6780 4568 6956
rect 10152 6956 12164 6984
rect 4801 6919 4859 6925
rect 4801 6885 4813 6919
rect 4847 6916 4859 6919
rect 5442 6916 5448 6928
rect 4847 6888 5448 6916
rect 4847 6885 4859 6888
rect 4801 6879 4859 6885
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 6822 6916 6828 6928
rect 5960 6888 6828 6916
rect 5960 6876 5966 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5592 6820 5641 6848
rect 5592 6808 5598 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 6730 6848 6736 6860
rect 6691 6820 6736 6848
rect 5629 6811 5687 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 5902 6780 5908 6792
rect 4540 6752 5908 6780
rect 4212 6740 4218 6752
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7926 6780 7932 6792
rect 7055 6752 7932 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9950 6780 9956 6792
rect 9815 6752 9956 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 2958 6712 2964 6724
rect 2884 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 8297 6715 8355 6721
rect 5132 6684 5488 6712
rect 5132 6672 5138 6684
rect 5460 6656 5488 6684
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 10152 6712 10180 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12526 6984 12532 6996
rect 12268 6956 12532 6984
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 10468 6888 11468 6916
rect 10468 6876 10474 6888
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11440 6857 11468 6888
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 11885 6919 11943 6925
rect 11885 6916 11897 6919
rect 11664 6888 11897 6916
rect 11664 6876 11670 6888
rect 11885 6885 11897 6888
rect 11931 6916 11943 6919
rect 12268 6916 12296 6956
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 14274 6984 14280 6996
rect 12860 6956 14280 6984
rect 12860 6944 12866 6956
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17552 6956 17601 6984
rect 17552 6944 17558 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 17589 6947 17647 6953
rect 12710 6916 12716 6928
rect 11931 6888 12296 6916
rect 12544 6888 12716 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 12544 6860 12572 6888
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 17126 6916 17132 6928
rect 16224 6888 17132 6916
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11112 6820 11161 6848
rect 11112 6808 11118 6820
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 8343 6684 10180 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 3050 6644 3056 6656
rect 2792 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6644 3114 6656
rect 3510 6644 3516 6656
rect 3108 6616 3516 6644
rect 3108 6604 3114 6616
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5500 6616 5825 6644
rect 5500 6604 5506 6616
rect 5813 6613 5825 6616
rect 5859 6613 5871 6647
rect 11164 6644 11192 6811
rect 11440 6780 11468 6811
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 13354 6848 13360 6860
rect 12636 6820 13360 6848
rect 12636 6780 12664 6820
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 15933 6851 15991 6857
rect 15933 6817 15945 6851
rect 15979 6848 15991 6851
rect 16224 6848 16252 6888
rect 17126 6876 17132 6888
rect 17184 6876 17190 6928
rect 15979 6820 16252 6848
rect 16301 6851 16359 6857
rect 15979 6817 15991 6820
rect 15933 6811 15991 6817
rect 16301 6817 16313 6851
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 16531 6820 17325 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 11440 6752 12664 6780
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12989 6783 13047 6789
rect 12768 6752 12813 6780
rect 12768 6740 12774 6752
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13170 6780 13176 6792
rect 13035 6752 13176 6780
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14182 6780 14188 6792
rect 13964 6752 14188 6780
rect 13964 6740 13970 6752
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6780 16083 6783
rect 16114 6780 16120 6792
rect 16071 6752 16120 6780
rect 16071 6749 16083 6752
rect 16025 6743 16083 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16316 6780 16344 6811
rect 16574 6780 16580 6792
rect 16316 6752 16580 6780
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 17328 6780 17356 6811
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17460 6820 17509 6848
rect 17460 6808 17466 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 18966 6780 18972 6792
rect 17328 6752 18972 6780
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 11241 6715 11299 6721
rect 11241 6681 11253 6715
rect 11287 6712 11299 6715
rect 11330 6712 11336 6724
rect 11287 6684 11336 6712
rect 11287 6681 11299 6684
rect 11241 6675 11299 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 13906 6644 13912 6656
rect 11164 6616 13912 6644
rect 5813 6607 5871 6613
rect 13906 6604 13912 6616
rect 13964 6644 13970 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13964 6616 14105 6644
rect 13964 6604 13970 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 14093 6607 14151 6613
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 1104 6554 24840 6576
rect 1104 6502 4947 6554
rect 4999 6502 5011 6554
rect 5063 6502 5075 6554
rect 5127 6502 5139 6554
rect 5191 6502 12878 6554
rect 12930 6502 12942 6554
rect 12994 6502 13006 6554
rect 13058 6502 13070 6554
rect 13122 6502 20808 6554
rect 20860 6502 20872 6554
rect 20924 6502 20936 6554
rect 20988 6502 21000 6554
rect 21052 6502 24840 6554
rect 1104 6480 24840 6502
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11606 6440 11612 6452
rect 10008 6412 11612 6440
rect 10008 6400 10014 6412
rect 11606 6400 11612 6412
rect 11664 6440 11670 6452
rect 11882 6440 11888 6452
rect 11664 6412 11888 6440
rect 11664 6400 11670 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12989 6443 13047 6449
rect 12989 6409 13001 6443
rect 13035 6440 13047 6443
rect 13170 6440 13176 6452
rect 13035 6412 13176 6440
rect 13035 6409 13047 6412
rect 12989 6403 13047 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 15194 6440 15200 6452
rect 13320 6412 15200 6440
rect 13320 6400 13326 6412
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 16574 6440 16580 6452
rect 16535 6412 16580 6440
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 2958 6372 2964 6384
rect 2919 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 7926 6372 7932 6384
rect 4304 6344 5120 6372
rect 7887 6344 7932 6372
rect 4304 6332 4310 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 2976 6304 3004 6332
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 2976 6276 4353 6304
rect 4341 6273 4353 6276
rect 4387 6304 4399 6307
rect 4430 6304 4436 6316
rect 4387 6276 4436 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 1394 6236 1400 6248
rect 1307 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 1762 6236 1768 6248
rect 1452 6208 1768 6236
rect 1452 6196 1458 6208
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4304 6208 4537 6236
rect 4304 6196 4310 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6236 4951 6239
rect 4982 6236 4988 6248
rect 4939 6208 4988 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5092 6245 5120 6344
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 10686 6372 10692 6384
rect 10152 6344 10692 6372
rect 10152 6316 10180 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 6086 6304 6092 6316
rect 5684 6276 6092 6304
rect 5684 6264 5690 6276
rect 6086 6264 6092 6276
rect 6144 6304 6150 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6144 6276 6929 6304
rect 6144 6264 6150 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 10134 6304 10140 6316
rect 10095 6276 10140 6304
rect 6917 6267 6975 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 11146 6304 11152 6316
rect 10612 6276 11152 6304
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 7006 6236 7012 6248
rect 6967 6208 7012 6236
rect 5077 6199 5135 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 7156 6208 7481 6236
rect 7156 6196 7162 6208
rect 7469 6205 7481 6208
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 2406 6128 2412 6180
rect 2464 6168 2470 6180
rect 6914 6168 6920 6180
rect 2464 6140 6920 6168
rect 2464 6128 2470 6140
rect 6914 6128 6920 6140
rect 6972 6168 6978 6180
rect 7576 6168 7604 6199
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10612 6245 10640 6276
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 13412 6276 13461 6304
rect 13412 6264 13418 6276
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 13998 6304 14004 6316
rect 13959 6276 14004 6304
rect 13449 6267 13507 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14332 6276 15025 6304
rect 14332 6264 14338 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15378 6304 15384 6316
rect 15335 6276 15384 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9916 6208 10241 6236
rect 9916 6196 9922 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10778 6236 10784 6248
rect 10739 6208 10784 6236
rect 10597 6199 10655 6205
rect 6972 6140 7604 6168
rect 9585 6171 9643 6177
rect 6972 6128 6978 6140
rect 9585 6137 9597 6171
rect 9631 6168 9643 6171
rect 9950 6168 9956 6180
rect 9631 6140 9956 6168
rect 9631 6137 9643 6140
rect 9585 6131 9643 6137
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10244 6168 10272 6199
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 13906 6236 13912 6248
rect 13867 6208 13912 6236
rect 13541 6199 13599 6205
rect 13446 6168 13452 6180
rect 10244 6140 13452 6168
rect 13446 6128 13452 6140
rect 13504 6128 13510 6180
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4430 6100 4436 6112
rect 4203 6072 4436 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4982 6100 4988 6112
rect 4580 6072 4988 6100
rect 4580 6060 4586 6072
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 11054 6100 11060 6112
rect 7524 6072 11060 6100
rect 7524 6060 7530 6072
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 13556 6100 13584 6199
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 15160 6208 18061 6236
rect 15160 6196 15166 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 15378 6100 15384 6112
rect 13556 6072 15384 6100
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 18138 6100 18144 6112
rect 18099 6072 18144 6100
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 1104 6010 24840 6032
rect 1104 5958 8912 6010
rect 8964 5958 8976 6010
rect 9028 5958 9040 6010
rect 9092 5958 9104 6010
rect 9156 5958 16843 6010
rect 16895 5958 16907 6010
rect 16959 5958 16971 6010
rect 17023 5958 17035 6010
rect 17087 5958 24840 6010
rect 1104 5936 24840 5958
rect 3050 5896 3056 5908
rect 3011 5868 3056 5896
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4890 5896 4896 5908
rect 4295 5868 4896 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4890 5856 4896 5868
rect 4948 5896 4954 5908
rect 5258 5896 5264 5908
rect 4948 5868 5264 5896
rect 4948 5856 4954 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 10962 5896 10968 5908
rect 9640 5868 10968 5896
rect 9640 5856 9646 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 18138 5896 18144 5908
rect 11112 5868 18144 5896
rect 11112 5856 11118 5868
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 4430 5828 4436 5840
rect 4391 5800 4436 5828
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 4798 5828 4804 5840
rect 4759 5800 4804 5828
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 5813 5831 5871 5837
rect 5813 5828 5825 5831
rect 5408 5800 5825 5828
rect 5408 5788 5414 5800
rect 5813 5797 5825 5800
rect 5859 5797 5871 5831
rect 6362 5828 6368 5840
rect 6323 5800 6368 5828
rect 5813 5791 5871 5797
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 7116 5800 7512 5828
rect 1486 5760 1492 5772
rect 1447 5732 1492 5760
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 2915 5732 4200 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4172 5692 4200 5732
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 5902 5760 5908 5772
rect 4396 5732 4441 5760
rect 5815 5732 5908 5760
rect 4396 5720 4402 5732
rect 5902 5720 5908 5732
rect 5960 5760 5966 5772
rect 7116 5760 7144 5800
rect 7484 5772 7512 5800
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11333 5831 11391 5837
rect 11333 5828 11345 5831
rect 11204 5800 11345 5828
rect 11204 5788 11210 5800
rect 11333 5797 11345 5800
rect 11379 5797 11391 5831
rect 16393 5831 16451 5837
rect 16393 5828 16405 5831
rect 11333 5791 11391 5797
rect 13648 5800 16405 5828
rect 5960 5732 7144 5760
rect 7377 5763 7435 5769
rect 5960 5720 5966 5732
rect 7377 5729 7389 5763
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 4430 5692 4436 5704
rect 4172 5664 4436 5692
rect 4065 5655 4123 5661
rect 4080 5624 4108 5655
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 7392 5692 7420 5723
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7929 5763 7987 5769
rect 7524 5732 7569 5760
rect 7524 5720 7530 5732
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 9950 5760 9956 5772
rect 7975 5732 9812 5760
rect 9911 5732 9956 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 5500 5664 7420 5692
rect 5500 5652 5506 5664
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9640 5664 9689 5692
rect 9640 5652 9646 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9784 5692 9812 5732
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 13262 5720 13268 5772
rect 13320 5720 13326 5772
rect 13648 5769 13676 5800
rect 16393 5797 16405 5800
rect 16439 5797 16451 5831
rect 16393 5791 16451 5797
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5729 13691 5763
rect 14001 5763 14059 5769
rect 14001 5760 14013 5763
rect 13633 5723 13691 5729
rect 13740 5732 14013 5760
rect 13280 5692 13308 5720
rect 9784 5664 13308 5692
rect 9677 5655 9735 5661
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 13412 5664 13553 5692
rect 13412 5652 13418 5664
rect 13541 5661 13553 5664
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 5350 5624 5356 5636
rect 4080 5596 5356 5624
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 5592 5596 7205 5624
rect 5592 5584 5598 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 13740 5624 13768 5732
rect 14001 5729 14013 5732
rect 14047 5729 14059 5763
rect 14001 5723 14059 5729
rect 14185 5763 14243 5769
rect 14185 5729 14197 5763
rect 14231 5760 14243 5763
rect 15194 5760 15200 5772
rect 14231 5732 15200 5760
rect 14231 5729 14243 5732
rect 14185 5723 14243 5729
rect 14016 5692 14044 5723
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 14458 5692 14464 5704
rect 14016 5664 14464 5692
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 15304 5692 15332 5723
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 16301 5763 16359 5769
rect 15436 5732 15481 5760
rect 15436 5720 15442 5732
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 14608 5664 15332 5692
rect 14608 5652 14614 5664
rect 7193 5587 7251 5593
rect 13004 5596 13768 5624
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 5626 5556 5632 5568
rect 5587 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 13004 5556 13032 5596
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 16316 5624 16344 5723
rect 14056 5596 16344 5624
rect 14056 5584 14062 5596
rect 10468 5528 13032 5556
rect 13081 5559 13139 5565
rect 10468 5516 10474 5528
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13354 5556 13360 5568
rect 13127 5528 13360 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 1104 5466 24840 5488
rect 1104 5414 4947 5466
rect 4999 5414 5011 5466
rect 5063 5414 5075 5466
rect 5127 5414 5139 5466
rect 5191 5414 12878 5466
rect 12930 5414 12942 5466
rect 12994 5414 13006 5466
rect 13058 5414 13070 5466
rect 13122 5414 20808 5466
rect 20860 5414 20872 5466
rect 20924 5414 20936 5466
rect 20988 5414 21000 5466
rect 21052 5414 24840 5466
rect 1104 5392 24840 5414
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 4338 5352 4344 5364
rect 3467 5324 4344 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6880 5324 7021 5352
rect 6880 5312 6886 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 7009 5315 7067 5321
rect 7116 5324 13001 5352
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 3694 5284 3700 5296
rect 2271 5256 3700 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 4154 5284 4160 5296
rect 3896 5256 4160 5284
rect 2958 5216 2964 5228
rect 2019 5188 2964 5216
rect 2019 5157 2047 5188
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3896 5225 3924 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 5166 5284 5172 5296
rect 4264 5256 5172 5284
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 3881 5179 3939 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 2019 5151 2087 5157
rect 2019 5120 2041 5151
rect 2029 5117 2041 5120
rect 2075 5117 2087 5151
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 2029 5111 2087 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4264 5148 4292 5256
rect 5166 5244 5172 5256
rect 5224 5284 5230 5296
rect 5534 5284 5540 5296
rect 5224 5256 5540 5284
rect 5224 5244 5230 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 5994 5244 6000 5296
rect 6052 5284 6058 5296
rect 7116 5284 7144 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 15657 5355 15715 5361
rect 15657 5352 15669 5355
rect 13504 5324 15669 5352
rect 13504 5312 13510 5324
rect 15657 5321 15669 5324
rect 15703 5321 15715 5355
rect 15657 5315 15715 5321
rect 6052 5256 7144 5284
rect 6052 5244 6058 5256
rect 8754 5244 8760 5296
rect 8812 5244 8818 5296
rect 14458 5284 14464 5296
rect 14419 5256 14464 5284
rect 14458 5244 14464 5256
rect 14516 5244 14522 5296
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5216 5963 5219
rect 8772 5216 8800 5244
rect 5951 5188 8800 5216
rect 9125 5219 9183 5225
rect 5951 5185 5963 5188
rect 5905 5179 5963 5185
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 11057 5219 11115 5225
rect 11057 5216 11069 5219
rect 9171 5188 11069 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 11057 5185 11069 5188
rect 11103 5216 11115 5219
rect 13354 5216 13360 5228
rect 11103 5188 13216 5216
rect 13315 5188 13360 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 4203 5120 4292 5148
rect 5169 5151 5227 5157
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5350 5148 5356 5160
rect 5311 5120 5356 5148
rect 5169 5111 5227 5117
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 5184 5080 5212 5111
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 5258 5080 5264 5092
rect 2648 5052 5264 5080
rect 2648 5040 2654 5052
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 5460 5080 5488 5111
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5592 5120 6837 5148
rect 5592 5108 5598 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 8803 5120 10272 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 5902 5080 5908 5092
rect 5460 5052 5908 5080
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5049 8631 5083
rect 8573 5043 8631 5049
rect 9953 5083 10011 5089
rect 9953 5049 9965 5083
rect 9999 5080 10011 5083
rect 10134 5080 10140 5092
rect 9999 5052 10140 5080
rect 9999 5049 10011 5052
rect 9953 5043 10011 5049
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4338 5012 4344 5024
rect 3936 4984 4344 5012
rect 3936 4972 3942 4984
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 8588 5012 8616 5043
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 10244 5080 10272 5120
rect 10318 5108 10324 5160
rect 10376 5148 10382 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10376 5120 10609 5148
rect 10376 5108 10382 5120
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 10965 5151 11023 5157
rect 10744 5120 10789 5148
rect 10744 5108 10750 5120
rect 10965 5117 10977 5151
rect 11011 5148 11023 5151
rect 11238 5148 11244 5160
rect 11011 5120 11244 5148
rect 11011 5117 11023 5120
rect 10965 5111 11023 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12710 5148 12716 5160
rect 12400 5120 12716 5148
rect 12400 5108 12406 5120
rect 12710 5108 12716 5120
rect 12768 5148 12774 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12768 5120 13093 5148
rect 12768 5108 12774 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13188 5148 13216 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 13188 5120 15577 5148
rect 13081 5111 13139 5117
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 11054 5080 11060 5092
rect 10244 5052 11060 5080
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 18598 5080 18604 5092
rect 14016 5052 18604 5080
rect 10778 5012 10784 5024
rect 8588 4984 10784 5012
rect 10778 4972 10784 4984
rect 10836 5012 10842 5024
rect 12158 5012 12164 5024
rect 10836 4984 12164 5012
rect 10836 4972 10842 4984
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 14016 5012 14044 5052
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 13035 4984 14044 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 1104 4922 24840 4944
rect 1104 4870 8912 4922
rect 8964 4870 8976 4922
rect 9028 4870 9040 4922
rect 9092 4870 9104 4922
rect 9156 4870 16843 4922
rect 16895 4870 16907 4922
rect 16959 4870 16971 4922
rect 17023 4870 17035 4922
rect 17087 4870 24840 4922
rect 1104 4848 24840 4870
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9824 4780 9873 4808
rect 9824 4768 9830 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12032 4780 12357 4808
rect 12032 4768 12038 4780
rect 12345 4777 12357 4780
rect 12391 4777 12403 4811
rect 12345 4771 12403 4777
rect 4709 4743 4767 4749
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 5261 4743 5319 4749
rect 4755 4712 5212 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 2958 4672 2964 4684
rect 2919 4644 2964 4672
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 4154 4672 4160 4684
rect 3191 4644 4160 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 5184 4672 5212 4712
rect 5261 4709 5273 4743
rect 5307 4740 5319 4743
rect 5534 4740 5540 4752
rect 5307 4712 5540 4740
rect 5307 4709 5319 4712
rect 5261 4703 5319 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 12360 4740 12388 4771
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13228 4780 14228 4808
rect 13228 4768 13234 4780
rect 14200 4752 14228 4780
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14826 4808 14832 4820
rect 14424 4780 14832 4808
rect 14424 4768 14430 4780
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15565 4811 15623 4817
rect 15565 4808 15577 4811
rect 15252 4780 15577 4808
rect 15252 4768 15258 4780
rect 15565 4777 15577 4780
rect 15611 4808 15623 4811
rect 16022 4808 16028 4820
rect 15611 4780 16028 4808
rect 15611 4777 15623 4780
rect 15565 4771 15623 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 13449 4743 13507 4749
rect 7064 4712 9720 4740
rect 12360 4712 13032 4740
rect 7064 4700 7070 4712
rect 5350 4672 5356 4684
rect 4856 4644 4901 4672
rect 5184 4644 5356 4672
rect 4856 4632 4862 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6638 4672 6644 4684
rect 6512 4644 6644 4672
rect 6512 4632 6518 4644
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 6914 4672 6920 4684
rect 6871 4644 6920 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 6914 4632 6920 4644
rect 6972 4672 6978 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6972 4644 7389 4672
rect 6972 4632 6978 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 8478 4672 8484 4684
rect 7607 4644 8484 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9692 4681 9720 4712
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 13004 4672 13032 4712
rect 13449 4709 13461 4743
rect 13495 4740 13507 4743
rect 13722 4740 13728 4752
rect 13495 4712 13728 4740
rect 13495 4709 13507 4712
rect 13449 4703 13507 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 15289 4743 15347 4749
rect 15289 4740 15301 4743
rect 14240 4712 15301 4740
rect 14240 4700 14246 4712
rect 15289 4709 15301 4712
rect 15335 4709 15347 4743
rect 15289 4703 15347 4709
rect 13354 4672 13360 4684
rect 13004 4644 13360 4672
rect 9677 4635 9735 4641
rect 13354 4632 13360 4644
rect 13412 4672 13418 4684
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13412 4644 13645 4672
rect 13412 4632 13418 4644
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 13872 4644 15485 4672
rect 13872 4632 13878 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 23017 4675 23075 4681
rect 23017 4641 23029 4675
rect 23063 4672 23075 4675
rect 23934 4672 23940 4684
rect 23063 4644 23940 4672
rect 23063 4641 23075 4644
rect 23017 4635 23075 4641
rect 23934 4632 23940 4644
rect 23992 4632 23998 4684
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 3844 4576 4537 4604
rect 3844 4564 3850 4576
rect 4525 4573 4537 4576
rect 4571 4604 4583 4607
rect 5626 4604 5632 4616
rect 4571 4576 5632 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 10962 4604 10968 4616
rect 10923 4576 10968 4604
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11238 4604 11244 4616
rect 11199 4576 11244 4604
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12158 4564 12164 4616
rect 12216 4604 12222 4616
rect 13998 4604 14004 4616
rect 12216 4576 14004 4604
rect 12216 4564 12222 4576
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4604 23443 4607
rect 23566 4604 23572 4616
rect 23431 4576 23572 4604
rect 23431 4573 23443 4576
rect 23385 4567 23443 4573
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 23182 4539 23240 4545
rect 23182 4505 23194 4539
rect 23228 4536 23240 4539
rect 24302 4536 24308 4548
rect 23228 4508 24308 4536
rect 23228 4505 23240 4508
rect 23182 4499 23240 4505
rect 24302 4496 24308 4508
rect 24360 4496 24366 4548
rect 7834 4468 7840 4480
rect 7795 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 23290 4468 23296 4480
rect 23251 4440 23296 4468
rect 23290 4428 23296 4440
rect 23348 4428 23354 4480
rect 23382 4428 23388 4480
rect 23440 4468 23446 4480
rect 23477 4471 23535 4477
rect 23477 4468 23489 4471
rect 23440 4440 23489 4468
rect 23440 4428 23446 4440
rect 23477 4437 23489 4440
rect 23523 4437 23535 4471
rect 23477 4431 23535 4437
rect 1104 4378 24840 4400
rect 1104 4326 4947 4378
rect 4999 4326 5011 4378
rect 5063 4326 5075 4378
rect 5127 4326 5139 4378
rect 5191 4326 12878 4378
rect 12930 4326 12942 4378
rect 12994 4326 13006 4378
rect 13058 4326 13070 4378
rect 13122 4326 20808 4378
rect 20860 4326 20872 4378
rect 20924 4326 20936 4378
rect 20988 4326 21000 4378
rect 21052 4326 24840 4378
rect 1104 4304 24840 4326
rect 3421 4267 3479 4273
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 4154 4264 4160 4276
rect 3467 4236 4160 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 18598 4264 18604 4276
rect 18559 4236 18604 4264
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 22278 4196 22284 4208
rect 3752 4168 4752 4196
rect 22239 4168 22284 4196
rect 3752 4156 3758 4168
rect 750 4088 756 4140
rect 808 4128 814 4140
rect 1486 4128 1492 4140
rect 808 4100 1492 4128
rect 808 4088 814 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 3786 4128 3792 4140
rect 2280 4100 3792 4128
rect 2280 4088 2286 4100
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 4724 4128 4752 4168
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 4724 4100 4936 4128
rect 106 4020 112 4072
rect 164 4060 170 4072
rect 1302 4060 1308 4072
rect 164 4032 1308 4060
rect 164 4020 170 4032
rect 1302 4020 1308 4032
rect 1360 4020 1366 4072
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 4724 4069 4752 4100
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4908 4060 4936 4100
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 6880 4100 7573 4128
rect 6880 4088 6886 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7834 4128 7840 4140
rect 7795 4100 7840 4128
rect 7561 4091 7619 4097
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9858 4128 9864 4140
rect 9263 4100 9864 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 10410 4128 10416 4140
rect 9916 4100 10416 4128
rect 9916 4088 9922 4100
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 11296 4100 12449 4128
rect 11296 4088 11302 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12437 4091 12495 4097
rect 12986 4088 12992 4100
rect 13044 4128 13050 4140
rect 13262 4128 13268 4140
rect 13044 4100 13268 4128
rect 13044 4088 13050 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 14550 4088 14556 4140
rect 14608 4137 14614 4140
rect 14608 4131 14666 4137
rect 14608 4097 14620 4131
rect 14654 4097 14666 4131
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 14608 4091 14666 4097
rect 14608 4088 14614 4091
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15102 4128 15108 4140
rect 15063 4100 15108 4128
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 22186 4137 22192 4140
rect 22152 4131 22192 4137
rect 22152 4097 22164 4131
rect 22152 4091 22192 4097
rect 22186 4088 22192 4091
rect 22244 4088 22250 4140
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 5261 4063 5319 4069
rect 5261 4060 5273 4063
rect 4908 4032 5273 4060
rect 4801 4023 4859 4029
rect 5261 4029 5273 4032
rect 5307 4029 5319 4063
rect 5261 4023 5319 4029
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5718 4060 5724 4072
rect 5491 4032 5724 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 4816 3992 4844 4023
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 8720 4032 10057 4060
rect 8720 4020 8726 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10275 4032 10793 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11606 4060 11612 4072
rect 11011 4032 11612 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 6362 3992 6368 4004
rect 4816 3964 6368 3992
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 10244 3992 10272 4023
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13412 4032 13461 4060
rect 13412 4020 13418 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 13722 4060 13728 4072
rect 13679 4032 13728 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14691 4063 14749 4069
rect 14691 4029 14703 4063
rect 14737 4060 14749 4063
rect 14918 4060 14924 4072
rect 14737 4032 14924 4060
rect 14737 4029 14749 4032
rect 14691 4023 14749 4029
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4060 18567 4063
rect 22480 4060 22508 4091
rect 18555 4032 22508 4060
rect 18555 4029 18567 4032
rect 18509 4023 18567 4029
rect 9824 3964 10272 3992
rect 14461 3995 14519 4001
rect 9824 3952 9830 3964
rect 14461 3961 14473 3995
rect 14507 3992 14519 3995
rect 15010 3992 15016 4004
rect 14507 3964 15016 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 18325 3995 18383 4001
rect 18325 3961 18337 3995
rect 18371 3961 18383 3995
rect 18325 3955 18383 3961
rect 22005 3995 22063 4001
rect 22005 3961 22017 3995
rect 22051 3992 22063 3995
rect 23382 3992 23388 4004
rect 22051 3964 23388 3992
rect 22051 3961 22063 3964
rect 22005 3955 22063 3961
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10008 3896 11253 3924
rect 10008 3884 10014 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 11241 3887 11299 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 18340 3924 18368 3955
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 18506 3924 18512 3936
rect 18340 3896 18512 3924
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 23014 3924 23020 3936
rect 22244 3896 23020 3924
rect 22244 3884 22250 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 1104 3834 24840 3856
rect 1104 3782 8912 3834
rect 8964 3782 8976 3834
rect 9028 3782 9040 3834
rect 9092 3782 9104 3834
rect 9156 3782 16843 3834
rect 16895 3782 16907 3834
rect 16959 3782 16971 3834
rect 17023 3782 17035 3834
rect 17087 3782 24840 3834
rect 1104 3760 24840 3782
rect 4525 3723 4583 3729
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 4798 3720 4804 3732
rect 4571 3692 4804 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 8113 3723 8171 3729
rect 8113 3720 8125 3723
rect 4908 3692 8125 3720
rect 4908 3652 4936 3692
rect 8113 3689 8125 3692
rect 8159 3720 8171 3723
rect 8202 3720 8208 3732
rect 8159 3692 8208 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11204 3692 11253 3720
rect 11204 3680 11210 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 13136 3692 14289 3720
rect 13136 3680 13142 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 22370 3680 22376 3732
rect 22428 3720 22434 3732
rect 22833 3723 22891 3729
rect 22833 3720 22845 3723
rect 22428 3692 22845 3720
rect 22428 3680 22434 3692
rect 22833 3689 22845 3692
rect 22879 3689 22891 3723
rect 22833 3683 22891 3689
rect 2976 3624 4936 3652
rect 7101 3655 7159 3661
rect 2682 3584 2688 3596
rect 2643 3556 2688 3584
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 2976 3593 3004 3624
rect 7101 3621 7113 3655
rect 7147 3652 7159 3655
rect 7282 3652 7288 3664
rect 7147 3624 7288 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 16114 3652 16120 3664
rect 12820 3624 16120 3652
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3584 3203 3587
rect 4062 3584 4068 3596
rect 3191 3556 4068 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4522 3584 4528 3596
rect 4387 3556 4528 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 9766 3544 9772 3596
rect 9824 3544 9830 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 12820 3593 12848 3624
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 22189 3655 22247 3661
rect 22189 3621 22201 3655
rect 22235 3652 22247 3655
rect 22554 3652 22560 3664
rect 22235 3624 22560 3652
rect 22235 3621 22247 3624
rect 22189 3615 22247 3621
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 12986 3584 12992 3596
rect 12943 3556 12992 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 13814 3584 13820 3596
rect 13219 3556 13820 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 6822 3516 6828 3528
rect 5491 3488 6828 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 9784 3516 9812 3544
rect 10870 3516 10876 3528
rect 9723 3488 10876 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11330 3516 11336 3528
rect 11020 3488 11336 3516
rect 11020 3476 11026 3488
rect 11330 3476 11336 3488
rect 11388 3516 11394 3528
rect 13188 3516 13216 3547
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 14056 3556 14197 3584
rect 14056 3544 14062 3556
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 14550 3544 14556 3596
rect 14608 3584 14614 3596
rect 15286 3584 15292 3596
rect 14608 3556 15292 3584
rect 14608 3544 14614 3556
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 16666 3584 16672 3596
rect 16627 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 18230 3584 18236 3596
rect 18191 3556 18236 3584
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 11388 3488 13216 3516
rect 11388 3476 11394 3488
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13320 3488 13365 3516
rect 13320 3476 13326 3488
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16540 3488 17049 3516
rect 16540 3476 16546 3488
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 18380 3519 18438 3525
rect 18380 3485 18392 3519
rect 18426 3516 18438 3519
rect 18506 3516 18512 3528
rect 18426 3488 18512 3516
rect 18426 3485 18438 3488
rect 18380 3479 18438 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 16834 3451 16892 3457
rect 16834 3417 16846 3451
rect 16880 3448 16892 3451
rect 17218 3448 17224 3460
rect 16880 3420 17224 3448
rect 16880 3417 16892 3420
rect 16834 3411 16892 3417
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 18616 3448 18644 3479
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22152 3488 22569 3516
rect 22152 3476 22158 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 17920 3420 18644 3448
rect 17920 3408 17926 3420
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22465 3451 22523 3457
rect 22465 3448 22477 3451
rect 21876 3420 22477 3448
rect 21876 3408 21882 3420
rect 22465 3417 22477 3420
rect 22511 3417 22523 3451
rect 22465 3411 22523 3417
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 3602 3380 3608 3392
rect 1452 3352 3608 3380
rect 1452 3340 1458 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 10318 3380 10324 3392
rect 6512 3352 10324 3380
rect 6512 3340 6518 3352
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12710 3380 12716 3392
rect 12299 3352 12716 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 15378 3380 15384 3392
rect 15339 3352 15384 3380
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 16945 3383 17003 3389
rect 16945 3380 16957 3383
rect 16172 3352 16957 3380
rect 16172 3340 16178 3352
rect 16945 3349 16957 3352
rect 16991 3349 17003 3383
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 16945 3343 17003 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 17552 3352 18521 3380
rect 17552 3340 17558 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 18690 3380 18696 3392
rect 18651 3352 18696 3380
rect 18509 3343 18567 3349
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 22354 3383 22412 3389
rect 22354 3349 22366 3383
rect 22400 3380 22412 3383
rect 22922 3380 22928 3392
rect 22400 3352 22928 3380
rect 22400 3349 22412 3352
rect 22354 3343 22412 3349
rect 22922 3340 22928 3352
rect 22980 3340 22986 3392
rect 1104 3290 24840 3312
rect 1104 3238 4947 3290
rect 4999 3238 5011 3290
rect 5063 3238 5075 3290
rect 5127 3238 5139 3290
rect 5191 3238 12878 3290
rect 12930 3238 12942 3290
rect 12994 3238 13006 3290
rect 13058 3238 13070 3290
rect 13122 3238 20808 3290
rect 20860 3238 20872 3290
rect 20924 3238 20936 3290
rect 20988 3238 21000 3290
rect 21052 3238 24840 3290
rect 1104 3216 24840 3238
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 4062 3176 4068 3188
rect 3016 3148 3648 3176
rect 4023 3148 4068 3176
rect 3016 3136 3022 3148
rect 3620 3108 3648 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 5258 3176 5264 3188
rect 5215 3148 5264 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 5184 3108 5212 3139
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7340 3148 8432 3176
rect 7340 3136 7346 3148
rect 3620 3080 5212 3108
rect 8404 3108 8432 3148
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 8536 3148 10057 3176
rect 8536 3136 8542 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 15086 3179 15144 3185
rect 10376 3148 14007 3176
rect 10376 3136 10382 3148
rect 12434 3108 12440 3120
rect 8404 3080 12440 3108
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 13814 3108 13820 3120
rect 13775 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2188 3012 2973 3040
rect 2188 3000 2194 3012
rect 2961 3009 2973 3012
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5905 3043 5963 3049
rect 4856 3012 5488 3040
rect 4856 3000 4862 3012
rect 1118 2932 1124 2984
rect 1176 2972 1182 2984
rect 1489 2975 1547 2981
rect 1489 2972 1501 2975
rect 1176 2944 1501 2972
rect 1176 2932 1182 2944
rect 1489 2941 1501 2944
rect 1535 2941 1547 2975
rect 1489 2935 1547 2941
rect 1854 2932 1860 2984
rect 1912 2972 1918 2984
rect 5460 2981 5488 3012
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 7926 3040 7932 3052
rect 5951 3012 7932 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 12710 3040 12716 3052
rect 9171 3012 10971 3040
rect 12671 3012 12716 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 10943 2984 10971 3012
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 1912 2944 2697 2972
rect 1912 2932 1918 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 6880 2944 7481 2972
rect 6880 2932 6886 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7469 2935 7527 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9916 2944 9965 2972
rect 9916 2932 9922 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 10943 2972 10968 2984
rect 10875 2944 10968 2972
rect 9953 2935 10011 2941
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 13979 2972 14007 3148
rect 15086 3145 15098 3179
rect 15132 3176 15144 3179
rect 15378 3176 15384 3188
rect 15132 3148 15384 3176
rect 15132 3145 15144 3148
rect 15086 3139 15144 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19337 3179 19395 3185
rect 19337 3176 19349 3179
rect 19024 3148 19349 3176
rect 19024 3136 19030 3148
rect 19337 3145 19349 3148
rect 19383 3145 19395 3179
rect 19337 3139 19395 3145
rect 21545 3179 21603 3185
rect 21545 3145 21557 3179
rect 21591 3176 21603 3179
rect 22278 3176 22284 3188
rect 21591 3148 22284 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 14918 3108 14924 3120
rect 14700 3080 14924 3108
rect 14700 3068 14706 3080
rect 14918 3068 14924 3080
rect 14976 3108 14982 3120
rect 15197 3111 15255 3117
rect 15197 3108 15209 3111
rect 14976 3080 15209 3108
rect 14976 3068 14982 3080
rect 15197 3077 15209 3080
rect 15243 3077 15255 3111
rect 15197 3071 15255 3077
rect 19226 3111 19284 3117
rect 19226 3077 19238 3111
rect 19272 3108 19284 3111
rect 20070 3108 20076 3120
rect 19272 3080 20076 3108
rect 19272 3077 19284 3080
rect 19226 3071 19284 3077
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 20346 3068 20352 3120
rect 20404 3108 20410 3120
rect 21177 3111 21235 3117
rect 21177 3108 21189 3111
rect 20404 3080 21189 3108
rect 20404 3068 20410 3080
rect 21177 3077 21189 3080
rect 21223 3077 21235 3111
rect 21177 3071 21235 3077
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 15102 3040 15108 3052
rect 14884 3012 15108 3040
rect 14884 3000 14890 3012
rect 15102 3000 15108 3012
rect 15160 3040 15166 3052
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15160 3012 15301 3040
rect 15160 3000 15166 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3009 15439 3043
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 15381 3003 15439 3009
rect 19352 3012 19441 3040
rect 15396 2972 15424 3003
rect 19352 2984 19380 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20772 3012 21281 3040
rect 20772 3000 20778 3012
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 13979 2944 15424 2972
rect 12437 2935 12495 2941
rect 19334 2932 19340 2984
rect 19392 2932 19398 2984
rect 21048 2975 21106 2981
rect 21048 2941 21060 2975
rect 21094 2972 21106 2975
rect 21450 2972 21456 2984
rect 21094 2944 21456 2972
rect 21094 2941 21106 2944
rect 21048 2935 21106 2941
rect 21450 2932 21456 2944
rect 21508 2932 21514 2984
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2972 22615 2975
rect 24670 2972 24676 2984
rect 22603 2944 24676 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 24670 2932 24676 2944
rect 24728 2932 24734 2984
rect 5350 2904 5356 2916
rect 5311 2876 5356 2904
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 14921 2907 14979 2913
rect 14921 2873 14933 2907
rect 14967 2904 14979 2907
rect 15378 2904 15384 2916
rect 14967 2876 15384 2904
rect 14967 2873 14979 2876
rect 14921 2867 14979 2873
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 19061 2907 19119 2913
rect 19061 2873 19073 2907
rect 19107 2904 19119 2907
rect 19610 2904 19616 2916
rect 19107 2876 19616 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 20901 2907 20959 2913
rect 20901 2873 20913 2907
rect 20947 2904 20959 2907
rect 21174 2904 21180 2916
rect 20947 2876 21180 2904
rect 20947 2873 20959 2876
rect 20901 2867 20959 2873
rect 21174 2864 21180 2876
rect 21232 2864 21238 2916
rect 22370 2864 22376 2916
rect 22428 2904 22434 2916
rect 25406 2904 25412 2916
rect 22428 2876 25412 2904
rect 22428 2864 22434 2876
rect 25406 2864 25412 2876
rect 25464 2864 25470 2916
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 1946 2836 1952 2848
rect 1627 2808 1952 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 1946 2796 1952 2808
rect 2004 2796 2010 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 11057 2839 11115 2845
rect 11057 2836 11069 2839
rect 8076 2808 11069 2836
rect 8076 2796 8082 2808
rect 11057 2805 11069 2808
rect 11103 2805 11115 2839
rect 11057 2799 11115 2805
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 15286 2836 15292 2848
rect 13964 2808 15292 2836
rect 13964 2796 13970 2808
rect 15286 2796 15292 2808
rect 15344 2836 15350 2848
rect 15746 2836 15752 2848
rect 15344 2808 15752 2836
rect 15344 2796 15350 2808
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 19702 2836 19708 2848
rect 19663 2808 19708 2836
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 22649 2839 22707 2845
rect 22649 2805 22661 2839
rect 22695 2836 22707 2839
rect 22738 2836 22744 2848
rect 22695 2808 22744 2836
rect 22695 2805 22707 2808
rect 22649 2799 22707 2805
rect 22738 2796 22744 2808
rect 22796 2796 22802 2848
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 25774 2836 25780 2848
rect 23440 2808 25780 2836
rect 23440 2796 23446 2808
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 1104 2746 24840 2768
rect 1104 2694 8912 2746
rect 8964 2694 8976 2746
rect 9028 2694 9040 2746
rect 9092 2694 9104 2746
rect 9156 2694 16843 2746
rect 16895 2694 16907 2746
rect 16959 2694 16971 2746
rect 17023 2694 17035 2746
rect 17087 2694 24840 2746
rect 1104 2672 24840 2694
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7800 2604 8125 2632
rect 7800 2592 7806 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 8220 2604 10916 2632
rect 1578 2524 1584 2576
rect 1636 2564 1642 2576
rect 1857 2567 1915 2573
rect 1857 2564 1869 2567
rect 1636 2536 1869 2564
rect 1636 2524 1642 2536
rect 1857 2533 1869 2536
rect 1903 2533 1915 2567
rect 1857 2527 1915 2533
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2564 4491 2567
rect 5350 2564 5356 2576
rect 4479 2536 5356 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 5350 2524 5356 2536
rect 5408 2524 5414 2576
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 8220 2564 8248 2604
rect 5684 2536 8248 2564
rect 10888 2564 10916 2604
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 11204 2604 11253 2632
rect 11204 2592 11210 2604
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 12713 2635 12771 2641
rect 12713 2632 12725 2635
rect 11241 2595 11299 2601
rect 11348 2604 12725 2632
rect 11348 2564 11376 2604
rect 12713 2601 12725 2604
rect 12759 2601 12771 2635
rect 12713 2595 12771 2601
rect 15010 2592 15016 2644
rect 15068 2632 15074 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15068 2604 15577 2632
rect 15068 2592 15074 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 18969 2635 19027 2641
rect 18969 2632 18981 2635
rect 18656 2604 18981 2632
rect 18656 2592 18662 2604
rect 18969 2601 18981 2604
rect 19015 2601 19027 2635
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 18969 2595 19027 2601
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 10888 2536 11376 2564
rect 13817 2567 13875 2573
rect 5684 2524 5690 2536
rect 13817 2533 13829 2567
rect 13863 2564 13875 2567
rect 18325 2567 18383 2573
rect 13863 2536 15424 2564
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 15396 2508 15424 2536
rect 18325 2533 18337 2567
rect 18371 2564 18383 2567
rect 18690 2564 18696 2576
rect 18371 2536 18696 2564
rect 18371 2533 18383 2536
rect 18325 2527 18383 2533
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 22370 2564 22376 2576
rect 22331 2536 22376 2564
rect 22370 2524 22376 2536
rect 22428 2524 22434 2576
rect 1946 2456 1952 2508
rect 2004 2505 2010 2508
rect 2004 2499 2062 2505
rect 2004 2465 2016 2499
rect 2050 2465 2062 2499
rect 4246 2496 4252 2508
rect 2004 2459 2062 2465
rect 2148 2468 4252 2496
rect 2004 2456 2010 2459
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 2148 2428 2176 2468
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 4522 2496 4528 2508
rect 4435 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6454 2496 6460 2508
rect 5859 2468 6460 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 7064 2468 7113 2496
rect 7064 2456 7070 2468
rect 7101 2465 7113 2468
rect 7147 2496 7159 2499
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 7147 2468 7665 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7653 2465 7665 2468
rect 7699 2465 7711 2499
rect 7653 2459 7711 2465
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8018 2496 8024 2508
rect 7883 2468 8024 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9824 2468 9873 2496
rect 9824 2456 9830 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 10134 2496 10140 2508
rect 10095 2468 10140 2496
rect 9861 2459 9919 2465
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12492 2468 12633 2496
rect 12492 2456 12498 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13906 2456 13912 2508
rect 13964 2505 13970 2508
rect 13964 2499 14022 2505
rect 13964 2465 13976 2499
rect 14010 2465 14022 2499
rect 13964 2459 14022 2465
rect 13964 2456 13970 2459
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15436 2468 15485 2496
rect 15436 2456 15442 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 18472 2499 18530 2505
rect 18472 2465 18484 2499
rect 18518 2496 18530 2499
rect 19702 2496 19708 2508
rect 18518 2468 19708 2496
rect 18518 2465 18530 2468
rect 18472 2459 18530 2465
rect 19702 2456 19708 2468
rect 19760 2456 19766 2508
rect 21361 2499 21419 2505
rect 21361 2465 21373 2499
rect 21407 2465 21419 2499
rect 21361 2459 21419 2465
rect 22520 2499 22578 2505
rect 22520 2465 22532 2499
rect 22566 2496 22578 2499
rect 23382 2496 23388 2508
rect 22566 2468 23388 2496
rect 22566 2465 22578 2468
rect 22520 2459 22578 2465
rect 1912 2400 2176 2428
rect 2225 2431 2283 2437
rect 1912 2388 1918 2400
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2314 2428 2320 2440
rect 2271 2400 2320 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 4540 2428 4568 2456
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 4540 2400 5917 2428
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6420 2400 6929 2428
rect 6420 2388 6426 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2428 14243 2431
rect 15102 2428 15108 2440
rect 14231 2400 15108 2428
rect 14231 2397 14243 2400
rect 14185 2391 14243 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 17310 2388 17316 2440
rect 17368 2428 17374 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 17368 2400 18705 2428
rect 17368 2388 17374 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 2038 2320 2044 2372
rect 2096 2360 2102 2372
rect 2133 2363 2191 2369
rect 2133 2360 2145 2363
rect 2096 2332 2145 2360
rect 2096 2320 2102 2332
rect 2133 2329 2145 2332
rect 2179 2329 2191 2363
rect 2133 2323 2191 2329
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2360 14151 2363
rect 14642 2360 14648 2372
rect 14139 2332 14648 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4488 2264 4721 2292
rect 4488 2252 4494 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 14274 2292 14280 2304
rect 14235 2264 14280 2292
rect 4709 2255 4767 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 18598 2292 18604 2304
rect 18559 2264 18604 2292
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 21376 2292 21404 2459
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 22738 2428 22744 2440
rect 22699 2400 22744 2428
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 21453 2363 21511 2369
rect 21453 2329 21465 2363
rect 21499 2360 21511 2363
rect 22649 2363 22707 2369
rect 22649 2360 22661 2363
rect 21499 2332 22661 2360
rect 21499 2329 21511 2332
rect 21453 2323 21511 2329
rect 22649 2329 22661 2332
rect 22695 2329 22707 2363
rect 22649 2323 22707 2329
rect 25038 2292 25044 2304
rect 21376 2264 25044 2292
rect 25038 2252 25044 2264
rect 25096 2252 25102 2304
rect 1104 2202 24840 2224
rect 1104 2150 4947 2202
rect 4999 2150 5011 2202
rect 5063 2150 5075 2202
rect 5127 2150 5139 2202
rect 5191 2150 12878 2202
rect 12930 2150 12942 2202
rect 12994 2150 13006 2202
rect 13058 2150 13070 2202
rect 13122 2150 20808 2202
rect 20860 2150 20872 2202
rect 20924 2150 20936 2202
rect 20988 2150 21000 2202
rect 21052 2150 24840 2202
rect 1104 2128 24840 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 14274 2088 14280 2100
rect 2924 2060 14280 2088
rect 2924 2048 2930 2060
rect 14274 2048 14280 2060
rect 14332 2048 14338 2100
rect 2498 1980 2504 2032
rect 2556 2020 2562 2032
rect 18598 2020 18604 2032
rect 2556 1992 18604 2020
rect 2556 1980 2562 1992
rect 18598 1980 18604 1992
rect 18656 1980 18662 2032
rect 4614 1912 4620 1964
rect 4672 1952 4678 1964
rect 5074 1952 5080 1964
rect 4672 1924 5080 1952
rect 4672 1912 4678 1924
rect 5074 1912 5080 1924
rect 5132 1912 5138 1964
rect 12710 1300 12716 1352
rect 12768 1340 12774 1352
rect 13262 1340 13268 1352
rect 12768 1312 13268 1340
rect 12768 1300 12774 1312
rect 13262 1300 13268 1312
rect 13320 1300 13326 1352
rect 11146 960 11152 1012
rect 11204 1000 11210 1012
rect 12066 1000 12072 1012
rect 11204 972 12072 1000
rect 11204 960 11210 972
rect 12066 960 12072 972
rect 12124 960 12130 1012
<< via1 >>
rect 22100 49104 22152 49156
rect 23204 49104 23256 49156
rect 8912 47302 8964 47354
rect 8976 47302 9028 47354
rect 9040 47302 9092 47354
rect 9104 47302 9156 47354
rect 16843 47302 16895 47354
rect 16907 47302 16959 47354
rect 16971 47302 17023 47354
rect 17035 47302 17087 47354
rect 8208 47064 8260 47116
rect 11244 47200 11296 47252
rect 12164 47200 12216 47252
rect 21180 47200 21232 47252
rect 21640 47200 21692 47252
rect 3056 46928 3108 46980
rect 6276 46928 6328 46980
rect 12532 47064 12584 47116
rect 13820 47132 13872 47184
rect 14556 47132 14608 47184
rect 14004 47107 14056 47116
rect 14004 47073 14013 47107
rect 14013 47073 14047 47107
rect 14047 47073 14056 47107
rect 14004 47064 14056 47073
rect 14188 47107 14240 47116
rect 14188 47073 14197 47107
rect 14197 47073 14231 47107
rect 14231 47073 14240 47107
rect 14188 47064 14240 47073
rect 15660 47107 15712 47116
rect 15660 47073 15669 47107
rect 15669 47073 15703 47107
rect 15703 47073 15712 47107
rect 15660 47064 15712 47073
rect 15752 47107 15804 47116
rect 15752 47073 15761 47107
rect 15761 47073 15795 47107
rect 15795 47073 15804 47107
rect 15752 47064 15804 47073
rect 12440 46996 12492 47048
rect 16212 47039 16264 47048
rect 16212 47005 16221 47039
rect 16221 47005 16255 47039
rect 16255 47005 16264 47039
rect 16212 46996 16264 47005
rect 2688 46860 2740 46912
rect 3332 46860 3384 46912
rect 10048 46903 10100 46912
rect 10048 46869 10057 46903
rect 10057 46869 10091 46903
rect 10091 46869 10100 46903
rect 10048 46860 10100 46869
rect 11428 46903 11480 46912
rect 11428 46869 11437 46903
rect 11437 46869 11471 46903
rect 11471 46869 11480 46903
rect 11428 46860 11480 46869
rect 12348 46860 12400 46912
rect 13728 46860 13780 46912
rect 14280 46903 14332 46912
rect 14280 46869 14289 46903
rect 14289 46869 14323 46903
rect 14323 46869 14332 46903
rect 14280 46860 14332 46869
rect 15476 46903 15528 46912
rect 15476 46869 15485 46903
rect 15485 46869 15519 46903
rect 15519 46869 15528 46903
rect 15476 46860 15528 46869
rect 19984 46860 20036 46912
rect 24032 46860 24084 46912
rect 4947 46758 4999 46810
rect 5011 46758 5063 46810
rect 5075 46758 5127 46810
rect 5139 46758 5191 46810
rect 12878 46758 12930 46810
rect 12942 46758 12994 46810
rect 13006 46758 13058 46810
rect 13070 46758 13122 46810
rect 20808 46758 20860 46810
rect 20872 46758 20924 46810
rect 20936 46758 20988 46810
rect 21000 46758 21052 46810
rect 1952 46656 2004 46708
rect 4344 46656 4396 46708
rect 10600 46656 10652 46708
rect 14188 46656 14240 46708
rect 17684 46656 17736 46708
rect 18420 46656 18472 46708
rect 25596 46656 25648 46708
rect 1124 46588 1176 46640
rect 5724 46588 5776 46640
rect 14832 46520 14884 46572
rect 5908 46452 5960 46504
rect 7656 46452 7708 46504
rect 8760 46452 8812 46504
rect 11152 46495 11204 46504
rect 11152 46461 11161 46495
rect 11161 46461 11195 46495
rect 11195 46461 11204 46495
rect 11152 46452 11204 46461
rect 14096 46495 14148 46504
rect 5448 46384 5500 46436
rect 12532 46384 12584 46436
rect 13176 46384 13228 46436
rect 5632 46359 5684 46368
rect 5632 46325 5641 46359
rect 5641 46325 5675 46359
rect 5675 46325 5684 46359
rect 5632 46316 5684 46325
rect 11336 46359 11388 46368
rect 11336 46325 11345 46359
rect 11345 46325 11379 46359
rect 11379 46325 11388 46359
rect 11336 46316 11388 46325
rect 12716 46359 12768 46368
rect 12716 46325 12725 46359
rect 12725 46325 12759 46359
rect 12759 46325 12768 46359
rect 12716 46316 12768 46325
rect 14096 46461 14105 46495
rect 14105 46461 14139 46495
rect 14139 46461 14148 46495
rect 14096 46452 14148 46461
rect 15476 46452 15528 46504
rect 17132 46452 17184 46504
rect 15384 46384 15436 46436
rect 16672 46384 16724 46436
rect 17960 46384 18012 46436
rect 20076 46384 20128 46436
rect 21364 46384 21416 46436
rect 24768 46384 24820 46436
rect 16120 46316 16172 46368
rect 8912 46214 8964 46266
rect 8976 46214 9028 46266
rect 9040 46214 9092 46266
rect 9104 46214 9156 46266
rect 16843 46214 16895 46266
rect 16907 46214 16959 46266
rect 16971 46214 17023 46266
rect 17035 46214 17087 46266
rect 5908 46112 5960 46164
rect 18512 46112 18564 46164
rect 22468 46112 22520 46164
rect 8208 46087 8260 46096
rect 8208 46053 8217 46087
rect 8217 46053 8251 46087
rect 8251 46053 8260 46087
rect 8208 46044 8260 46053
rect 12348 46087 12400 46096
rect 12348 46053 12357 46087
rect 12357 46053 12391 46087
rect 12391 46053 12400 46087
rect 12348 46044 12400 46053
rect 14280 46044 14332 46096
rect 10600 45976 10652 46028
rect 10784 45976 10836 46028
rect 13912 46019 13964 46028
rect 13912 45985 13921 46019
rect 13921 45985 13955 46019
rect 13955 45985 13964 46019
rect 13912 45976 13964 45985
rect 14832 45976 14884 46028
rect 16672 45976 16724 46028
rect 388 45908 440 45960
rect 2688 45908 2740 45960
rect 4804 45908 4856 45960
rect 5356 45908 5408 45960
rect 10968 45951 11020 45960
rect 10968 45917 10977 45951
rect 10977 45917 11011 45951
rect 11011 45917 11020 45951
rect 10968 45908 11020 45917
rect 15476 45840 15528 45892
rect 8484 45815 8536 45824
rect 8484 45781 8493 45815
rect 8493 45781 8527 45815
rect 8527 45781 8536 45815
rect 8484 45772 8536 45781
rect 13636 45815 13688 45824
rect 13636 45781 13645 45815
rect 13645 45781 13679 45815
rect 13679 45781 13688 45815
rect 13636 45772 13688 45781
rect 14096 45815 14148 45824
rect 14096 45781 14105 45815
rect 14105 45781 14139 45815
rect 14139 45781 14148 45815
rect 14096 45772 14148 45781
rect 15936 45772 15988 45824
rect 18236 46044 18288 46096
rect 4947 45670 4999 45722
rect 5011 45670 5063 45722
rect 5075 45670 5127 45722
rect 5139 45670 5191 45722
rect 12878 45670 12930 45722
rect 12942 45670 12994 45722
rect 13006 45670 13058 45722
rect 13070 45670 13122 45722
rect 20808 45670 20860 45722
rect 20872 45670 20924 45722
rect 20936 45670 20988 45722
rect 21000 45670 21052 45722
rect 5356 45568 5408 45620
rect 8760 45611 8812 45620
rect 8760 45577 8769 45611
rect 8769 45577 8803 45611
rect 8803 45577 8812 45611
rect 8760 45568 8812 45577
rect 13820 45611 13872 45620
rect 13820 45577 13829 45611
rect 13829 45577 13863 45611
rect 13863 45577 13872 45611
rect 13820 45568 13872 45577
rect 16120 45568 16172 45620
rect 11244 45543 11296 45552
rect 11244 45509 11253 45543
rect 11253 45509 11287 45543
rect 11287 45509 11296 45543
rect 11244 45500 11296 45509
rect 10784 45432 10836 45484
rect 13360 45432 13412 45484
rect 15660 45432 15712 45484
rect 4712 45364 4764 45416
rect 5264 45407 5316 45416
rect 5264 45373 5273 45407
rect 5273 45373 5307 45407
rect 5307 45373 5316 45407
rect 5264 45364 5316 45373
rect 5448 45364 5500 45416
rect 7472 45364 7524 45416
rect 7748 45364 7800 45416
rect 8484 45407 8536 45416
rect 8484 45373 8493 45407
rect 8493 45373 8527 45407
rect 8527 45373 8536 45407
rect 8484 45364 8536 45373
rect 10140 45407 10192 45416
rect 5632 45296 5684 45348
rect 8392 45296 8444 45348
rect 10140 45373 10149 45407
rect 10149 45373 10183 45407
rect 10183 45373 10192 45407
rect 10140 45364 10192 45373
rect 12532 45364 12584 45416
rect 14832 45364 14884 45416
rect 15200 45407 15252 45416
rect 15200 45373 15209 45407
rect 15209 45373 15243 45407
rect 15243 45373 15252 45407
rect 15200 45364 15252 45373
rect 18144 45364 18196 45416
rect 18328 45364 18380 45416
rect 18052 45339 18104 45348
rect 18052 45305 18061 45339
rect 18061 45305 18095 45339
rect 18095 45305 18104 45339
rect 18052 45296 18104 45305
rect 4804 45228 4856 45280
rect 8912 45126 8964 45178
rect 8976 45126 9028 45178
rect 9040 45126 9092 45178
rect 9104 45126 9156 45178
rect 16843 45126 16895 45178
rect 16907 45126 16959 45178
rect 16971 45126 17023 45178
rect 17035 45126 17087 45178
rect 7472 45024 7524 45076
rect 4804 44999 4856 45008
rect 4804 44965 4813 44999
rect 4813 44965 4847 44999
rect 4847 44965 4856 44999
rect 4804 44956 4856 44965
rect 10048 44956 10100 45008
rect 12440 45024 12492 45076
rect 12532 44956 12584 45008
rect 12716 44956 12768 45008
rect 15200 44956 15252 45008
rect 18144 44956 18196 45008
rect 4712 44931 4764 44940
rect 4712 44897 4721 44931
rect 4721 44897 4755 44931
rect 4755 44897 4764 44931
rect 4712 44888 4764 44897
rect 9220 44888 9272 44940
rect 11336 44931 11388 44940
rect 11336 44897 11345 44931
rect 11345 44897 11379 44931
rect 11379 44897 11388 44931
rect 11336 44888 11388 44897
rect 11520 44931 11572 44940
rect 11520 44897 11529 44931
rect 11529 44897 11563 44931
rect 11563 44897 11572 44931
rect 11520 44888 11572 44897
rect 12624 44888 12676 44940
rect 16212 44888 16264 44940
rect 5448 44820 5500 44872
rect 4160 44752 4212 44804
rect 4896 44752 4948 44804
rect 14832 44820 14884 44872
rect 10140 44727 10192 44736
rect 10140 44693 10149 44727
rect 10149 44693 10183 44727
rect 10183 44693 10192 44727
rect 10140 44684 10192 44693
rect 12716 44684 12768 44736
rect 13636 44684 13688 44736
rect 4947 44582 4999 44634
rect 5011 44582 5063 44634
rect 5075 44582 5127 44634
rect 5139 44582 5191 44634
rect 12878 44582 12930 44634
rect 12942 44582 12994 44634
rect 13006 44582 13058 44634
rect 13070 44582 13122 44634
rect 20808 44582 20860 44634
rect 20872 44582 20924 44634
rect 20936 44582 20988 44634
rect 21000 44582 21052 44634
rect 5356 44480 5408 44532
rect 9772 44480 9824 44532
rect 10968 44480 11020 44532
rect 11336 44412 11388 44464
rect 7656 44387 7708 44396
rect 7656 44353 7665 44387
rect 7665 44353 7699 44387
rect 7699 44353 7708 44387
rect 7656 44344 7708 44353
rect 4160 44276 4212 44328
rect 4804 44276 4856 44328
rect 5356 44276 5408 44328
rect 5540 44276 5592 44328
rect 7932 44319 7984 44328
rect 7932 44285 7941 44319
rect 7941 44285 7975 44319
rect 7975 44285 7984 44319
rect 7932 44276 7984 44285
rect 10416 44276 10468 44328
rect 15200 44480 15252 44532
rect 15476 44480 15528 44532
rect 13912 44319 13964 44328
rect 13912 44285 13921 44319
rect 13921 44285 13955 44319
rect 13955 44285 13964 44319
rect 13912 44276 13964 44285
rect 15936 44412 15988 44464
rect 15384 44344 15436 44396
rect 18328 44344 18380 44396
rect 15660 44276 15712 44328
rect 17868 44276 17920 44328
rect 3424 44251 3476 44260
rect 3424 44217 3433 44251
rect 3433 44217 3467 44251
rect 3467 44217 3476 44251
rect 3424 44208 3476 44217
rect 11428 44208 11480 44260
rect 12440 44208 12492 44260
rect 13176 44208 13228 44260
rect 5356 44140 5408 44192
rect 12808 44183 12860 44192
rect 12808 44149 12817 44183
rect 12817 44149 12851 44183
rect 12851 44149 12860 44183
rect 12808 44140 12860 44149
rect 16304 44208 16356 44260
rect 8912 44038 8964 44090
rect 8976 44038 9028 44090
rect 9040 44038 9092 44090
rect 9104 44038 9156 44090
rect 16843 44038 16895 44090
rect 16907 44038 16959 44090
rect 16971 44038 17023 44090
rect 17035 44038 17087 44090
rect 8208 43936 8260 43988
rect 3424 43868 3476 43920
rect 7380 43868 7432 43920
rect 8116 43868 8168 43920
rect 4712 43800 4764 43852
rect 6368 43843 6420 43852
rect 6368 43809 6377 43843
rect 6377 43809 6411 43843
rect 6411 43809 6420 43843
rect 6368 43800 6420 43809
rect 7656 43843 7708 43852
rect 7656 43809 7665 43843
rect 7665 43809 7699 43843
rect 7699 43809 7708 43843
rect 7656 43800 7708 43809
rect 13544 43936 13596 43988
rect 12808 43868 12860 43920
rect 17960 43868 18012 43920
rect 7564 43732 7616 43784
rect 4620 43664 4672 43716
rect 11428 43800 11480 43852
rect 13544 43843 13596 43852
rect 13544 43809 13553 43843
rect 13553 43809 13587 43843
rect 13587 43809 13596 43843
rect 13544 43800 13596 43809
rect 16304 43843 16356 43852
rect 11336 43732 11388 43784
rect 12256 43775 12308 43784
rect 12256 43741 12265 43775
rect 12265 43741 12299 43775
rect 12299 43741 12308 43775
rect 12256 43732 12308 43741
rect 12532 43732 12584 43784
rect 16304 43809 16313 43843
rect 16313 43809 16347 43843
rect 16347 43809 16356 43843
rect 16304 43800 16356 43809
rect 14096 43775 14148 43784
rect 14096 43741 14105 43775
rect 14105 43741 14139 43775
rect 14139 43741 14148 43775
rect 14096 43732 14148 43741
rect 14832 43732 14884 43784
rect 12440 43664 12492 43716
rect 4804 43596 4856 43648
rect 6920 43596 6972 43648
rect 7748 43596 7800 43648
rect 7932 43639 7984 43648
rect 7932 43605 7941 43639
rect 7941 43605 7975 43639
rect 7975 43605 7984 43639
rect 7932 43596 7984 43605
rect 10508 43596 10560 43648
rect 12716 43596 12768 43648
rect 4947 43494 4999 43546
rect 5011 43494 5063 43546
rect 5075 43494 5127 43546
rect 5139 43494 5191 43546
rect 12878 43494 12930 43546
rect 12942 43494 12994 43546
rect 13006 43494 13058 43546
rect 13070 43494 13122 43546
rect 20808 43494 20860 43546
rect 20872 43494 20924 43546
rect 20936 43494 20988 43546
rect 21000 43494 21052 43546
rect 11336 43392 11388 43444
rect 15292 43392 15344 43444
rect 18328 43435 18380 43444
rect 18328 43401 18337 43435
rect 18337 43401 18371 43435
rect 18371 43401 18380 43435
rect 18328 43392 18380 43401
rect 3516 43256 3568 43308
rect 3700 43231 3752 43240
rect 3700 43197 3709 43231
rect 3709 43197 3743 43231
rect 3743 43197 3752 43231
rect 3700 43188 3752 43197
rect 5356 43231 5408 43240
rect 5356 43197 5365 43231
rect 5365 43197 5399 43231
rect 5399 43197 5408 43231
rect 5356 43188 5408 43197
rect 7380 43188 7432 43240
rect 9312 43256 9364 43308
rect 8208 43188 8260 43240
rect 11612 43256 11664 43308
rect 12256 43256 12308 43308
rect 14096 43256 14148 43308
rect 10600 43231 10652 43240
rect 10600 43197 10609 43231
rect 10609 43197 10643 43231
rect 10643 43197 10652 43231
rect 10600 43188 10652 43197
rect 12808 43188 12860 43240
rect 13360 43188 13412 43240
rect 14832 43188 14884 43240
rect 17960 43188 18012 43240
rect 2596 43120 2648 43172
rect 5908 43163 5960 43172
rect 5908 43129 5917 43163
rect 5917 43129 5951 43163
rect 5951 43129 5960 43163
rect 5908 43120 5960 43129
rect 9496 43163 9548 43172
rect 9496 43129 9505 43163
rect 9505 43129 9539 43163
rect 9539 43129 9548 43163
rect 9496 43120 9548 43129
rect 10508 43163 10560 43172
rect 10508 43129 10517 43163
rect 10517 43129 10551 43163
rect 10551 43129 10560 43163
rect 10508 43120 10560 43129
rect 18052 43163 18104 43172
rect 3148 43052 3200 43104
rect 7748 43052 7800 43104
rect 18052 43129 18061 43163
rect 18061 43129 18095 43163
rect 18095 43129 18104 43163
rect 18052 43120 18104 43129
rect 12440 43052 12492 43104
rect 14280 43052 14332 43104
rect 16488 43052 16540 43104
rect 8912 42950 8964 43002
rect 8976 42950 9028 43002
rect 9040 42950 9092 43002
rect 9104 42950 9156 43002
rect 16843 42950 16895 43002
rect 16907 42950 16959 43002
rect 16971 42950 17023 43002
rect 17035 42950 17087 43002
rect 13452 42848 13504 42900
rect 4436 42780 4488 42832
rect 5356 42780 5408 42832
rect 8208 42823 8260 42832
rect 8208 42789 8217 42823
rect 8217 42789 8251 42823
rect 8251 42789 8260 42823
rect 8208 42780 8260 42789
rect 9588 42712 9640 42764
rect 12440 42755 12492 42764
rect 5356 42644 5408 42696
rect 5816 42687 5868 42696
rect 4620 42576 4672 42628
rect 4804 42576 4856 42628
rect 5816 42653 5825 42687
rect 5825 42653 5859 42687
rect 5859 42653 5868 42687
rect 5816 42644 5868 42653
rect 6644 42644 6696 42696
rect 9956 42687 10008 42696
rect 9956 42653 9965 42687
rect 9965 42653 9999 42687
rect 9999 42653 10008 42687
rect 9956 42644 10008 42653
rect 11612 42644 11664 42696
rect 12440 42721 12449 42755
rect 12449 42721 12483 42755
rect 12483 42721 12492 42755
rect 12440 42712 12492 42721
rect 15384 42755 15436 42764
rect 15384 42721 15393 42755
rect 15393 42721 15427 42755
rect 15427 42721 15436 42755
rect 15384 42712 15436 42721
rect 18328 42712 18380 42764
rect 3976 42508 4028 42560
rect 6828 42508 6880 42560
rect 7656 42508 7708 42560
rect 12808 42644 12860 42696
rect 16120 42644 16172 42696
rect 17040 42687 17092 42696
rect 14832 42576 14884 42628
rect 16580 42576 16632 42628
rect 17040 42653 17049 42687
rect 17049 42653 17083 42687
rect 17083 42653 17092 42687
rect 17040 42644 17092 42653
rect 12440 42508 12492 42560
rect 15568 42508 15620 42560
rect 21272 42712 21324 42764
rect 4947 42406 4999 42458
rect 5011 42406 5063 42458
rect 5075 42406 5127 42458
rect 5139 42406 5191 42458
rect 12878 42406 12930 42458
rect 12942 42406 12994 42458
rect 13006 42406 13058 42458
rect 13070 42406 13122 42458
rect 20808 42406 20860 42458
rect 20872 42406 20924 42458
rect 20936 42406 20988 42458
rect 21000 42406 21052 42458
rect 3700 42304 3752 42356
rect 4620 42304 4672 42356
rect 5816 42304 5868 42356
rect 9312 42304 9364 42356
rect 4160 42236 4212 42288
rect 4804 42236 4856 42288
rect 3424 42100 3476 42152
rect 3976 42100 4028 42152
rect 6920 42168 6972 42220
rect 7012 42168 7064 42220
rect 7472 42168 7524 42220
rect 11520 42168 11572 42220
rect 5356 42143 5408 42152
rect 5356 42109 5365 42143
rect 5365 42109 5399 42143
rect 5399 42109 5408 42143
rect 5356 42100 5408 42109
rect 5540 42100 5592 42152
rect 7840 42143 7892 42152
rect 7840 42109 7849 42143
rect 7849 42109 7883 42143
rect 7883 42109 7892 42143
rect 7840 42100 7892 42109
rect 10692 42100 10744 42152
rect 11336 42143 11388 42152
rect 11336 42109 11345 42143
rect 11345 42109 11379 42143
rect 11379 42109 11388 42143
rect 11336 42100 11388 42109
rect 13912 42304 13964 42356
rect 18052 42304 18104 42356
rect 15476 42236 15528 42288
rect 16028 42236 16080 42288
rect 13544 42211 13596 42220
rect 13544 42177 13553 42211
rect 13553 42177 13587 42211
rect 13587 42177 13596 42211
rect 13544 42168 13596 42177
rect 17040 42168 17092 42220
rect 14280 42100 14332 42152
rect 14648 42143 14700 42152
rect 14648 42109 14657 42143
rect 14657 42109 14691 42143
rect 14691 42109 14700 42143
rect 14648 42100 14700 42109
rect 16212 42143 16264 42152
rect 16212 42109 16221 42143
rect 16221 42109 16255 42143
rect 16255 42109 16264 42143
rect 16212 42100 16264 42109
rect 17868 42100 17920 42152
rect 14556 42075 14608 42084
rect 14556 42041 14565 42075
rect 14565 42041 14599 42075
rect 14599 42041 14608 42075
rect 14556 42032 14608 42041
rect 16120 42075 16172 42084
rect 16120 42041 16129 42075
rect 16129 42041 16163 42075
rect 16163 42041 16172 42075
rect 16120 42032 16172 42041
rect 16672 42075 16724 42084
rect 16672 42041 16681 42075
rect 16681 42041 16715 42075
rect 16715 42041 16724 42075
rect 16672 42032 16724 42041
rect 8912 41862 8964 41914
rect 8976 41862 9028 41914
rect 9040 41862 9092 41914
rect 9104 41862 9156 41914
rect 16843 41862 16895 41914
rect 16907 41862 16959 41914
rect 16971 41862 17023 41914
rect 17035 41862 17087 41914
rect 4252 41760 4304 41812
rect 14556 41760 14608 41812
rect 1952 41624 2004 41676
rect 2596 41667 2648 41676
rect 2596 41633 2605 41667
rect 2605 41633 2639 41667
rect 2639 41633 2648 41667
rect 2596 41624 2648 41633
rect 7748 41735 7800 41744
rect 7748 41701 7757 41735
rect 7757 41701 7791 41735
rect 7791 41701 7800 41735
rect 7748 41692 7800 41701
rect 9496 41692 9548 41744
rect 11336 41692 11388 41744
rect 7472 41624 7524 41676
rect 9680 41624 9732 41676
rect 11796 41667 11848 41676
rect 11796 41633 11805 41667
rect 11805 41633 11839 41667
rect 11839 41633 11848 41667
rect 11796 41624 11848 41633
rect 18328 41692 18380 41744
rect 21180 41692 21232 41744
rect 13176 41624 13228 41676
rect 4068 41556 4120 41608
rect 4160 41556 4212 41608
rect 4528 41599 4580 41608
rect 4528 41565 4537 41599
rect 4537 41565 4571 41599
rect 4571 41565 4580 41599
rect 4528 41556 4580 41565
rect 6920 41556 6972 41608
rect 7196 41556 7248 41608
rect 12532 41556 12584 41608
rect 14464 41624 14516 41676
rect 15384 41667 15436 41676
rect 15384 41633 15393 41667
rect 15393 41633 15427 41667
rect 15427 41633 15436 41667
rect 15384 41624 15436 41633
rect 15568 41667 15620 41676
rect 15568 41633 15577 41667
rect 15577 41633 15611 41667
rect 15611 41633 15620 41667
rect 15568 41624 15620 41633
rect 16672 41624 16724 41676
rect 14648 41556 14700 41608
rect 16580 41556 16632 41608
rect 14280 41488 14332 41540
rect 14832 41488 14884 41540
rect 4160 41420 4212 41472
rect 4436 41420 4488 41472
rect 7840 41420 7892 41472
rect 9956 41420 10008 41472
rect 4947 41318 4999 41370
rect 5011 41318 5063 41370
rect 5075 41318 5127 41370
rect 5139 41318 5191 41370
rect 12878 41318 12930 41370
rect 12942 41318 12994 41370
rect 13006 41318 13058 41370
rect 13070 41318 13122 41370
rect 20808 41318 20860 41370
rect 20872 41318 20924 41370
rect 20936 41318 20988 41370
rect 21000 41318 21052 41370
rect 3424 41259 3476 41268
rect 3424 41225 3433 41259
rect 3433 41225 3467 41259
rect 3467 41225 3476 41259
rect 3424 41216 3476 41225
rect 4620 41216 4672 41268
rect 7380 41216 7432 41268
rect 12716 41216 12768 41268
rect 17132 41216 17184 41268
rect 16212 41148 16264 41200
rect 4528 41080 4580 41132
rect 6828 41080 6880 41132
rect 2964 41055 3016 41064
rect 2964 41021 2973 41055
rect 2973 41021 3007 41055
rect 3007 41021 3016 41055
rect 2964 41012 3016 41021
rect 3148 41055 3200 41064
rect 3148 41021 3157 41055
rect 3157 41021 3191 41055
rect 3191 41021 3200 41055
rect 3148 41012 3200 41021
rect 3700 41012 3752 41064
rect 4804 41055 4856 41064
rect 4804 41021 4813 41055
rect 4813 41021 4847 41055
rect 4847 41021 4856 41055
rect 4804 41012 4856 41021
rect 7012 41055 7064 41064
rect 7012 41021 7021 41055
rect 7021 41021 7055 41055
rect 7055 41021 7064 41055
rect 7012 41012 7064 41021
rect 7288 41055 7340 41064
rect 7288 41021 7297 41055
rect 7297 41021 7331 41055
rect 7331 41021 7340 41055
rect 7288 41012 7340 41021
rect 12624 41080 12676 41132
rect 9864 41012 9916 41064
rect 11060 41012 11112 41064
rect 11336 41012 11388 41064
rect 11520 41055 11572 41064
rect 11520 41021 11529 41055
rect 11529 41021 11563 41055
rect 11563 41021 11572 41055
rect 11520 41012 11572 41021
rect 13268 41012 13320 41064
rect 14372 41055 14424 41064
rect 4068 40944 4120 40996
rect 11152 40944 11204 40996
rect 14372 41021 14381 41055
rect 14381 41021 14415 41055
rect 14415 41021 14424 41055
rect 14372 41012 14424 41021
rect 14464 41012 14516 41064
rect 16028 41055 16080 41064
rect 16028 41021 16037 41055
rect 16037 41021 16071 41055
rect 16071 41021 16080 41055
rect 16028 41012 16080 41021
rect 16212 41055 16264 41064
rect 16212 41021 16221 41055
rect 16221 41021 16255 41055
rect 16255 41021 16264 41055
rect 16212 41012 16264 41021
rect 16120 40987 16172 40996
rect 16120 40953 16129 40987
rect 16129 40953 16163 40987
rect 16163 40953 16172 40987
rect 16120 40944 16172 40953
rect 16672 40987 16724 40996
rect 16672 40953 16681 40987
rect 16681 40953 16715 40987
rect 16715 40953 16724 40987
rect 16672 40944 16724 40953
rect 8912 40774 8964 40826
rect 8976 40774 9028 40826
rect 9040 40774 9092 40826
rect 9104 40774 9156 40826
rect 16843 40774 16895 40826
rect 16907 40774 16959 40826
rect 16971 40774 17023 40826
rect 17035 40774 17087 40826
rect 4160 40672 4212 40724
rect 5908 40604 5960 40656
rect 7288 40604 7340 40656
rect 15384 40647 15436 40656
rect 15384 40613 15393 40647
rect 15393 40613 15427 40647
rect 15427 40613 15436 40647
rect 15384 40604 15436 40613
rect 3148 40536 3200 40588
rect 4436 40579 4488 40588
rect 4436 40545 4445 40579
rect 4445 40545 4479 40579
rect 4479 40545 4488 40579
rect 4436 40536 4488 40545
rect 4804 40579 4856 40588
rect 4804 40545 4813 40579
rect 4813 40545 4847 40579
rect 4847 40545 4856 40579
rect 4804 40536 4856 40545
rect 5356 40536 5408 40588
rect 6736 40579 6788 40588
rect 6736 40545 6745 40579
rect 6745 40545 6779 40579
rect 6779 40545 6788 40579
rect 6736 40536 6788 40545
rect 8208 40579 8260 40588
rect 8208 40545 8217 40579
rect 8217 40545 8251 40579
rect 8251 40545 8260 40579
rect 8208 40536 8260 40545
rect 8760 40579 8812 40588
rect 8760 40545 8769 40579
rect 8769 40545 8803 40579
rect 8803 40545 8812 40579
rect 8760 40536 8812 40545
rect 9864 40579 9916 40588
rect 9864 40545 9873 40579
rect 9873 40545 9907 40579
rect 9907 40545 9916 40579
rect 9864 40536 9916 40545
rect 11152 40579 11204 40588
rect 11152 40545 11161 40579
rect 11161 40545 11195 40579
rect 11195 40545 11204 40579
rect 11152 40536 11204 40545
rect 11520 40579 11572 40588
rect 11520 40545 11529 40579
rect 11529 40545 11563 40579
rect 11563 40545 11572 40579
rect 11520 40536 11572 40545
rect 12440 40536 12492 40588
rect 18512 40672 18564 40724
rect 16120 40604 16172 40656
rect 16672 40536 16724 40588
rect 7196 40468 7248 40520
rect 9680 40468 9732 40520
rect 12716 40468 12768 40520
rect 16580 40468 16632 40520
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 10048 40375 10100 40384
rect 10048 40341 10057 40375
rect 10057 40341 10091 40375
rect 10091 40341 10100 40375
rect 10048 40332 10100 40341
rect 13820 40332 13872 40384
rect 13912 40375 13964 40384
rect 13912 40341 13921 40375
rect 13921 40341 13955 40375
rect 13955 40341 13964 40375
rect 13912 40332 13964 40341
rect 14924 40332 14976 40384
rect 17868 40332 17920 40384
rect 4947 40230 4999 40282
rect 5011 40230 5063 40282
rect 5075 40230 5127 40282
rect 5139 40230 5191 40282
rect 12878 40230 12930 40282
rect 12942 40230 12994 40282
rect 13006 40230 13058 40282
rect 13070 40230 13122 40282
rect 20808 40230 20860 40282
rect 20872 40230 20924 40282
rect 20936 40230 20988 40282
rect 21000 40230 21052 40282
rect 5264 40128 5316 40180
rect 9220 40128 9272 40180
rect 10416 40128 10468 40180
rect 12716 40128 12768 40180
rect 15384 40128 15436 40180
rect 3516 40035 3568 40044
rect 3516 40001 3525 40035
rect 3525 40001 3559 40035
rect 3559 40001 3568 40035
rect 3516 39992 3568 40001
rect 6368 39992 6420 40044
rect 11428 40060 11480 40112
rect 2504 39924 2556 39976
rect 4804 39967 4856 39976
rect 4804 39933 4813 39967
rect 4813 39933 4847 39967
rect 4847 39933 4856 39967
rect 4804 39924 4856 39933
rect 5356 39967 5408 39976
rect 5356 39933 5365 39967
rect 5365 39933 5399 39967
rect 5399 39933 5408 39967
rect 5356 39924 5408 39933
rect 7748 39856 7800 39908
rect 8760 39924 8812 39976
rect 9220 39967 9272 39976
rect 9220 39933 9229 39967
rect 9229 39933 9263 39967
rect 9263 39933 9272 39967
rect 9220 39924 9272 39933
rect 9864 39967 9916 39976
rect 9864 39933 9873 39967
rect 9873 39933 9907 39967
rect 9907 39933 9916 39967
rect 9864 39924 9916 39933
rect 10232 39856 10284 39908
rect 15200 39992 15252 40044
rect 10968 39967 11020 39976
rect 10968 39933 10977 39967
rect 10977 39933 11011 39967
rect 11011 39933 11020 39967
rect 10968 39924 11020 39933
rect 11428 39967 11480 39976
rect 11428 39933 11437 39967
rect 11437 39933 11471 39967
rect 11471 39933 11480 39967
rect 11428 39924 11480 39933
rect 11612 39924 11664 39976
rect 13544 39967 13596 39976
rect 13544 39933 13553 39967
rect 13553 39933 13587 39967
rect 13587 39933 13596 39967
rect 13820 39967 13872 39976
rect 13544 39924 13596 39933
rect 13820 39933 13829 39967
rect 13829 39933 13863 39967
rect 13863 39933 13872 39967
rect 13820 39924 13872 39933
rect 14924 39967 14976 39976
rect 14924 39933 14933 39967
rect 14933 39933 14967 39967
rect 14967 39933 14976 39967
rect 14924 39924 14976 39933
rect 16120 39967 16172 39976
rect 16120 39933 16129 39967
rect 16129 39933 16163 39967
rect 16163 39933 16172 39967
rect 16120 39924 16172 39933
rect 16304 39967 16356 39976
rect 16304 39933 16313 39967
rect 16313 39933 16347 39967
rect 16347 39933 16356 39967
rect 16304 39924 16356 39933
rect 18328 39924 18380 39976
rect 22100 39924 22152 39976
rect 15384 39856 15436 39908
rect 16488 39856 16540 39908
rect 16672 39856 16724 39908
rect 4252 39788 4304 39840
rect 5264 39788 5316 39840
rect 8912 39686 8964 39738
rect 8976 39686 9028 39738
rect 9040 39686 9092 39738
rect 9104 39686 9156 39738
rect 16843 39686 16895 39738
rect 16907 39686 16959 39738
rect 16971 39686 17023 39738
rect 17035 39686 17087 39738
rect 13820 39584 13872 39636
rect 18328 39627 18380 39636
rect 2688 39516 2740 39568
rect 4620 39491 4672 39500
rect 4620 39457 4629 39491
rect 4629 39457 4663 39491
rect 4663 39457 4672 39491
rect 4620 39448 4672 39457
rect 4712 39448 4764 39500
rect 5356 39448 5408 39500
rect 6828 39516 6880 39568
rect 18328 39593 18337 39627
rect 18337 39593 18371 39627
rect 18371 39593 18380 39627
rect 18328 39584 18380 39593
rect 7748 39491 7800 39500
rect 7748 39457 7757 39491
rect 7757 39457 7791 39491
rect 7791 39457 7800 39491
rect 7748 39448 7800 39457
rect 8392 39491 8444 39500
rect 6552 39380 6604 39432
rect 6368 39312 6420 39364
rect 8392 39457 8401 39491
rect 8401 39457 8435 39491
rect 8435 39457 8444 39491
rect 8392 39448 8444 39457
rect 8760 39491 8812 39500
rect 8760 39457 8769 39491
rect 8769 39457 8803 39491
rect 8803 39457 8812 39491
rect 8760 39448 8812 39457
rect 9864 39448 9916 39500
rect 10876 39448 10928 39500
rect 12440 39448 12492 39500
rect 13176 39491 13228 39500
rect 13176 39457 13185 39491
rect 13185 39457 13219 39491
rect 13219 39457 13228 39491
rect 13176 39448 13228 39457
rect 10784 39423 10836 39432
rect 10784 39389 10793 39423
rect 10793 39389 10827 39423
rect 10827 39389 10836 39423
rect 10784 39380 10836 39389
rect 8392 39312 8444 39364
rect 12624 39312 12676 39364
rect 14464 39448 14516 39500
rect 15200 39448 15252 39500
rect 15384 39448 15436 39500
rect 16672 39448 16724 39500
rect 15660 39380 15712 39432
rect 16580 39380 16632 39432
rect 14832 39312 14884 39364
rect 4528 39244 4580 39296
rect 7012 39244 7064 39296
rect 7840 39244 7892 39296
rect 14096 39244 14148 39296
rect 4947 39142 4999 39194
rect 5011 39142 5063 39194
rect 5075 39142 5127 39194
rect 5139 39142 5191 39194
rect 12878 39142 12930 39194
rect 12942 39142 12994 39194
rect 13006 39142 13058 39194
rect 13070 39142 13122 39194
rect 20808 39142 20860 39194
rect 20872 39142 20924 39194
rect 20936 39142 20988 39194
rect 21000 39142 21052 39194
rect 2504 39083 2556 39092
rect 2504 39049 2513 39083
rect 2513 39049 2547 39083
rect 2547 39049 2556 39083
rect 2504 39040 2556 39049
rect 3700 39083 3752 39092
rect 3700 39049 3709 39083
rect 3709 39049 3743 39083
rect 3743 39049 3752 39083
rect 3700 39040 3752 39049
rect 11612 39040 11664 39092
rect 9588 38972 9640 39024
rect 10048 38972 10100 39024
rect 12072 38972 12124 39024
rect 2412 38904 2464 38956
rect 3424 38836 3476 38888
rect 3700 38879 3752 38888
rect 3700 38845 3709 38879
rect 3709 38845 3743 38879
rect 3743 38845 3752 38879
rect 3700 38836 3752 38845
rect 4528 38904 4580 38956
rect 5356 38904 5408 38956
rect 5540 38947 5592 38956
rect 5540 38913 5549 38947
rect 5549 38913 5583 38947
rect 5583 38913 5592 38947
rect 5540 38904 5592 38913
rect 7472 38947 7524 38956
rect 7472 38913 7481 38947
rect 7481 38913 7515 38947
rect 7515 38913 7524 38947
rect 7472 38904 7524 38913
rect 10600 38904 10652 38956
rect 12624 38947 12676 38956
rect 12624 38913 12633 38947
rect 12633 38913 12667 38947
rect 12667 38913 12676 38947
rect 12624 38904 12676 38913
rect 16212 38904 16264 38956
rect 5908 38879 5960 38888
rect 3516 38768 3568 38820
rect 5908 38845 5917 38879
rect 5917 38845 5951 38879
rect 5951 38845 5960 38879
rect 5908 38836 5960 38845
rect 6828 38836 6880 38888
rect 7656 38879 7708 38888
rect 7656 38845 7665 38879
rect 7665 38845 7699 38879
rect 7699 38845 7708 38879
rect 7656 38836 7708 38845
rect 5816 38768 5868 38820
rect 5540 38700 5592 38752
rect 9864 38836 9916 38888
rect 11336 38879 11388 38888
rect 11336 38845 11337 38879
rect 11337 38845 11371 38879
rect 11371 38845 11388 38879
rect 11336 38836 11388 38845
rect 12716 38836 12768 38888
rect 15844 38879 15896 38888
rect 10600 38768 10652 38820
rect 15844 38845 15853 38879
rect 15853 38845 15887 38879
rect 15887 38845 15896 38879
rect 15844 38836 15896 38845
rect 16672 38879 16724 38888
rect 16672 38845 16681 38879
rect 16681 38845 16715 38879
rect 16715 38845 16724 38879
rect 16672 38836 16724 38845
rect 16396 38768 16448 38820
rect 8760 38700 8812 38752
rect 13820 38700 13872 38752
rect 16120 38700 16172 38752
rect 8912 38598 8964 38650
rect 8976 38598 9028 38650
rect 9040 38598 9092 38650
rect 9104 38598 9156 38650
rect 16843 38598 16895 38650
rect 16907 38598 16959 38650
rect 16971 38598 17023 38650
rect 17035 38598 17087 38650
rect 3516 38496 3568 38548
rect 7748 38496 7800 38548
rect 9864 38539 9916 38548
rect 9864 38505 9873 38539
rect 9873 38505 9907 38539
rect 9907 38505 9916 38539
rect 9864 38496 9916 38505
rect 1952 38428 2004 38480
rect 3608 38428 3660 38480
rect 4068 38403 4120 38412
rect 4068 38369 4077 38403
rect 4077 38369 4111 38403
rect 4111 38369 4120 38403
rect 4068 38360 4120 38369
rect 8760 38428 8812 38480
rect 6000 38360 6052 38412
rect 5908 38292 5960 38344
rect 6644 38360 6696 38412
rect 7564 38360 7616 38412
rect 7656 38403 7708 38412
rect 7656 38369 7665 38403
rect 7665 38369 7699 38403
rect 7699 38369 7708 38403
rect 7656 38360 7708 38369
rect 8668 38360 8720 38412
rect 10876 38360 10928 38412
rect 13820 38428 13872 38480
rect 11336 38360 11388 38412
rect 15752 38428 15804 38480
rect 16488 38428 16540 38480
rect 11244 38335 11296 38344
rect 11244 38301 11253 38335
rect 11253 38301 11287 38335
rect 11287 38301 11296 38335
rect 11244 38292 11296 38301
rect 14464 38360 14516 38412
rect 15568 38403 15620 38412
rect 15568 38369 15577 38403
rect 15577 38369 15611 38403
rect 15611 38369 15620 38403
rect 15568 38360 15620 38369
rect 15844 38403 15896 38412
rect 15844 38369 15853 38403
rect 15853 38369 15887 38403
rect 15887 38369 15896 38403
rect 15844 38360 15896 38369
rect 19984 38360 20036 38412
rect 14556 38292 14608 38344
rect 16304 38292 16356 38344
rect 5448 38224 5500 38276
rect 8760 38156 8812 38208
rect 10968 38156 11020 38208
rect 13176 38156 13228 38208
rect 16212 38156 16264 38208
rect 4947 38054 4999 38106
rect 5011 38054 5063 38106
rect 5075 38054 5127 38106
rect 5139 38054 5191 38106
rect 12878 38054 12930 38106
rect 12942 38054 12994 38106
rect 13006 38054 13058 38106
rect 13070 38054 13122 38106
rect 20808 38054 20860 38106
rect 20872 38054 20924 38106
rect 20936 38054 20988 38106
rect 21000 38054 21052 38106
rect 3424 37952 3476 38004
rect 6368 37952 6420 38004
rect 6736 37952 6788 38004
rect 10968 37995 11020 38004
rect 6276 37884 6328 37936
rect 10968 37961 10977 37995
rect 10977 37961 11011 37995
rect 11011 37961 11020 37995
rect 10968 37952 11020 37961
rect 11428 37995 11480 38004
rect 11428 37961 11437 37995
rect 11437 37961 11471 37995
rect 11471 37961 11480 37995
rect 11428 37952 11480 37961
rect 12716 37952 12768 38004
rect 12256 37884 12308 37936
rect 7840 37816 7892 37868
rect 10876 37816 10928 37868
rect 12072 37816 12124 37868
rect 13452 37859 13504 37868
rect 13452 37825 13461 37859
rect 13461 37825 13495 37859
rect 13495 37825 13504 37859
rect 13452 37816 13504 37825
rect 3884 37791 3936 37800
rect 3884 37757 3893 37791
rect 3893 37757 3927 37791
rect 3927 37757 3936 37791
rect 3884 37748 3936 37757
rect 4528 37791 4580 37800
rect 4528 37757 4537 37791
rect 4537 37757 4571 37791
rect 4571 37757 4580 37791
rect 4528 37748 4580 37757
rect 5540 37748 5592 37800
rect 6368 37748 6420 37800
rect 7656 37748 7708 37800
rect 8760 37791 8812 37800
rect 8760 37757 8769 37791
rect 8769 37757 8803 37791
rect 8803 37757 8812 37791
rect 8760 37748 8812 37757
rect 8024 37680 8076 37732
rect 11336 37748 11388 37800
rect 11612 37680 11664 37732
rect 13820 37748 13872 37800
rect 14096 37791 14148 37800
rect 14096 37757 14105 37791
rect 14105 37757 14139 37791
rect 14139 37757 14148 37791
rect 14096 37748 14148 37757
rect 15108 37748 15160 37800
rect 16028 37791 16080 37800
rect 15292 37680 15344 37732
rect 10048 37655 10100 37664
rect 10048 37621 10057 37655
rect 10057 37621 10091 37655
rect 10091 37621 10100 37655
rect 10048 37612 10100 37621
rect 11520 37612 11572 37664
rect 13176 37612 13228 37664
rect 15752 37612 15804 37664
rect 16028 37757 16037 37791
rect 16037 37757 16071 37791
rect 16071 37757 16080 37791
rect 16028 37748 16080 37757
rect 16304 37791 16356 37800
rect 16304 37757 16313 37791
rect 16313 37757 16347 37791
rect 16347 37757 16356 37791
rect 16304 37748 16356 37757
rect 16212 37723 16264 37732
rect 16212 37689 16221 37723
rect 16221 37689 16255 37723
rect 16255 37689 16264 37723
rect 16212 37680 16264 37689
rect 16672 37680 16724 37732
rect 8912 37510 8964 37562
rect 8976 37510 9028 37562
rect 9040 37510 9092 37562
rect 9104 37510 9156 37562
rect 16843 37510 16895 37562
rect 16907 37510 16959 37562
rect 16971 37510 17023 37562
rect 17035 37510 17087 37562
rect 5632 37408 5684 37460
rect 5724 37408 5776 37460
rect 8024 37408 8076 37460
rect 12072 37451 12124 37460
rect 2412 37315 2464 37324
rect 2412 37281 2421 37315
rect 2421 37281 2455 37315
rect 2455 37281 2464 37315
rect 2412 37272 2464 37281
rect 4160 37272 4212 37324
rect 4252 37204 4304 37256
rect 7104 37272 7156 37324
rect 7564 37315 7616 37324
rect 7564 37281 7573 37315
rect 7573 37281 7607 37315
rect 7607 37281 7616 37315
rect 7564 37272 7616 37281
rect 8024 37315 8076 37324
rect 5448 37204 5500 37256
rect 8024 37281 8033 37315
rect 8033 37281 8067 37315
rect 8067 37281 8076 37315
rect 8024 37272 8076 37281
rect 8760 37340 8812 37392
rect 10416 37340 10468 37392
rect 11244 37340 11296 37392
rect 10324 37272 10376 37324
rect 11520 37272 11572 37324
rect 12072 37417 12081 37451
rect 12081 37417 12115 37451
rect 12115 37417 12124 37451
rect 12072 37408 12124 37417
rect 14464 37408 14516 37460
rect 11704 37340 11756 37392
rect 14924 37340 14976 37392
rect 11244 37204 11296 37256
rect 13176 37315 13228 37324
rect 13176 37281 13185 37315
rect 13185 37281 13219 37315
rect 13219 37281 13228 37315
rect 13176 37272 13228 37281
rect 13820 37272 13872 37324
rect 15292 37315 15344 37324
rect 15292 37281 15301 37315
rect 15301 37281 15335 37315
rect 15335 37281 15344 37315
rect 15292 37272 15344 37281
rect 19984 37340 20036 37392
rect 16764 37315 16816 37324
rect 16764 37281 16773 37315
rect 16773 37281 16807 37315
rect 16807 37281 16816 37315
rect 16764 37272 16816 37281
rect 3056 37068 3108 37120
rect 8116 37068 8168 37120
rect 16028 37068 16080 37120
rect 4947 36966 4999 37018
rect 5011 36966 5063 37018
rect 5075 36966 5127 37018
rect 5139 36966 5191 37018
rect 12878 36966 12930 37018
rect 12942 36966 12994 37018
rect 13006 36966 13058 37018
rect 13070 36966 13122 37018
rect 20808 36966 20860 37018
rect 20872 36966 20924 37018
rect 20936 36966 20988 37018
rect 21000 36966 21052 37018
rect 4344 36907 4396 36916
rect 4344 36873 4353 36907
rect 4353 36873 4387 36907
rect 4387 36873 4396 36907
rect 4344 36864 4396 36873
rect 5632 36864 5684 36916
rect 7104 36907 7156 36916
rect 7104 36873 7113 36907
rect 7113 36873 7147 36907
rect 7147 36873 7156 36907
rect 7104 36864 7156 36873
rect 8116 36864 8168 36916
rect 10784 36907 10836 36916
rect 10784 36873 10793 36907
rect 10793 36873 10827 36907
rect 10827 36873 10836 36907
rect 10784 36864 10836 36873
rect 10968 36864 11020 36916
rect 15200 36864 15252 36916
rect 15936 36864 15988 36916
rect 16304 36864 16356 36916
rect 3056 36771 3108 36780
rect 3056 36737 3065 36771
rect 3065 36737 3099 36771
rect 3099 36737 3108 36771
rect 3056 36728 3108 36737
rect 4252 36728 4304 36780
rect 4068 36660 4120 36712
rect 5356 36660 5408 36712
rect 9680 36771 9732 36780
rect 9680 36737 9689 36771
rect 9689 36737 9723 36771
rect 9723 36737 9732 36771
rect 9680 36728 9732 36737
rect 6920 36703 6972 36712
rect 6920 36669 6929 36703
rect 6929 36669 6963 36703
rect 6963 36669 6972 36703
rect 6920 36660 6972 36669
rect 7932 36660 7984 36712
rect 9772 36703 9824 36712
rect 9772 36669 9781 36703
rect 9781 36669 9815 36703
rect 9815 36669 9824 36703
rect 9772 36660 9824 36669
rect 10324 36703 10376 36712
rect 10324 36669 10333 36703
rect 10333 36669 10367 36703
rect 10367 36669 10376 36703
rect 10324 36660 10376 36669
rect 11336 36660 11388 36712
rect 12440 36728 12492 36780
rect 14464 36728 14516 36780
rect 15108 36771 15160 36780
rect 15108 36737 15117 36771
rect 15117 36737 15151 36771
rect 15151 36737 15160 36771
rect 15108 36728 15160 36737
rect 13360 36660 13412 36712
rect 14648 36703 14700 36712
rect 14648 36669 14657 36703
rect 14657 36669 14691 36703
rect 14691 36669 14700 36703
rect 14648 36660 14700 36669
rect 14740 36703 14792 36712
rect 14740 36669 14749 36703
rect 14749 36669 14783 36703
rect 14783 36669 14792 36703
rect 15016 36703 15068 36712
rect 14740 36660 14792 36669
rect 15016 36669 15025 36703
rect 15025 36669 15059 36703
rect 15059 36669 15068 36703
rect 15016 36660 15068 36669
rect 15476 36660 15528 36712
rect 13636 36592 13688 36644
rect 15108 36592 15160 36644
rect 15752 36592 15804 36644
rect 3148 36524 3200 36576
rect 5540 36524 5592 36576
rect 8760 36524 8812 36576
rect 9772 36524 9824 36576
rect 10324 36524 10376 36576
rect 11612 36524 11664 36576
rect 13544 36524 13596 36576
rect 8912 36422 8964 36474
rect 8976 36422 9028 36474
rect 9040 36422 9092 36474
rect 9104 36422 9156 36474
rect 16843 36422 16895 36474
rect 16907 36422 16959 36474
rect 16971 36422 17023 36474
rect 17035 36422 17087 36474
rect 6460 36320 6512 36372
rect 10692 36320 10744 36372
rect 15384 36320 15436 36372
rect 3148 36252 3200 36304
rect 6920 36252 6972 36304
rect 5172 36227 5224 36236
rect 5172 36193 5181 36227
rect 5181 36193 5215 36227
rect 5215 36193 5224 36227
rect 5172 36184 5224 36193
rect 3240 35980 3292 36032
rect 5356 36184 5408 36236
rect 5724 36227 5776 36236
rect 5724 36193 5733 36227
rect 5733 36193 5767 36227
rect 5767 36193 5776 36227
rect 5724 36184 5776 36193
rect 6460 36184 6512 36236
rect 11244 36252 11296 36304
rect 11520 36252 11572 36304
rect 13820 36252 13872 36304
rect 11428 36184 11480 36236
rect 13360 36227 13412 36236
rect 13360 36193 13369 36227
rect 13369 36193 13403 36227
rect 13403 36193 13412 36227
rect 13360 36184 13412 36193
rect 13636 36184 13688 36236
rect 14096 36184 14148 36236
rect 15016 36184 15068 36236
rect 15936 36184 15988 36236
rect 5540 36116 5592 36168
rect 7380 36159 7432 36168
rect 7380 36125 7389 36159
rect 7389 36125 7423 36159
rect 7423 36125 7432 36159
rect 7380 36116 7432 36125
rect 8668 36116 8720 36168
rect 13452 36116 13504 36168
rect 14740 36116 14792 36168
rect 11336 36048 11388 36100
rect 15292 36048 15344 36100
rect 8852 35980 8904 36032
rect 12716 35980 12768 36032
rect 17132 36023 17184 36032
rect 17132 35989 17141 36023
rect 17141 35989 17175 36023
rect 17175 35989 17184 36023
rect 17132 35980 17184 35989
rect 4947 35878 4999 35930
rect 5011 35878 5063 35930
rect 5075 35878 5127 35930
rect 5139 35878 5191 35930
rect 12878 35878 12930 35930
rect 12942 35878 12994 35930
rect 13006 35878 13058 35930
rect 13070 35878 13122 35930
rect 20808 35878 20860 35930
rect 20872 35878 20924 35930
rect 20936 35878 20988 35930
rect 21000 35878 21052 35930
rect 2044 35640 2096 35692
rect 2688 35640 2740 35692
rect 8852 35776 8904 35828
rect 11428 35776 11480 35828
rect 11704 35776 11756 35828
rect 7380 35708 7432 35760
rect 12716 35683 12768 35692
rect 4436 35572 4488 35624
rect 4712 35615 4764 35624
rect 4712 35581 4721 35615
rect 4721 35581 4755 35615
rect 4755 35581 4764 35615
rect 4712 35572 4764 35581
rect 2688 35504 2740 35556
rect 4712 35436 4764 35488
rect 5632 35572 5684 35624
rect 12716 35649 12725 35683
rect 12725 35649 12759 35683
rect 12759 35649 12768 35683
rect 12716 35640 12768 35649
rect 12808 35640 12860 35692
rect 8668 35615 8720 35624
rect 6092 35504 6144 35556
rect 7012 35479 7064 35488
rect 7012 35445 7021 35479
rect 7021 35445 7055 35479
rect 7055 35445 7064 35479
rect 7012 35436 7064 35445
rect 8668 35581 8677 35615
rect 8677 35581 8711 35615
rect 8711 35581 8720 35615
rect 8668 35572 8720 35581
rect 8484 35504 8536 35556
rect 10968 35572 11020 35624
rect 11888 35572 11940 35624
rect 8852 35504 8904 35556
rect 11612 35504 11664 35556
rect 9680 35436 9732 35488
rect 11428 35479 11480 35488
rect 11428 35445 11437 35479
rect 11437 35445 11471 35479
rect 11471 35445 11480 35479
rect 11428 35436 11480 35445
rect 15108 35776 15160 35828
rect 15200 35683 15252 35692
rect 15200 35649 15209 35683
rect 15209 35649 15243 35683
rect 15243 35649 15252 35683
rect 15200 35640 15252 35649
rect 14924 35615 14976 35624
rect 14924 35581 14933 35615
rect 14933 35581 14967 35615
rect 14967 35581 14976 35615
rect 14924 35572 14976 35581
rect 18420 35572 18472 35624
rect 19616 35504 19668 35556
rect 14924 35436 14976 35488
rect 16580 35436 16632 35488
rect 8912 35334 8964 35386
rect 8976 35334 9028 35386
rect 9040 35334 9092 35386
rect 9104 35334 9156 35386
rect 16843 35334 16895 35386
rect 16907 35334 16959 35386
rect 16971 35334 17023 35386
rect 17035 35334 17087 35386
rect 4252 35139 4304 35148
rect 4252 35105 4261 35139
rect 4261 35105 4295 35139
rect 4295 35105 4304 35139
rect 4252 35096 4304 35105
rect 5356 35232 5408 35284
rect 7012 35232 7064 35284
rect 11704 35232 11756 35284
rect 11980 35232 12032 35284
rect 8116 35164 8168 35216
rect 5724 35096 5776 35148
rect 14648 35232 14700 35284
rect 14464 35164 14516 35216
rect 21364 35164 21416 35216
rect 2044 35028 2096 35080
rect 4160 34935 4212 34944
rect 4160 34901 4169 34935
rect 4169 34901 4203 34935
rect 4203 34901 4212 34935
rect 4160 34892 4212 34901
rect 7288 35028 7340 35080
rect 10232 35071 10284 35080
rect 10232 35037 10241 35071
rect 10241 35037 10275 35071
rect 10275 35037 10284 35071
rect 10232 35028 10284 35037
rect 12532 35139 12584 35148
rect 12532 35105 12547 35139
rect 12547 35105 12581 35139
rect 12581 35105 12584 35139
rect 13636 35139 13688 35148
rect 12532 35096 12584 35105
rect 13636 35105 13645 35139
rect 13645 35105 13679 35139
rect 13679 35105 13688 35139
rect 13636 35096 13688 35105
rect 16672 35096 16724 35148
rect 17132 35096 17184 35148
rect 13820 35028 13872 35080
rect 14464 35028 14516 35080
rect 14740 35028 14792 35080
rect 11888 34960 11940 35012
rect 11336 34892 11388 34944
rect 11980 34892 12032 34944
rect 12532 34960 12584 35012
rect 15292 34960 15344 35012
rect 13360 34892 13412 34944
rect 13820 34935 13872 34944
rect 13820 34901 13844 34935
rect 13844 34901 13872 34935
rect 13820 34892 13872 34901
rect 18512 35028 18564 35080
rect 17224 34892 17276 34944
rect 4947 34790 4999 34842
rect 5011 34790 5063 34842
rect 5075 34790 5127 34842
rect 5139 34790 5191 34842
rect 12878 34790 12930 34842
rect 12942 34790 12994 34842
rect 13006 34790 13058 34842
rect 13070 34790 13122 34842
rect 20808 34790 20860 34842
rect 20872 34790 20924 34842
rect 20936 34790 20988 34842
rect 21000 34790 21052 34842
rect 4344 34688 4396 34740
rect 6460 34688 6512 34740
rect 6828 34688 6880 34740
rect 2596 34484 2648 34536
rect 5632 34620 5684 34672
rect 3056 34552 3108 34604
rect 2964 34348 3016 34400
rect 4068 34484 4120 34536
rect 4528 34527 4580 34536
rect 4528 34493 4537 34527
rect 4537 34493 4571 34527
rect 4571 34493 4580 34527
rect 4528 34484 4580 34493
rect 4712 34527 4764 34536
rect 4712 34493 4721 34527
rect 4721 34493 4755 34527
rect 4755 34493 4764 34527
rect 4712 34484 4764 34493
rect 6460 34552 6512 34604
rect 9312 34688 9364 34740
rect 10232 34731 10284 34740
rect 10232 34697 10241 34731
rect 10241 34697 10275 34731
rect 10275 34697 10284 34731
rect 10232 34688 10284 34697
rect 11428 34688 11480 34740
rect 13176 34688 13228 34740
rect 16028 34688 16080 34740
rect 18512 34731 18564 34740
rect 18512 34697 18521 34731
rect 18521 34697 18555 34731
rect 18555 34697 18564 34731
rect 18512 34688 18564 34697
rect 5264 34527 5316 34536
rect 5264 34493 5273 34527
rect 5273 34493 5307 34527
rect 5307 34493 5316 34527
rect 8300 34620 8352 34672
rect 5264 34484 5316 34493
rect 7472 34527 7524 34536
rect 7472 34493 7481 34527
rect 7481 34493 7515 34527
rect 7515 34493 7524 34527
rect 7472 34484 7524 34493
rect 7564 34527 7616 34536
rect 7564 34493 7573 34527
rect 7573 34493 7607 34527
rect 7607 34493 7616 34527
rect 7564 34484 7616 34493
rect 8484 34484 8536 34536
rect 9864 34620 9916 34672
rect 12808 34595 12860 34604
rect 12808 34561 12817 34595
rect 12817 34561 12851 34595
rect 12851 34561 12860 34595
rect 12808 34552 12860 34561
rect 9312 34527 9364 34536
rect 9312 34493 9321 34527
rect 9321 34493 9355 34527
rect 9355 34493 9364 34527
rect 9312 34484 9364 34493
rect 9772 34527 9824 34536
rect 9772 34493 9781 34527
rect 9781 34493 9815 34527
rect 9815 34493 9824 34527
rect 9772 34484 9824 34493
rect 9956 34484 10008 34536
rect 11336 34527 11388 34536
rect 11336 34493 11345 34527
rect 11345 34493 11379 34527
rect 11379 34493 11388 34527
rect 11336 34484 11388 34493
rect 10140 34416 10192 34468
rect 12624 34484 12676 34536
rect 16304 34552 16356 34604
rect 16396 34552 16448 34604
rect 14004 34527 14056 34536
rect 14004 34493 14013 34527
rect 14013 34493 14047 34527
rect 14047 34493 14056 34527
rect 14004 34484 14056 34493
rect 15660 34484 15712 34536
rect 15752 34527 15804 34536
rect 15752 34493 15761 34527
rect 15761 34493 15795 34527
rect 15795 34493 15804 34527
rect 15752 34484 15804 34493
rect 21364 34484 21416 34536
rect 19616 34459 19668 34468
rect 5540 34348 5592 34400
rect 7748 34348 7800 34400
rect 19616 34425 19625 34459
rect 19625 34425 19659 34459
rect 19659 34425 19668 34459
rect 19616 34416 19668 34425
rect 8912 34246 8964 34298
rect 8976 34246 9028 34298
rect 9040 34246 9092 34298
rect 9104 34246 9156 34298
rect 16843 34246 16895 34298
rect 16907 34246 16959 34298
rect 16971 34246 17023 34298
rect 17035 34246 17087 34298
rect 3700 34144 3752 34196
rect 7472 34144 7524 34196
rect 8484 34187 8536 34196
rect 8484 34153 8493 34187
rect 8493 34153 8527 34187
rect 8527 34153 8536 34187
rect 8484 34144 8536 34153
rect 9956 34187 10008 34196
rect 9956 34153 9965 34187
rect 9965 34153 9999 34187
rect 9999 34153 10008 34187
rect 9956 34144 10008 34153
rect 11060 34187 11112 34196
rect 11060 34153 11069 34187
rect 11069 34153 11103 34187
rect 11103 34153 11112 34187
rect 11060 34144 11112 34153
rect 12440 34144 12492 34196
rect 11428 34076 11480 34128
rect 2596 34051 2648 34060
rect 2596 34017 2605 34051
rect 2605 34017 2639 34051
rect 2639 34017 2648 34051
rect 2596 34008 2648 34017
rect 2964 34051 3016 34060
rect 2964 34017 2973 34051
rect 2973 34017 3007 34051
rect 3007 34017 3016 34051
rect 2964 34008 3016 34017
rect 3148 34051 3200 34060
rect 3148 34017 3157 34051
rect 3157 34017 3191 34051
rect 3191 34017 3200 34051
rect 3148 34008 3200 34017
rect 5908 34008 5960 34060
rect 6092 34051 6144 34060
rect 6092 34017 6101 34051
rect 6101 34017 6135 34051
rect 6135 34017 6144 34051
rect 6092 34008 6144 34017
rect 8300 34051 8352 34060
rect 8300 34017 8309 34051
rect 8309 34017 8343 34051
rect 8343 34017 8352 34051
rect 8300 34008 8352 34017
rect 9864 34008 9916 34060
rect 10416 34008 10468 34060
rect 11244 34008 11296 34060
rect 18420 34076 18472 34128
rect 2688 33983 2740 33992
rect 2688 33949 2697 33983
rect 2697 33949 2731 33983
rect 2731 33949 2740 33983
rect 2688 33940 2740 33949
rect 5724 33940 5776 33992
rect 10600 33940 10652 33992
rect 10048 33872 10100 33924
rect 11060 33872 11112 33924
rect 12440 34008 12492 34060
rect 12808 34008 12860 34060
rect 11888 33940 11940 33992
rect 12164 33872 12216 33924
rect 15752 34008 15804 34060
rect 16396 33940 16448 33992
rect 14740 33872 14792 33924
rect 15292 33872 15344 33924
rect 17224 34008 17276 34060
rect 16764 33940 16816 33992
rect 1952 33804 2004 33856
rect 7196 33847 7248 33856
rect 7196 33813 7205 33847
rect 7205 33813 7239 33847
rect 7239 33813 7248 33847
rect 7196 33804 7248 33813
rect 4947 33702 4999 33754
rect 5011 33702 5063 33754
rect 5075 33702 5127 33754
rect 5139 33702 5191 33754
rect 12878 33702 12930 33754
rect 12942 33702 12994 33754
rect 13006 33702 13058 33754
rect 13070 33702 13122 33754
rect 20808 33702 20860 33754
rect 20872 33702 20924 33754
rect 20936 33702 20988 33754
rect 21000 33702 21052 33754
rect 5908 33600 5960 33652
rect 14004 33643 14056 33652
rect 1492 33464 1544 33516
rect 5724 33532 5776 33584
rect 14004 33609 14013 33643
rect 14013 33609 14047 33643
rect 14047 33609 14056 33643
rect 14004 33600 14056 33609
rect 16028 33643 16080 33652
rect 16028 33609 16037 33643
rect 16037 33609 16071 33643
rect 16071 33609 16080 33643
rect 16028 33600 16080 33609
rect 11520 33532 11572 33584
rect 4620 33464 4672 33516
rect 3976 33396 4028 33448
rect 4160 33396 4212 33448
rect 7748 33507 7800 33516
rect 7748 33473 7757 33507
rect 7757 33473 7791 33507
rect 7791 33473 7800 33507
rect 7748 33464 7800 33473
rect 16764 33507 16816 33516
rect 16764 33473 16773 33507
rect 16773 33473 16807 33507
rect 16807 33473 16816 33507
rect 16764 33464 16816 33473
rect 5540 33396 5592 33448
rect 5632 33328 5684 33380
rect 3700 33260 3752 33312
rect 5356 33260 5408 33312
rect 5540 33260 5592 33312
rect 6184 33396 6236 33448
rect 10048 33396 10100 33448
rect 10232 33439 10284 33448
rect 10232 33405 10241 33439
rect 10241 33405 10275 33439
rect 10275 33405 10284 33439
rect 10600 33439 10652 33448
rect 10232 33396 10284 33405
rect 10600 33405 10609 33439
rect 10609 33405 10643 33439
rect 10643 33405 10652 33439
rect 10600 33396 10652 33405
rect 12532 33396 12584 33448
rect 12716 33439 12768 33448
rect 12716 33405 12725 33439
rect 12725 33405 12759 33439
rect 12759 33405 12768 33439
rect 12716 33396 12768 33405
rect 14924 33439 14976 33448
rect 14924 33405 14933 33439
rect 14933 33405 14967 33439
rect 14967 33405 14976 33439
rect 14924 33396 14976 33405
rect 16304 33439 16356 33448
rect 16304 33405 16313 33439
rect 16313 33405 16347 33439
rect 16347 33405 16356 33439
rect 16304 33396 16356 33405
rect 16580 33328 16632 33380
rect 5908 33260 5960 33312
rect 8760 33260 8812 33312
rect 9680 33260 9732 33312
rect 15016 33303 15068 33312
rect 15016 33269 15025 33303
rect 15025 33269 15059 33303
rect 15059 33269 15068 33303
rect 15016 33260 15068 33269
rect 8912 33158 8964 33210
rect 8976 33158 9028 33210
rect 9040 33158 9092 33210
rect 9104 33158 9156 33210
rect 16843 33158 16895 33210
rect 16907 33158 16959 33210
rect 16971 33158 17023 33210
rect 17035 33158 17087 33210
rect 2688 33056 2740 33108
rect 3056 33099 3108 33108
rect 3056 33065 3065 33099
rect 3065 33065 3099 33099
rect 3099 33065 3108 33099
rect 3056 33056 3108 33065
rect 4068 33056 4120 33108
rect 7380 33099 7432 33108
rect 7380 33065 7389 33099
rect 7389 33065 7423 33099
rect 7423 33065 7432 33099
rect 7380 33056 7432 33065
rect 10600 33056 10652 33108
rect 12716 33056 12768 33108
rect 1952 32963 2004 32972
rect 1952 32929 1961 32963
rect 1961 32929 1995 32963
rect 1995 32929 2004 32963
rect 1952 32920 2004 32929
rect 15200 32988 15252 33040
rect 3700 32920 3752 32972
rect 5908 32963 5960 32972
rect 5908 32929 5917 32963
rect 5917 32929 5951 32963
rect 5951 32929 5960 32963
rect 5908 32920 5960 32929
rect 4528 32852 4580 32904
rect 4712 32852 4764 32904
rect 6184 32852 6236 32904
rect 6460 32852 6512 32904
rect 9772 32920 9824 32972
rect 9956 32852 10008 32904
rect 10232 32920 10284 32972
rect 10692 32920 10744 32972
rect 11336 32963 11388 32972
rect 11336 32929 11345 32963
rect 11345 32929 11379 32963
rect 11379 32929 11388 32963
rect 11336 32920 11388 32929
rect 12440 32920 12492 32972
rect 13544 32963 13596 32972
rect 13544 32929 13553 32963
rect 13553 32929 13587 32963
rect 13587 32929 13596 32963
rect 13544 32920 13596 32929
rect 10968 32852 11020 32904
rect 14188 32920 14240 32972
rect 15016 32920 15068 32972
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 13912 32827 13964 32836
rect 13912 32793 13921 32827
rect 13921 32793 13955 32827
rect 13955 32793 13964 32827
rect 13912 32784 13964 32793
rect 15384 32852 15436 32904
rect 15844 32895 15896 32904
rect 15844 32861 15853 32895
rect 15853 32861 15887 32895
rect 15887 32861 15896 32895
rect 15844 32852 15896 32861
rect 16672 32920 16724 32972
rect 16580 32852 16632 32904
rect 5724 32759 5776 32768
rect 5724 32725 5733 32759
rect 5733 32725 5767 32759
rect 5767 32725 5776 32759
rect 5724 32716 5776 32725
rect 9864 32716 9916 32768
rect 13360 32759 13412 32768
rect 13360 32725 13369 32759
rect 13369 32725 13403 32759
rect 13403 32725 13412 32759
rect 13360 32716 13412 32725
rect 13820 32759 13872 32768
rect 13820 32725 13844 32759
rect 13844 32725 13872 32759
rect 15384 32759 15436 32768
rect 13820 32716 13872 32725
rect 15384 32725 15393 32759
rect 15393 32725 15427 32759
rect 15427 32725 15436 32759
rect 15384 32716 15436 32725
rect 4947 32614 4999 32666
rect 5011 32614 5063 32666
rect 5075 32614 5127 32666
rect 5139 32614 5191 32666
rect 12878 32614 12930 32666
rect 12942 32614 12994 32666
rect 13006 32614 13058 32666
rect 13070 32614 13122 32666
rect 20808 32614 20860 32666
rect 20872 32614 20924 32666
rect 20936 32614 20988 32666
rect 21000 32614 21052 32666
rect 14096 32512 14148 32564
rect 3976 32487 4028 32496
rect 3976 32453 3985 32487
rect 3985 32453 4019 32487
rect 4019 32453 4028 32487
rect 3976 32444 4028 32453
rect 5816 32444 5868 32496
rect 7472 32376 7524 32428
rect 8024 32376 8076 32428
rect 9680 32376 9732 32428
rect 9956 32376 10008 32428
rect 10324 32376 10376 32428
rect 12532 32376 12584 32428
rect 13544 32376 13596 32428
rect 15384 32376 15436 32428
rect 3056 32351 3108 32360
rect 1584 32215 1636 32224
rect 1584 32181 1593 32215
rect 1593 32181 1627 32215
rect 1627 32181 1636 32215
rect 1584 32172 1636 32181
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 3792 32351 3844 32360
rect 3792 32317 3801 32351
rect 3801 32317 3835 32351
rect 3835 32317 3844 32351
rect 3792 32308 3844 32317
rect 4068 32308 4120 32360
rect 4804 32308 4856 32360
rect 5724 32308 5776 32360
rect 6460 32308 6512 32360
rect 7104 32240 7156 32292
rect 8116 32308 8168 32360
rect 10140 32308 10192 32360
rect 10416 32308 10468 32360
rect 16304 32351 16356 32360
rect 16304 32317 16313 32351
rect 16313 32317 16347 32351
rect 16347 32317 16356 32351
rect 16304 32308 16356 32317
rect 7932 32240 7984 32292
rect 4712 32172 4764 32224
rect 5264 32215 5316 32224
rect 5264 32181 5273 32215
rect 5273 32181 5307 32215
rect 5307 32181 5316 32215
rect 5264 32172 5316 32181
rect 9220 32172 9272 32224
rect 16212 32240 16264 32292
rect 16488 32240 16540 32292
rect 10600 32172 10652 32224
rect 11704 32172 11756 32224
rect 14188 32172 14240 32224
rect 16580 32172 16632 32224
rect 8912 32070 8964 32122
rect 8976 32070 9028 32122
rect 9040 32070 9092 32122
rect 9104 32070 9156 32122
rect 16843 32070 16895 32122
rect 16907 32070 16959 32122
rect 16971 32070 17023 32122
rect 17035 32070 17087 32122
rect 5724 31968 5776 32020
rect 2780 31900 2832 31952
rect 7932 31968 7984 32020
rect 10048 31968 10100 32020
rect 10968 31968 11020 32020
rect 15292 31968 15344 32020
rect 16028 31968 16080 32020
rect 16304 31968 16356 32020
rect 2964 31875 3016 31884
rect 2964 31841 2973 31875
rect 2973 31841 3007 31875
rect 3007 31841 3016 31875
rect 4804 31875 4856 31884
rect 2964 31832 3016 31841
rect 4804 31841 4813 31875
rect 4813 31841 4847 31875
rect 4847 31841 4856 31875
rect 4804 31832 4856 31841
rect 7380 31900 7432 31952
rect 5816 31832 5868 31884
rect 6276 31832 6328 31884
rect 8300 31832 8352 31884
rect 13452 31900 13504 31952
rect 11336 31875 11388 31884
rect 6184 31807 6236 31816
rect 6184 31773 6193 31807
rect 6193 31773 6227 31807
rect 6227 31773 6236 31807
rect 6184 31764 6236 31773
rect 11336 31841 11345 31875
rect 11345 31841 11379 31875
rect 11379 31841 11388 31875
rect 11336 31832 11388 31841
rect 11704 31832 11756 31884
rect 12072 31875 12124 31884
rect 12072 31841 12081 31875
rect 12081 31841 12115 31875
rect 12115 31841 12124 31875
rect 12072 31832 12124 31841
rect 12532 31832 12584 31884
rect 13360 31832 13412 31884
rect 13636 31875 13688 31884
rect 13636 31841 13645 31875
rect 13645 31841 13679 31875
rect 13679 31841 13688 31875
rect 13636 31832 13688 31841
rect 14924 31832 14976 31884
rect 16212 31832 16264 31884
rect 16304 31832 16356 31884
rect 16488 31832 16540 31884
rect 4528 31696 4580 31748
rect 5448 31696 5500 31748
rect 8760 31764 8812 31816
rect 9496 31696 9548 31748
rect 10324 31764 10376 31816
rect 11060 31696 11112 31748
rect 14188 31764 14240 31816
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 15568 31807 15620 31816
rect 15568 31773 15577 31807
rect 15577 31773 15611 31807
rect 15611 31773 15620 31807
rect 15568 31764 15620 31773
rect 13820 31739 13872 31748
rect 13820 31705 13844 31739
rect 13844 31705 13872 31739
rect 13820 31696 13872 31705
rect 13912 31739 13964 31748
rect 13912 31705 13921 31739
rect 13921 31705 13955 31739
rect 13955 31705 13964 31739
rect 13912 31696 13964 31705
rect 5356 31628 5408 31680
rect 5816 31628 5868 31680
rect 8024 31628 8076 31680
rect 10232 31628 10284 31680
rect 12348 31671 12400 31680
rect 12348 31637 12357 31671
rect 12357 31637 12391 31671
rect 12391 31637 12400 31671
rect 12348 31628 12400 31637
rect 17868 31671 17920 31680
rect 17868 31637 17877 31671
rect 17877 31637 17911 31671
rect 17911 31637 17920 31671
rect 17868 31628 17920 31637
rect 4947 31526 4999 31578
rect 5011 31526 5063 31578
rect 5075 31526 5127 31578
rect 5139 31526 5191 31578
rect 12878 31526 12930 31578
rect 12942 31526 12994 31578
rect 13006 31526 13058 31578
rect 13070 31526 13122 31578
rect 20808 31526 20860 31578
rect 20872 31526 20924 31578
rect 20936 31526 20988 31578
rect 21000 31526 21052 31578
rect 4436 31424 4488 31476
rect 9680 31424 9732 31476
rect 10416 31424 10468 31476
rect 1492 31331 1544 31340
rect 1492 31297 1501 31331
rect 1501 31297 1535 31331
rect 1535 31297 1544 31331
rect 1492 31288 1544 31297
rect 5172 31356 5224 31408
rect 1768 31084 1820 31136
rect 3056 31220 3108 31272
rect 4896 31263 4948 31272
rect 4896 31229 4905 31263
rect 4905 31229 4939 31263
rect 4939 31229 4948 31263
rect 4896 31220 4948 31229
rect 9772 31288 9824 31340
rect 10324 31288 10376 31340
rect 8024 31220 8076 31272
rect 10416 31220 10468 31272
rect 10600 31263 10652 31272
rect 10600 31229 10609 31263
rect 10609 31229 10643 31263
rect 10643 31229 10652 31263
rect 10600 31220 10652 31229
rect 9220 31152 9272 31204
rect 9404 31084 9456 31136
rect 13544 31424 13596 31476
rect 14188 31424 14240 31476
rect 15568 31424 15620 31476
rect 12348 31288 12400 31340
rect 12440 31263 12492 31272
rect 12440 31229 12449 31263
rect 12449 31229 12483 31263
rect 12483 31229 12492 31263
rect 17868 31356 17920 31408
rect 16212 31331 16264 31340
rect 16212 31297 16221 31331
rect 16221 31297 16255 31331
rect 16255 31297 16264 31331
rect 16212 31288 16264 31297
rect 12440 31220 12492 31229
rect 15844 31263 15896 31272
rect 15844 31229 15853 31263
rect 15853 31229 15887 31263
rect 15887 31229 15896 31263
rect 15844 31220 15896 31229
rect 12532 31152 12584 31204
rect 15384 31152 15436 31204
rect 16028 31152 16080 31204
rect 13912 31084 13964 31136
rect 8912 30982 8964 31034
rect 8976 30982 9028 31034
rect 9040 30982 9092 31034
rect 9104 30982 9156 31034
rect 16843 30982 16895 31034
rect 16907 30982 16959 31034
rect 16971 30982 17023 31034
rect 17035 30982 17087 31034
rect 3056 30923 3108 30932
rect 3056 30889 3065 30923
rect 3065 30889 3099 30923
rect 3099 30889 3108 30923
rect 3056 30880 3108 30889
rect 3608 30880 3660 30932
rect 4804 30880 4856 30932
rect 6184 30923 6236 30932
rect 6184 30889 6193 30923
rect 6193 30889 6227 30923
rect 6227 30889 6236 30923
rect 6184 30880 6236 30889
rect 5816 30812 5868 30864
rect 7196 30812 7248 30864
rect 2964 30744 3016 30796
rect 5264 30744 5316 30796
rect 5356 30744 5408 30796
rect 5724 30787 5776 30796
rect 5724 30753 5733 30787
rect 5733 30753 5767 30787
rect 5767 30753 5776 30787
rect 5724 30744 5776 30753
rect 4436 30676 4488 30728
rect 6460 30744 6512 30796
rect 10324 30880 10376 30932
rect 10416 30880 10468 30932
rect 11428 30880 11480 30932
rect 9404 30812 9456 30864
rect 9956 30787 10008 30796
rect 9956 30753 9965 30787
rect 9965 30753 9999 30787
rect 9999 30753 10008 30787
rect 9956 30744 10008 30753
rect 10324 30744 10376 30796
rect 11796 30812 11848 30864
rect 12164 30812 12216 30864
rect 14464 30880 14516 30932
rect 14648 30880 14700 30932
rect 15200 30880 15252 30932
rect 14004 30787 14056 30796
rect 7012 30676 7064 30728
rect 12072 30676 12124 30728
rect 14004 30753 14013 30787
rect 14013 30753 14047 30787
rect 14047 30753 14056 30787
rect 14004 30744 14056 30753
rect 16580 30744 16632 30796
rect 16028 30676 16080 30728
rect 3976 30608 4028 30660
rect 5356 30608 5408 30660
rect 5908 30608 5960 30660
rect 7196 30583 7248 30592
rect 7196 30549 7205 30583
rect 7205 30549 7239 30583
rect 7239 30549 7248 30583
rect 8024 30608 8076 30660
rect 9956 30608 10008 30660
rect 11060 30608 11112 30660
rect 11520 30608 11572 30660
rect 13452 30608 13504 30660
rect 15292 30608 15344 30660
rect 7196 30540 7248 30549
rect 7840 30540 7892 30592
rect 14096 30583 14148 30592
rect 14096 30549 14105 30583
rect 14105 30549 14139 30583
rect 14139 30549 14148 30583
rect 14096 30540 14148 30549
rect 15384 30540 15436 30592
rect 16488 30540 16540 30592
rect 4947 30438 4999 30490
rect 5011 30438 5063 30490
rect 5075 30438 5127 30490
rect 5139 30438 5191 30490
rect 12878 30438 12930 30490
rect 12942 30438 12994 30490
rect 13006 30438 13058 30490
rect 13070 30438 13122 30490
rect 20808 30438 20860 30490
rect 20872 30438 20924 30490
rect 20936 30438 20988 30490
rect 21000 30438 21052 30490
rect 3516 30336 3568 30388
rect 5540 30336 5592 30388
rect 2872 30268 2924 30320
rect 2504 30132 2556 30184
rect 3056 30132 3108 30184
rect 3516 30132 3568 30184
rect 4068 30132 4120 30184
rect 4160 30132 4212 30184
rect 11152 30268 11204 30320
rect 11796 30268 11848 30320
rect 4344 30064 4396 30116
rect 5724 30064 5776 30116
rect 5908 30107 5960 30116
rect 5908 30073 5917 30107
rect 5917 30073 5951 30107
rect 5951 30073 5960 30107
rect 5908 30064 5960 30073
rect 6460 30132 6512 30184
rect 8024 30175 8076 30184
rect 8024 30141 8033 30175
rect 8033 30141 8067 30175
rect 8067 30141 8076 30175
rect 8024 30132 8076 30141
rect 8760 30200 8812 30252
rect 12624 30243 12676 30252
rect 12624 30209 12633 30243
rect 12633 30209 12667 30243
rect 12667 30209 12676 30243
rect 12624 30200 12676 30209
rect 9220 30132 9272 30184
rect 7380 30064 7432 30116
rect 8668 30107 8720 30116
rect 8668 30073 8677 30107
rect 8677 30073 8711 30107
rect 8711 30073 8720 30107
rect 8668 30064 8720 30073
rect 4160 30039 4212 30048
rect 4160 30005 4169 30039
rect 4169 30005 4203 30039
rect 4203 30005 4212 30039
rect 4160 29996 4212 30005
rect 6920 30039 6972 30048
rect 6920 30005 6929 30039
rect 6929 30005 6963 30039
rect 6963 30005 6972 30039
rect 6920 29996 6972 30005
rect 11428 30132 11480 30184
rect 12164 30132 12216 30184
rect 13176 30132 13228 30184
rect 14004 30268 14056 30320
rect 13636 30200 13688 30252
rect 15844 30243 15896 30252
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 16212 30200 16264 30252
rect 15936 30175 15988 30184
rect 15936 30141 15945 30175
rect 15945 30141 15979 30175
rect 15979 30141 15988 30175
rect 15936 30132 15988 30141
rect 16488 30132 16540 30184
rect 12072 30064 12124 30116
rect 15568 30064 15620 30116
rect 11060 29996 11112 30048
rect 17592 29996 17644 30048
rect 8912 29894 8964 29946
rect 8976 29894 9028 29946
rect 9040 29894 9092 29946
rect 9104 29894 9156 29946
rect 16843 29894 16895 29946
rect 16907 29894 16959 29946
rect 16971 29894 17023 29946
rect 17035 29894 17087 29946
rect 3516 29792 3568 29844
rect 4436 29792 4488 29844
rect 5356 29792 5408 29844
rect 5724 29792 5776 29844
rect 3148 29724 3200 29776
rect 3424 29724 3476 29776
rect 8024 29724 8076 29776
rect 11520 29792 11572 29844
rect 9864 29767 9916 29776
rect 1492 29656 1544 29708
rect 4160 29656 4212 29708
rect 3424 29588 3476 29640
rect 3608 29588 3660 29640
rect 2504 29452 2556 29504
rect 7196 29656 7248 29708
rect 9404 29656 9456 29708
rect 9864 29733 9873 29767
rect 9873 29733 9907 29767
rect 9907 29733 9916 29767
rect 9864 29724 9916 29733
rect 11704 29699 11756 29708
rect 8024 29588 8076 29640
rect 11704 29665 11713 29699
rect 11713 29665 11747 29699
rect 11747 29665 11756 29699
rect 11704 29656 11756 29665
rect 12164 29699 12216 29708
rect 12164 29665 12173 29699
rect 12173 29665 12207 29699
rect 12207 29665 12216 29699
rect 12164 29656 12216 29665
rect 12624 29656 12676 29708
rect 13728 29699 13780 29708
rect 13728 29665 13737 29699
rect 13737 29665 13771 29699
rect 13771 29665 13780 29699
rect 13728 29656 13780 29665
rect 13912 29699 13964 29708
rect 13912 29665 13921 29699
rect 13921 29665 13955 29699
rect 13955 29665 13964 29699
rect 13912 29656 13964 29665
rect 15200 29656 15252 29708
rect 15568 29699 15620 29708
rect 15568 29665 15577 29699
rect 15577 29665 15611 29699
rect 15611 29665 15620 29699
rect 15568 29656 15620 29665
rect 10140 29588 10192 29640
rect 6184 29452 6236 29504
rect 8576 29452 8628 29504
rect 9772 29452 9824 29504
rect 12716 29495 12768 29504
rect 12716 29461 12725 29495
rect 12725 29461 12759 29495
rect 12759 29461 12768 29495
rect 12716 29452 12768 29461
rect 16488 29452 16540 29504
rect 4947 29350 4999 29402
rect 5011 29350 5063 29402
rect 5075 29350 5127 29402
rect 5139 29350 5191 29402
rect 12878 29350 12930 29402
rect 12942 29350 12994 29402
rect 13006 29350 13058 29402
rect 13070 29350 13122 29402
rect 20808 29350 20860 29402
rect 20872 29350 20924 29402
rect 20936 29350 20988 29402
rect 21000 29350 21052 29402
rect 8024 29291 8076 29300
rect 8024 29257 8033 29291
rect 8033 29257 8067 29291
rect 8067 29257 8076 29291
rect 8024 29248 8076 29257
rect 12164 29248 12216 29300
rect 1492 29044 1544 29096
rect 9680 29180 9732 29232
rect 12716 29180 12768 29232
rect 15200 29180 15252 29232
rect 4160 29112 4212 29164
rect 13176 29112 13228 29164
rect 16304 29112 16356 29164
rect 4068 29087 4120 29096
rect 4068 29053 4077 29087
rect 4077 29053 4111 29087
rect 4111 29053 4120 29087
rect 4068 29044 4120 29053
rect 4528 29087 4580 29096
rect 4528 29053 4537 29087
rect 4537 29053 4571 29087
rect 4571 29053 4580 29087
rect 4528 29044 4580 29053
rect 7012 29087 7064 29096
rect 3056 28976 3108 29028
rect 3608 28976 3660 29028
rect 4804 28976 4856 29028
rect 7012 29053 7021 29087
rect 7021 29053 7055 29087
rect 7055 29053 7064 29087
rect 7012 29044 7064 29053
rect 7196 29044 7248 29096
rect 8760 29044 8812 29096
rect 10140 29087 10192 29096
rect 10140 29053 10149 29087
rect 10149 29053 10183 29087
rect 10183 29053 10192 29087
rect 10140 29044 10192 29053
rect 10324 29087 10376 29096
rect 10324 29053 10333 29087
rect 10333 29053 10367 29087
rect 10367 29053 10376 29087
rect 10324 29044 10376 29053
rect 11060 29087 11112 29096
rect 11060 29053 11069 29087
rect 11069 29053 11103 29087
rect 11103 29053 11112 29087
rect 11060 29044 11112 29053
rect 12532 29044 12584 29096
rect 16488 29044 16540 29096
rect 11244 28976 11296 29028
rect 2780 28951 2832 28960
rect 2780 28917 2789 28951
rect 2789 28917 2823 28951
rect 2823 28917 2832 28951
rect 11336 28951 11388 28960
rect 2780 28908 2832 28917
rect 11336 28917 11345 28951
rect 11345 28917 11379 28951
rect 11379 28917 11388 28951
rect 11336 28908 11388 28917
rect 15292 28976 15344 29028
rect 15384 28976 15436 29028
rect 8912 28806 8964 28858
rect 8976 28806 9028 28858
rect 9040 28806 9092 28858
rect 9104 28806 9156 28858
rect 16843 28806 16895 28858
rect 16907 28806 16959 28858
rect 16971 28806 17023 28858
rect 17035 28806 17087 28858
rect 4068 28704 4120 28756
rect 3792 28636 3844 28688
rect 4344 28636 4396 28688
rect 2688 28568 2740 28620
rect 2964 28568 3016 28620
rect 1492 28500 1544 28552
rect 3056 28500 3108 28552
rect 5816 28704 5868 28756
rect 6828 28704 6880 28756
rect 15108 28704 15160 28756
rect 15384 28704 15436 28756
rect 17592 28747 17644 28756
rect 17592 28713 17601 28747
rect 17601 28713 17635 28747
rect 17635 28713 17644 28747
rect 17592 28704 17644 28713
rect 13728 28636 13780 28688
rect 6184 28568 6236 28620
rect 8300 28611 8352 28620
rect 8300 28577 8309 28611
rect 8309 28577 8343 28611
rect 8343 28577 8352 28611
rect 8300 28568 8352 28577
rect 11336 28568 11388 28620
rect 12624 28568 12676 28620
rect 15200 28568 15252 28620
rect 16120 28611 16172 28620
rect 16120 28577 16129 28611
rect 16129 28577 16163 28611
rect 16163 28577 16172 28611
rect 16120 28568 16172 28577
rect 4804 28500 4856 28552
rect 6828 28500 6880 28552
rect 12348 28500 12400 28552
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 15844 28500 15896 28552
rect 4528 28475 4580 28484
rect 4528 28441 4537 28475
rect 4537 28441 4571 28475
rect 4571 28441 4580 28475
rect 4528 28432 4580 28441
rect 5264 28432 5316 28484
rect 16028 28432 16080 28484
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 16580 28500 16632 28509
rect 3976 28364 4028 28416
rect 4344 28364 4396 28416
rect 4804 28364 4856 28416
rect 6460 28364 6512 28416
rect 7288 28364 7340 28416
rect 13912 28364 13964 28416
rect 15568 28407 15620 28416
rect 15568 28373 15577 28407
rect 15577 28373 15611 28407
rect 15611 28373 15620 28407
rect 15568 28364 15620 28373
rect 4947 28262 4999 28314
rect 5011 28262 5063 28314
rect 5075 28262 5127 28314
rect 5139 28262 5191 28314
rect 12878 28262 12930 28314
rect 12942 28262 12994 28314
rect 13006 28262 13058 28314
rect 13070 28262 13122 28314
rect 20808 28262 20860 28314
rect 20872 28262 20924 28314
rect 20936 28262 20988 28314
rect 21000 28262 21052 28314
rect 2780 28203 2832 28212
rect 2780 28169 2789 28203
rect 2789 28169 2823 28203
rect 2823 28169 2832 28203
rect 2780 28160 2832 28169
rect 3148 28160 3200 28212
rect 12624 28203 12676 28212
rect 12624 28169 12633 28203
rect 12633 28169 12667 28203
rect 12667 28169 12676 28203
rect 12624 28160 12676 28169
rect 15936 28160 15988 28212
rect 4620 28067 4672 28076
rect 4620 28033 4629 28067
rect 4629 28033 4663 28067
rect 4663 28033 4672 28067
rect 4620 28024 4672 28033
rect 1492 27956 1544 28008
rect 1676 27999 1728 28008
rect 1676 27965 1685 27999
rect 1685 27965 1719 27999
rect 1719 27965 1728 27999
rect 1676 27956 1728 27965
rect 2872 27956 2924 28008
rect 7196 28092 7248 28144
rect 8668 28092 8720 28144
rect 9680 28092 9732 28144
rect 5264 28024 5316 28076
rect 8024 28024 8076 28076
rect 5356 27956 5408 28008
rect 5632 27956 5684 28008
rect 7564 27999 7616 28008
rect 7564 27965 7573 27999
rect 7573 27965 7607 27999
rect 7607 27965 7616 27999
rect 7564 27956 7616 27965
rect 7748 27999 7800 28008
rect 7748 27965 7757 27999
rect 7757 27965 7791 27999
rect 7791 27965 7800 27999
rect 7748 27956 7800 27965
rect 9864 27956 9916 28008
rect 10876 27999 10928 28008
rect 10876 27965 10885 27999
rect 10885 27965 10919 27999
rect 10919 27965 10928 27999
rect 10876 27956 10928 27965
rect 13912 28067 13964 28076
rect 13912 28033 13921 28067
rect 13921 28033 13955 28067
rect 13955 28033 13964 28067
rect 13912 28024 13964 28033
rect 15384 27956 15436 28008
rect 16212 27999 16264 28008
rect 16212 27965 16221 27999
rect 16221 27965 16255 27999
rect 16255 27965 16264 27999
rect 16212 27956 16264 27965
rect 5908 27888 5960 27940
rect 10416 27888 10468 27940
rect 16488 27956 16540 28008
rect 16580 27956 16632 28008
rect 2412 27820 2464 27872
rect 2780 27820 2832 27872
rect 8300 27820 8352 27872
rect 8912 27718 8964 27770
rect 8976 27718 9028 27770
rect 9040 27718 9092 27770
rect 9104 27718 9156 27770
rect 16843 27718 16895 27770
rect 16907 27718 16959 27770
rect 16971 27718 17023 27770
rect 17035 27718 17087 27770
rect 4896 27616 4948 27668
rect 4068 27548 4120 27600
rect 3792 27480 3844 27532
rect 4896 27480 4948 27532
rect 5264 27480 5316 27532
rect 7012 27616 7064 27668
rect 8208 27616 8260 27668
rect 8484 27616 8536 27668
rect 6828 27548 6880 27600
rect 6920 27523 6972 27532
rect 6920 27489 6929 27523
rect 6929 27489 6963 27523
rect 6963 27489 6972 27523
rect 6920 27480 6972 27489
rect 7012 27523 7064 27532
rect 7012 27489 7021 27523
rect 7021 27489 7055 27523
rect 7055 27489 7064 27523
rect 7012 27480 7064 27489
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 9772 27523 9824 27532
rect 9772 27489 9781 27523
rect 9781 27489 9815 27523
rect 9815 27489 9824 27523
rect 9772 27480 9824 27489
rect 3976 27412 4028 27464
rect 4160 27455 4212 27464
rect 4160 27421 4169 27455
rect 4169 27421 4203 27455
rect 4203 27421 4212 27455
rect 4160 27412 4212 27421
rect 6276 27455 6328 27464
rect 6276 27421 6285 27455
rect 6285 27421 6319 27455
rect 6319 27421 6328 27455
rect 6276 27412 6328 27421
rect 8392 27412 8444 27464
rect 8944 27412 8996 27464
rect 9864 27412 9916 27464
rect 10876 27548 10928 27600
rect 13268 27548 13320 27600
rect 10232 27480 10284 27532
rect 11336 27480 11388 27532
rect 15292 27548 15344 27600
rect 11612 27412 11664 27464
rect 13268 27412 13320 27464
rect 12716 27344 12768 27396
rect 13820 27344 13872 27396
rect 2780 27276 2832 27328
rect 3148 27276 3200 27328
rect 5540 27276 5592 27328
rect 6828 27276 6880 27328
rect 7656 27276 7708 27328
rect 8668 27319 8720 27328
rect 8668 27285 8677 27319
rect 8677 27285 8711 27319
rect 8711 27285 8720 27319
rect 8668 27276 8720 27285
rect 11060 27276 11112 27328
rect 15200 27480 15252 27532
rect 15384 27480 15436 27532
rect 15568 27523 15620 27532
rect 15568 27489 15577 27523
rect 15577 27489 15611 27523
rect 15611 27489 15620 27523
rect 15568 27480 15620 27489
rect 16028 27412 16080 27464
rect 15568 27276 15620 27328
rect 16212 27276 16264 27328
rect 4947 27174 4999 27226
rect 5011 27174 5063 27226
rect 5075 27174 5127 27226
rect 5139 27174 5191 27226
rect 12878 27174 12930 27226
rect 12942 27174 12994 27226
rect 13006 27174 13058 27226
rect 13070 27174 13122 27226
rect 20808 27174 20860 27226
rect 20872 27174 20924 27226
rect 20936 27174 20988 27226
rect 21000 27174 21052 27226
rect 3056 27072 3108 27124
rect 4160 27072 4212 27124
rect 6276 27072 6328 27124
rect 6828 27072 6880 27124
rect 8852 27072 8904 27124
rect 9680 27072 9732 27124
rect 11428 27115 11480 27124
rect 11428 27081 11437 27115
rect 11437 27081 11471 27115
rect 11471 27081 11480 27115
rect 11428 27072 11480 27081
rect 11980 27072 12032 27124
rect 12348 27072 12400 27124
rect 16028 27072 16080 27124
rect 16120 27072 16172 27124
rect 3976 27004 4028 27056
rect 8300 27004 8352 27056
rect 12072 27004 12124 27056
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 3148 26979 3200 26988
rect 2872 26936 2924 26945
rect 3148 26945 3157 26979
rect 3157 26945 3191 26979
rect 3191 26945 3200 26979
rect 3148 26936 3200 26945
rect 3792 26936 3844 26988
rect 4068 26936 4120 26988
rect 4160 26936 4212 26988
rect 4528 26936 4580 26988
rect 4068 26800 4120 26852
rect 7748 26936 7800 26988
rect 6828 26911 6880 26920
rect 6828 26877 6837 26911
rect 6837 26877 6871 26911
rect 6871 26877 6880 26911
rect 6828 26868 6880 26877
rect 1952 26775 2004 26784
rect 1952 26741 1961 26775
rect 1961 26741 1995 26775
rect 1995 26741 2004 26775
rect 1952 26732 2004 26741
rect 3148 26732 3200 26784
rect 4436 26732 4488 26784
rect 4620 26732 4672 26784
rect 6460 26800 6512 26852
rect 7656 26868 7708 26920
rect 8024 26911 8076 26920
rect 8024 26877 8033 26911
rect 8033 26877 8067 26911
rect 8067 26877 8076 26911
rect 8024 26868 8076 26877
rect 8300 26911 8352 26920
rect 8300 26877 8329 26911
rect 8329 26877 8352 26911
rect 8300 26868 8352 26877
rect 8852 26868 8904 26920
rect 8208 26843 8260 26852
rect 8208 26809 8217 26843
rect 8217 26809 8251 26843
rect 8251 26809 8260 26843
rect 8208 26800 8260 26809
rect 8944 26800 8996 26852
rect 9680 26936 9732 26988
rect 9220 26868 9272 26920
rect 9772 26911 9824 26920
rect 9772 26877 9781 26911
rect 9781 26877 9815 26911
rect 9815 26877 9824 26911
rect 9772 26868 9824 26877
rect 14188 26936 14240 26988
rect 15384 26936 15436 26988
rect 15936 26936 15988 26988
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 12440 26868 12492 26877
rect 14004 26911 14056 26920
rect 14004 26877 14013 26911
rect 14013 26877 14047 26911
rect 14047 26877 14056 26911
rect 14004 26868 14056 26877
rect 16212 26911 16264 26920
rect 16212 26877 16221 26911
rect 16221 26877 16255 26911
rect 16255 26877 16264 26911
rect 16212 26868 16264 26877
rect 16488 26868 16540 26920
rect 7012 26775 7064 26784
rect 7012 26741 7021 26775
rect 7021 26741 7055 26775
rect 7055 26741 7064 26775
rect 7012 26732 7064 26741
rect 7564 26732 7616 26784
rect 8300 26732 8352 26784
rect 8392 26732 8444 26784
rect 15200 26732 15252 26784
rect 18144 26775 18196 26784
rect 18144 26741 18153 26775
rect 18153 26741 18187 26775
rect 18187 26741 18196 26775
rect 18144 26732 18196 26741
rect 8912 26630 8964 26682
rect 8976 26630 9028 26682
rect 9040 26630 9092 26682
rect 9104 26630 9156 26682
rect 16843 26630 16895 26682
rect 16907 26630 16959 26682
rect 16971 26630 17023 26682
rect 17035 26630 17087 26682
rect 1492 26528 1544 26580
rect 1768 26528 1820 26580
rect 3332 26528 3384 26580
rect 3976 26528 4028 26580
rect 6000 26571 6052 26580
rect 6000 26537 6009 26571
rect 6009 26537 6043 26571
rect 6043 26537 6052 26571
rect 6000 26528 6052 26537
rect 3792 26460 3844 26512
rect 2596 26392 2648 26444
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 2780 26392 2832 26401
rect 3148 26392 3200 26444
rect 4068 26435 4120 26444
rect 4068 26401 4077 26435
rect 4077 26401 4111 26435
rect 4111 26401 4120 26435
rect 4068 26392 4120 26401
rect 2228 26324 2280 26376
rect 2688 26324 2740 26376
rect 3056 26324 3108 26376
rect 5816 26392 5868 26444
rect 6000 26392 6052 26444
rect 6920 26528 6972 26580
rect 8208 26528 8260 26580
rect 8668 26528 8720 26580
rect 9220 26528 9272 26580
rect 9772 26528 9824 26580
rect 7288 26460 7340 26512
rect 10416 26503 10468 26512
rect 10416 26469 10425 26503
rect 10425 26469 10459 26503
rect 10459 26469 10468 26503
rect 10416 26460 10468 26469
rect 12716 26460 12768 26512
rect 16488 26460 16540 26512
rect 7564 26392 7616 26444
rect 7656 26392 7708 26444
rect 4068 26256 4120 26308
rect 5264 26256 5316 26308
rect 7012 26324 7064 26376
rect 9772 26392 9824 26444
rect 11980 26392 12032 26444
rect 13728 26435 13780 26444
rect 13728 26401 13737 26435
rect 13737 26401 13771 26435
rect 13771 26401 13780 26435
rect 13728 26392 13780 26401
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 12716 26324 12768 26376
rect 15200 26392 15252 26444
rect 18052 26392 18104 26444
rect 15384 26324 15436 26376
rect 16028 26324 16080 26376
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 8024 26299 8076 26308
rect 8024 26265 8033 26299
rect 8033 26265 8067 26299
rect 8067 26265 8076 26299
rect 8024 26256 8076 26265
rect 10600 26256 10652 26308
rect 1860 26231 1912 26240
rect 1860 26197 1869 26231
rect 1869 26197 1903 26231
rect 1903 26197 1912 26231
rect 1860 26188 1912 26197
rect 3516 26188 3568 26240
rect 4436 26188 4488 26240
rect 6460 26188 6512 26240
rect 6828 26188 6880 26240
rect 9864 26188 9916 26240
rect 10416 26188 10468 26240
rect 15568 26188 15620 26240
rect 17960 26231 18012 26240
rect 17960 26197 17969 26231
rect 17969 26197 18003 26231
rect 18003 26197 18012 26231
rect 17960 26188 18012 26197
rect 4947 26086 4999 26138
rect 5011 26086 5063 26138
rect 5075 26086 5127 26138
rect 5139 26086 5191 26138
rect 12878 26086 12930 26138
rect 12942 26086 12994 26138
rect 13006 26086 13058 26138
rect 13070 26086 13122 26138
rect 20808 26086 20860 26138
rect 20872 26086 20924 26138
rect 20936 26086 20988 26138
rect 21000 26086 21052 26138
rect 8024 26027 8076 26036
rect 8024 25993 8033 26027
rect 8033 25993 8067 26027
rect 8067 25993 8076 26027
rect 8024 25984 8076 25993
rect 9496 25984 9548 26036
rect 10600 26027 10652 26036
rect 10600 25993 10609 26027
rect 10609 25993 10643 26027
rect 10643 25993 10652 26027
rect 10600 25984 10652 25993
rect 14004 25984 14056 26036
rect 12072 25916 12124 25968
rect 18144 25916 18196 25968
rect 1860 25848 1912 25900
rect 3884 25848 3936 25900
rect 4344 25848 4396 25900
rect 2872 25780 2924 25832
rect 5356 25848 5408 25900
rect 11152 25848 11204 25900
rect 14556 25848 14608 25900
rect 15384 25891 15436 25900
rect 15384 25857 15393 25891
rect 15393 25857 15427 25891
rect 15427 25857 15436 25891
rect 15384 25848 15436 25857
rect 3148 25712 3200 25764
rect 5264 25780 5316 25832
rect 7840 25823 7892 25832
rect 7840 25789 7849 25823
rect 7849 25789 7883 25823
rect 7883 25789 7892 25823
rect 7840 25780 7892 25789
rect 8668 25780 8720 25832
rect 9404 25780 9456 25832
rect 11060 25780 11112 25832
rect 11428 25780 11480 25832
rect 12624 25823 12676 25832
rect 12624 25789 12633 25823
rect 12633 25789 12667 25823
rect 12667 25789 12676 25823
rect 12624 25780 12676 25789
rect 15292 25823 15344 25832
rect 1952 25644 2004 25696
rect 5632 25712 5684 25764
rect 7748 25755 7800 25764
rect 7748 25721 7757 25755
rect 7757 25721 7791 25755
rect 7791 25721 7800 25755
rect 7748 25712 7800 25721
rect 8576 25712 8628 25764
rect 9496 25712 9548 25764
rect 10692 25712 10744 25764
rect 15292 25789 15301 25823
rect 15301 25789 15335 25823
rect 15335 25789 15344 25823
rect 15292 25780 15344 25789
rect 15568 25780 15620 25832
rect 16212 25848 16264 25900
rect 16580 25780 16632 25832
rect 16120 25712 16172 25764
rect 7104 25644 7156 25696
rect 8024 25644 8076 25696
rect 9220 25687 9272 25696
rect 9220 25653 9229 25687
rect 9229 25653 9263 25687
rect 9263 25653 9272 25687
rect 9220 25644 9272 25653
rect 15200 25644 15252 25696
rect 16212 25644 16264 25696
rect 8912 25542 8964 25594
rect 8976 25542 9028 25594
rect 9040 25542 9092 25594
rect 9104 25542 9156 25594
rect 16843 25542 16895 25594
rect 16907 25542 16959 25594
rect 16971 25542 17023 25594
rect 17035 25542 17087 25594
rect 5724 25440 5776 25492
rect 1676 25372 1728 25424
rect 1768 25304 1820 25356
rect 3056 25372 3108 25424
rect 2412 25347 2464 25356
rect 2412 25313 2421 25347
rect 2421 25313 2455 25347
rect 2455 25313 2464 25347
rect 2412 25304 2464 25313
rect 2872 25304 2924 25356
rect 7104 25347 7156 25356
rect 7104 25313 7113 25347
rect 7113 25313 7147 25347
rect 7147 25313 7156 25347
rect 7104 25304 7156 25313
rect 11520 25440 11572 25492
rect 7656 25415 7708 25424
rect 7656 25381 7665 25415
rect 7665 25381 7699 25415
rect 7699 25381 7708 25415
rect 7656 25372 7708 25381
rect 15936 25440 15988 25492
rect 13268 25415 13320 25424
rect 8576 25304 8628 25356
rect 9680 25347 9732 25356
rect 9680 25313 9689 25347
rect 9689 25313 9723 25347
rect 9723 25313 9732 25347
rect 9680 25304 9732 25313
rect 11244 25347 11296 25356
rect 2228 25236 2280 25288
rect 4712 25279 4764 25288
rect 2412 25168 2464 25220
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 8208 25168 8260 25220
rect 11244 25313 11253 25347
rect 11253 25313 11287 25347
rect 11287 25313 11296 25347
rect 11244 25304 11296 25313
rect 11428 25304 11480 25356
rect 13268 25381 13277 25415
rect 13277 25381 13311 25415
rect 13311 25381 13320 25415
rect 13268 25372 13320 25381
rect 15384 25372 15436 25424
rect 17960 25372 18012 25424
rect 13636 25304 13688 25356
rect 16028 25347 16080 25356
rect 16028 25313 16037 25347
rect 16037 25313 16071 25347
rect 16071 25313 16080 25347
rect 16028 25304 16080 25313
rect 15384 25236 15436 25288
rect 15844 25236 15896 25288
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 7380 25100 7432 25152
rect 11060 25100 11112 25152
rect 4947 24998 4999 25050
rect 5011 24998 5063 25050
rect 5075 24998 5127 25050
rect 5139 24998 5191 25050
rect 12878 24998 12930 25050
rect 12942 24998 12994 25050
rect 13006 24998 13058 25050
rect 13070 24998 13122 25050
rect 20808 24998 20860 25050
rect 20872 24998 20924 25050
rect 20936 24998 20988 25050
rect 21000 24998 21052 25050
rect 4712 24939 4764 24948
rect 4712 24905 4721 24939
rect 4721 24905 4755 24939
rect 4755 24905 4764 24939
rect 4712 24896 4764 24905
rect 4068 24828 4120 24880
rect 17500 24896 17552 24948
rect 5724 24828 5776 24880
rect 5816 24828 5868 24880
rect 9864 24828 9916 24880
rect 11888 24828 11940 24880
rect 15936 24828 15988 24880
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 7748 24803 7800 24812
rect 2320 24735 2372 24744
rect 2320 24701 2329 24735
rect 2329 24701 2363 24735
rect 2363 24701 2372 24735
rect 2320 24692 2372 24701
rect 2412 24692 2464 24744
rect 3516 24735 3568 24744
rect 3516 24701 3525 24735
rect 3525 24701 3559 24735
rect 3559 24701 3568 24735
rect 3516 24692 3568 24701
rect 4068 24692 4120 24744
rect 4344 24692 4396 24744
rect 7012 24692 7064 24744
rect 7196 24692 7248 24744
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 7840 24760 7892 24812
rect 10416 24760 10468 24812
rect 10692 24760 10744 24812
rect 8576 24692 8628 24744
rect 10876 24692 10928 24744
rect 7840 24556 7892 24608
rect 9220 24624 9272 24676
rect 11336 24692 11388 24744
rect 12624 24735 12676 24744
rect 12624 24701 12633 24735
rect 12633 24701 12667 24735
rect 12667 24701 12676 24735
rect 12624 24692 12676 24701
rect 14188 24692 14240 24744
rect 14648 24692 14700 24744
rect 14740 24692 14792 24744
rect 19156 24735 19208 24744
rect 19156 24701 19165 24735
rect 19165 24701 19199 24735
rect 19199 24701 19208 24735
rect 19156 24692 19208 24701
rect 13452 24624 13504 24676
rect 16488 24624 16540 24676
rect 17592 24624 17644 24676
rect 9956 24556 10008 24608
rect 10232 24556 10284 24608
rect 11428 24556 11480 24608
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 8912 24454 8964 24506
rect 8976 24454 9028 24506
rect 9040 24454 9092 24506
rect 9104 24454 9156 24506
rect 16843 24454 16895 24506
rect 16907 24454 16959 24506
rect 16971 24454 17023 24506
rect 17035 24454 17087 24506
rect 1768 24352 1820 24404
rect 5540 24352 5592 24404
rect 6920 24352 6972 24404
rect 8576 24352 8628 24404
rect 9220 24352 9272 24404
rect 2688 24284 2740 24336
rect 9680 24284 9732 24336
rect 10140 24284 10192 24336
rect 11888 24284 11940 24336
rect 13728 24284 13780 24336
rect 16304 24352 16356 24404
rect 2504 24216 2556 24268
rect 2596 24259 2648 24268
rect 2596 24225 2605 24259
rect 2605 24225 2639 24259
rect 2639 24225 2648 24259
rect 2596 24216 2648 24225
rect 6920 24216 6972 24268
rect 2136 24148 2188 24200
rect 2688 24148 2740 24200
rect 5356 24148 5408 24200
rect 6828 24148 6880 24200
rect 7380 24216 7432 24268
rect 7564 24216 7616 24268
rect 7840 24216 7892 24268
rect 8300 24216 8352 24268
rect 8668 24216 8720 24268
rect 10692 24259 10744 24268
rect 8024 24148 8076 24200
rect 8208 24148 8260 24200
rect 10692 24225 10701 24259
rect 10701 24225 10735 24259
rect 10735 24225 10744 24259
rect 10692 24216 10744 24225
rect 11244 24216 11296 24268
rect 11428 24216 11480 24268
rect 11980 24259 12032 24268
rect 11980 24225 11989 24259
rect 11989 24225 12023 24259
rect 12023 24225 12032 24259
rect 11980 24216 12032 24225
rect 12072 24216 12124 24268
rect 14740 24216 14792 24268
rect 11060 24148 11112 24200
rect 11244 24080 11296 24132
rect 13912 24148 13964 24200
rect 14924 24148 14976 24200
rect 16672 24284 16724 24336
rect 17960 24284 18012 24336
rect 18420 24284 18472 24336
rect 15844 24216 15896 24268
rect 17132 24216 17184 24268
rect 18144 24259 18196 24268
rect 18144 24225 18153 24259
rect 18153 24225 18187 24259
rect 18187 24225 18196 24259
rect 18144 24216 18196 24225
rect 16488 24148 16540 24200
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 19156 24080 19208 24132
rect 2412 24012 2464 24064
rect 7012 24012 7064 24064
rect 9680 24055 9732 24064
rect 9680 24021 9689 24055
rect 9689 24021 9723 24055
rect 9723 24021 9732 24055
rect 10140 24055 10192 24064
rect 9680 24012 9732 24021
rect 10140 24021 10149 24055
rect 10149 24021 10183 24055
rect 10183 24021 10192 24055
rect 10140 24012 10192 24021
rect 10600 24012 10652 24064
rect 14372 24012 14424 24064
rect 4947 23910 4999 23962
rect 5011 23910 5063 23962
rect 5075 23910 5127 23962
rect 5139 23910 5191 23962
rect 12878 23910 12930 23962
rect 12942 23910 12994 23962
rect 13006 23910 13058 23962
rect 13070 23910 13122 23962
rect 20808 23910 20860 23962
rect 20872 23910 20924 23962
rect 20936 23910 20988 23962
rect 21000 23910 21052 23962
rect 1308 23808 1360 23860
rect 2136 23740 2188 23792
rect 2504 23808 2556 23860
rect 2688 23808 2740 23860
rect 7104 23808 7156 23860
rect 10692 23808 10744 23860
rect 11796 23808 11848 23860
rect 18512 23808 18564 23860
rect 5816 23740 5868 23792
rect 1768 23604 1820 23656
rect 2228 23647 2280 23656
rect 2228 23613 2237 23647
rect 2237 23613 2271 23647
rect 2271 23613 2280 23647
rect 2688 23672 2740 23724
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 4344 23672 4396 23724
rect 2228 23604 2280 23613
rect 2596 23647 2648 23656
rect 2596 23613 2605 23647
rect 2605 23613 2639 23647
rect 2639 23613 2648 23647
rect 2596 23604 2648 23613
rect 1676 23536 1728 23588
rect 4712 23604 4764 23656
rect 5540 23604 5592 23656
rect 5816 23604 5868 23656
rect 7012 23647 7064 23656
rect 7012 23613 7021 23647
rect 7021 23613 7055 23647
rect 7055 23613 7064 23647
rect 7012 23604 7064 23613
rect 7104 23647 7156 23656
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 4988 23536 5040 23588
rect 14372 23740 14424 23792
rect 14648 23783 14700 23792
rect 14648 23749 14657 23783
rect 14657 23749 14691 23783
rect 14691 23749 14700 23783
rect 14648 23740 14700 23749
rect 15108 23740 15160 23792
rect 16488 23740 16540 23792
rect 10876 23672 10928 23724
rect 11152 23672 11204 23724
rect 11612 23672 11664 23724
rect 8668 23604 8720 23656
rect 9496 23604 9548 23656
rect 12348 23604 12400 23656
rect 13912 23672 13964 23724
rect 15752 23715 15804 23724
rect 15752 23681 15761 23715
rect 15761 23681 15795 23715
rect 15795 23681 15804 23715
rect 15752 23672 15804 23681
rect 16212 23715 16264 23724
rect 16212 23681 16221 23715
rect 16221 23681 16255 23715
rect 16255 23681 16264 23715
rect 16212 23672 16264 23681
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 16488 23604 16540 23656
rect 16672 23604 16724 23656
rect 18328 23672 18380 23724
rect 17132 23604 17184 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18512 23604 18564 23656
rect 7380 23536 7432 23588
rect 9220 23536 9272 23588
rect 13084 23536 13136 23588
rect 14556 23536 14608 23588
rect 15108 23536 15160 23588
rect 18420 23536 18472 23588
rect 3516 23468 3568 23520
rect 3792 23468 3844 23520
rect 7012 23468 7064 23520
rect 7288 23468 7340 23520
rect 8300 23468 8352 23520
rect 11796 23468 11848 23520
rect 11888 23468 11940 23520
rect 12348 23468 12400 23520
rect 12624 23511 12676 23520
rect 12624 23477 12633 23511
rect 12633 23477 12667 23511
rect 12667 23477 12676 23511
rect 12624 23468 12676 23477
rect 13360 23468 13412 23520
rect 13820 23468 13872 23520
rect 17592 23468 17644 23520
rect 17868 23468 17920 23520
rect 8912 23366 8964 23418
rect 8976 23366 9028 23418
rect 9040 23366 9092 23418
rect 9104 23366 9156 23418
rect 16843 23366 16895 23418
rect 16907 23366 16959 23418
rect 16971 23366 17023 23418
rect 17035 23366 17087 23418
rect 2688 23264 2740 23316
rect 4068 23264 4120 23316
rect 8300 23264 8352 23316
rect 1676 23171 1728 23180
rect 1676 23137 1685 23171
rect 1685 23137 1719 23171
rect 1719 23137 1728 23171
rect 1676 23128 1728 23137
rect 3884 23128 3936 23180
rect 5356 23239 5408 23248
rect 5356 23205 5365 23239
rect 5365 23205 5399 23239
rect 5399 23205 5408 23239
rect 5356 23196 5408 23205
rect 9496 23196 9548 23248
rect 9864 23196 9916 23248
rect 11796 23264 11848 23316
rect 12256 23264 12308 23316
rect 13084 23264 13136 23316
rect 4988 23171 5040 23180
rect 4988 23137 4997 23171
rect 4997 23137 5031 23171
rect 5031 23137 5040 23171
rect 4988 23128 5040 23137
rect 7380 23171 7432 23180
rect 7380 23137 7389 23171
rect 7389 23137 7423 23171
rect 7423 23137 7432 23171
rect 7380 23128 7432 23137
rect 10140 23171 10192 23180
rect 10140 23137 10149 23171
rect 10149 23137 10183 23171
rect 10183 23137 10192 23171
rect 10140 23128 10192 23137
rect 11428 23128 11480 23180
rect 11888 23196 11940 23248
rect 12440 23196 12492 23248
rect 16488 23264 16540 23316
rect 16580 23196 16632 23248
rect 2504 23060 2556 23112
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 5908 23060 5960 23112
rect 12256 23128 12308 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 12716 23060 12768 23112
rect 13360 22992 13412 23044
rect 13452 22992 13504 23044
rect 13636 22992 13688 23044
rect 18144 23196 18196 23248
rect 17132 23128 17184 23180
rect 17868 23128 17920 23180
rect 17960 23128 18012 23180
rect 18696 23128 18748 23180
rect 19248 23060 19300 23112
rect 15200 22992 15252 23044
rect 1860 22924 1912 22976
rect 7564 22924 7616 22976
rect 9956 22924 10008 22976
rect 18236 22924 18288 22976
rect 19432 22924 19484 22976
rect 4947 22822 4999 22874
rect 5011 22822 5063 22874
rect 5075 22822 5127 22874
rect 5139 22822 5191 22874
rect 12878 22822 12930 22874
rect 12942 22822 12994 22874
rect 13006 22822 13058 22874
rect 13070 22822 13122 22874
rect 20808 22822 20860 22874
rect 20872 22822 20924 22874
rect 20936 22822 20988 22874
rect 21000 22822 21052 22874
rect 1860 22763 1912 22772
rect 1860 22729 1869 22763
rect 1869 22729 1903 22763
rect 1903 22729 1912 22763
rect 1860 22720 1912 22729
rect 2688 22720 2740 22772
rect 7104 22720 7156 22772
rect 2320 22652 2372 22704
rect 4068 22652 4120 22704
rect 4436 22652 4488 22704
rect 4712 22652 4764 22704
rect 4988 22652 5040 22704
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 7932 22584 7984 22636
rect 1676 22559 1728 22568
rect 1676 22525 1685 22559
rect 1685 22525 1719 22559
rect 1719 22525 1728 22559
rect 1676 22516 1728 22525
rect 2872 22380 2924 22432
rect 5632 22516 5684 22568
rect 6184 22516 6236 22568
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 7656 22516 7708 22568
rect 7564 22448 7616 22500
rect 8484 22516 8536 22568
rect 11704 22720 11756 22772
rect 13268 22720 13320 22772
rect 13636 22720 13688 22772
rect 18328 22720 18380 22772
rect 19248 22720 19300 22772
rect 10140 22652 10192 22704
rect 14004 22652 14056 22704
rect 15568 22652 15620 22704
rect 13176 22584 13228 22636
rect 10692 22559 10744 22568
rect 10692 22525 10701 22559
rect 10701 22525 10735 22559
rect 10735 22525 10744 22559
rect 10692 22516 10744 22525
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 11612 22516 11664 22568
rect 11888 22516 11940 22568
rect 14832 22584 14884 22636
rect 9680 22448 9732 22500
rect 10416 22448 10468 22500
rect 13728 22516 13780 22568
rect 14740 22448 14792 22500
rect 15936 22516 15988 22568
rect 16488 22652 16540 22704
rect 17684 22652 17736 22704
rect 19432 22652 19484 22704
rect 16304 22627 16356 22636
rect 16304 22593 16313 22627
rect 16313 22593 16347 22627
rect 16347 22593 16356 22627
rect 16304 22584 16356 22593
rect 18604 22627 18656 22636
rect 18604 22593 18613 22627
rect 18613 22593 18647 22627
rect 18647 22593 18656 22627
rect 18604 22584 18656 22593
rect 16672 22516 16724 22568
rect 17132 22516 17184 22568
rect 18236 22559 18288 22568
rect 18236 22525 18245 22559
rect 18245 22525 18279 22559
rect 18279 22525 18288 22559
rect 18236 22516 18288 22525
rect 16580 22448 16632 22500
rect 19156 22448 19208 22500
rect 7104 22423 7156 22432
rect 7104 22389 7113 22423
rect 7113 22389 7147 22423
rect 7147 22389 7156 22423
rect 7104 22380 7156 22389
rect 9404 22380 9456 22432
rect 9588 22380 9640 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 10140 22380 10192 22432
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 14372 22423 14424 22432
rect 14372 22389 14381 22423
rect 14381 22389 14415 22423
rect 14415 22389 14424 22423
rect 14372 22380 14424 22389
rect 14556 22380 14608 22432
rect 19524 22380 19576 22432
rect 8912 22278 8964 22330
rect 8976 22278 9028 22330
rect 9040 22278 9092 22330
rect 9104 22278 9156 22330
rect 16843 22278 16895 22330
rect 16907 22278 16959 22330
rect 16971 22278 17023 22330
rect 17035 22278 17087 22330
rect 8484 22176 8536 22228
rect 13544 22176 13596 22228
rect 14556 22176 14608 22228
rect 15568 22176 15620 22228
rect 17684 22176 17736 22228
rect 7196 22108 7248 22160
rect 2320 22040 2372 22092
rect 4068 21972 4120 22024
rect 3424 21904 3476 21956
rect 2228 21836 2280 21888
rect 4988 22040 5040 22092
rect 5264 22083 5316 22092
rect 5264 22049 5273 22083
rect 5273 22049 5307 22083
rect 5307 22049 5316 22083
rect 5264 22040 5316 22049
rect 8024 22040 8076 22092
rect 11244 22108 11296 22160
rect 5080 21972 5132 22024
rect 5448 21972 5500 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 9680 22040 9732 22092
rect 10140 22040 10192 22092
rect 11152 22040 11204 22092
rect 12256 22040 12308 22092
rect 14372 22040 14424 22092
rect 18236 22040 18288 22092
rect 18696 22083 18748 22092
rect 18696 22049 18705 22083
rect 18705 22049 18739 22083
rect 18739 22049 18748 22083
rect 18696 22040 18748 22049
rect 19524 22040 19576 22092
rect 9864 21972 9916 22024
rect 11428 21972 11480 22024
rect 16120 21972 16172 22024
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 16580 21972 16632 22024
rect 4620 21904 4672 21956
rect 6828 21904 6880 21956
rect 9772 21904 9824 21956
rect 4712 21836 4764 21888
rect 7564 21836 7616 21888
rect 11336 21836 11388 21888
rect 11980 21836 12032 21888
rect 14188 21836 14240 21888
rect 15292 21836 15344 21888
rect 15752 21836 15804 21888
rect 4947 21734 4999 21786
rect 5011 21734 5063 21786
rect 5075 21734 5127 21786
rect 5139 21734 5191 21786
rect 12878 21734 12930 21786
rect 12942 21734 12994 21786
rect 13006 21734 13058 21786
rect 13070 21734 13122 21786
rect 20808 21734 20860 21786
rect 20872 21734 20924 21786
rect 20936 21734 20988 21786
rect 21000 21734 21052 21786
rect 3976 21632 4028 21684
rect 11336 21632 11388 21684
rect 11612 21632 11664 21684
rect 14188 21675 14240 21684
rect 7564 21564 7616 21616
rect 8116 21564 8168 21616
rect 8484 21564 8536 21616
rect 9220 21564 9272 21616
rect 11152 21564 11204 21616
rect 11888 21564 11940 21616
rect 5816 21496 5868 21548
rect 7748 21496 7800 21548
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 3884 21471 3936 21480
rect 3884 21437 3893 21471
rect 3893 21437 3927 21471
rect 3927 21437 3936 21471
rect 4068 21471 4120 21480
rect 3884 21428 3936 21437
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 6552 21428 6604 21480
rect 6920 21428 6972 21480
rect 13176 21539 13228 21548
rect 13176 21505 13185 21539
rect 13185 21505 13219 21539
rect 13219 21505 13228 21539
rect 13176 21496 13228 21505
rect 5724 21360 5776 21412
rect 8116 21403 8168 21412
rect 4344 21335 4396 21344
rect 4344 21301 4353 21335
rect 4353 21301 4387 21335
rect 4387 21301 4396 21335
rect 4344 21292 4396 21301
rect 4712 21292 4764 21344
rect 7656 21292 7708 21344
rect 8116 21369 8125 21403
rect 8125 21369 8159 21403
rect 8159 21369 8168 21403
rect 8116 21360 8168 21369
rect 9588 21471 9640 21480
rect 9588 21437 9597 21471
rect 9597 21437 9631 21471
rect 9631 21437 9640 21471
rect 9772 21471 9824 21480
rect 9588 21428 9640 21437
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 10968 21428 11020 21480
rect 11152 21428 11204 21480
rect 12716 21471 12768 21480
rect 12716 21437 12725 21471
rect 12725 21437 12759 21471
rect 12759 21437 12768 21471
rect 12716 21428 12768 21437
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 16488 21632 16540 21684
rect 14740 21496 14792 21548
rect 17592 21496 17644 21548
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 15844 21428 15896 21437
rect 16304 21428 16356 21480
rect 19248 21496 19300 21548
rect 19064 21471 19116 21480
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 19156 21471 19208 21480
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 10416 21360 10468 21412
rect 13176 21360 13228 21412
rect 18052 21403 18104 21412
rect 18052 21369 18061 21403
rect 18061 21369 18095 21403
rect 18095 21369 18104 21403
rect 18052 21360 18104 21369
rect 18328 21360 18380 21412
rect 11152 21292 11204 21344
rect 11980 21292 12032 21344
rect 20168 21335 20220 21344
rect 20168 21301 20177 21335
rect 20177 21301 20211 21335
rect 20211 21301 20220 21335
rect 20168 21292 20220 21301
rect 8912 21190 8964 21242
rect 8976 21190 9028 21242
rect 9040 21190 9092 21242
rect 9104 21190 9156 21242
rect 16843 21190 16895 21242
rect 16907 21190 16959 21242
rect 16971 21190 17023 21242
rect 17035 21190 17087 21242
rect 4068 21088 4120 21140
rect 20168 21088 20220 21140
rect 3056 21063 3108 21072
rect 3056 21029 3065 21063
rect 3065 21029 3099 21063
rect 3099 21029 3108 21063
rect 3056 21020 3108 21029
rect 3700 21020 3752 21072
rect 6552 21063 6604 21072
rect 6552 21029 6561 21063
rect 6561 21029 6595 21063
rect 6595 21029 6604 21063
rect 6552 21020 6604 21029
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 1676 20927 1728 20936
rect 1676 20893 1685 20927
rect 1685 20893 1719 20927
rect 1719 20893 1728 20927
rect 1676 20884 1728 20893
rect 2320 20952 2372 21004
rect 4344 20995 4396 21004
rect 2504 20884 2556 20936
rect 4344 20961 4353 20995
rect 4353 20961 4387 20995
rect 4387 20961 4396 20995
rect 4344 20952 4396 20961
rect 8484 21020 8536 21072
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 10416 21063 10468 21072
rect 10416 21029 10425 21063
rect 10425 21029 10459 21063
rect 10459 21029 10468 21063
rect 10416 21020 10468 21029
rect 12716 21020 12768 21072
rect 7104 20995 7156 21004
rect 7104 20961 7113 20995
rect 7113 20961 7147 20995
rect 7147 20961 7156 20995
rect 7104 20952 7156 20961
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 7932 20995 7984 21004
rect 6828 20884 6880 20936
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 9128 20952 9180 21004
rect 10600 20952 10652 21004
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 7748 20884 7800 20936
rect 12808 20952 12860 21004
rect 13360 20952 13412 21004
rect 15292 20995 15344 21004
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 15568 20952 15620 21004
rect 18052 20952 18104 21004
rect 19064 20952 19116 21004
rect 7104 20816 7156 20868
rect 9128 20816 9180 20868
rect 6828 20748 6880 20800
rect 11612 20816 11664 20868
rect 16120 20884 16172 20936
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 12532 20816 12584 20868
rect 12624 20816 12676 20868
rect 15568 20816 15620 20868
rect 11336 20791 11388 20800
rect 11336 20757 11345 20791
rect 11345 20757 11379 20791
rect 11379 20757 11388 20791
rect 11336 20748 11388 20757
rect 11888 20748 11940 20800
rect 16304 20748 16356 20800
rect 18236 20748 18288 20800
rect 4947 20646 4999 20698
rect 5011 20646 5063 20698
rect 5075 20646 5127 20698
rect 5139 20646 5191 20698
rect 12878 20646 12930 20698
rect 12942 20646 12994 20698
rect 13006 20646 13058 20698
rect 13070 20646 13122 20698
rect 20808 20646 20860 20698
rect 20872 20646 20924 20698
rect 20936 20646 20988 20698
rect 21000 20646 21052 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 2044 20476 2096 20528
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 2320 20383 2372 20392
rect 2320 20349 2329 20383
rect 2329 20349 2363 20383
rect 2363 20349 2372 20383
rect 3056 20408 3108 20460
rect 2320 20340 2372 20349
rect 4712 20383 4764 20392
rect 2504 20272 2556 20324
rect 4712 20349 4721 20383
rect 4721 20349 4755 20383
rect 4755 20349 4764 20383
rect 4712 20340 4764 20349
rect 4804 20340 4856 20392
rect 7104 20476 7156 20528
rect 7196 20408 7248 20460
rect 8208 20476 8260 20528
rect 8852 20340 8904 20392
rect 9588 20544 9640 20596
rect 15108 20544 15160 20596
rect 18328 20587 18380 20596
rect 18328 20553 18337 20587
rect 18337 20553 18371 20587
rect 18371 20553 18380 20587
rect 18328 20544 18380 20553
rect 11336 20476 11388 20528
rect 11704 20408 11756 20460
rect 11980 20408 12032 20460
rect 13360 20408 13412 20460
rect 15660 20451 15712 20460
rect 9588 20340 9640 20392
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 11152 20340 11204 20392
rect 11336 20340 11388 20392
rect 6920 20272 6972 20324
rect 7564 20315 7616 20324
rect 7564 20281 7573 20315
rect 7573 20281 7607 20315
rect 7607 20281 7616 20315
rect 7564 20272 7616 20281
rect 10968 20272 11020 20324
rect 7012 20204 7064 20256
rect 14372 20340 14424 20392
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 16028 20408 16080 20460
rect 16580 20451 16632 20460
rect 16580 20417 16589 20451
rect 16589 20417 16623 20451
rect 16623 20417 16632 20451
rect 16580 20408 16632 20417
rect 17132 20408 17184 20460
rect 17776 20408 17828 20460
rect 18420 20451 18472 20460
rect 18420 20417 18429 20451
rect 18429 20417 18463 20451
rect 18463 20417 18472 20451
rect 18420 20408 18472 20417
rect 15292 20272 15344 20324
rect 17224 20272 17276 20324
rect 15568 20204 15620 20256
rect 16120 20204 16172 20256
rect 18696 20247 18748 20256
rect 18696 20213 18705 20247
rect 18705 20213 18739 20247
rect 18739 20213 18748 20247
rect 18696 20204 18748 20213
rect 8912 20102 8964 20154
rect 8976 20102 9028 20154
rect 9040 20102 9092 20154
rect 9104 20102 9156 20154
rect 16843 20102 16895 20154
rect 16907 20102 16959 20154
rect 16971 20102 17023 20154
rect 17035 20102 17087 20154
rect 3608 20000 3660 20052
rect 2136 19932 2188 19984
rect 2596 19932 2648 19984
rect 1492 19864 1544 19916
rect 2044 19864 2096 19916
rect 6920 20000 6972 20052
rect 7748 20000 7800 20052
rect 8116 20000 8168 20052
rect 8392 19932 8444 19984
rect 9588 19932 9640 19984
rect 13176 20000 13228 20052
rect 14648 20000 14700 20052
rect 5724 19907 5776 19916
rect 5724 19873 5733 19907
rect 5733 19873 5767 19907
rect 5767 19873 5776 19907
rect 5724 19864 5776 19873
rect 8024 19907 8076 19916
rect 8024 19873 8033 19907
rect 8033 19873 8067 19907
rect 8067 19873 8076 19907
rect 8024 19864 8076 19873
rect 8208 19864 8260 19916
rect 9772 19864 9824 19916
rect 13544 19932 13596 19984
rect 13636 19932 13688 19984
rect 11060 19864 11112 19916
rect 11428 19864 11480 19916
rect 12624 19864 12676 19916
rect 2688 19796 2740 19848
rect 3056 19796 3108 19848
rect 5908 19796 5960 19848
rect 2136 19728 2188 19780
rect 8116 19771 8168 19780
rect 8116 19737 8125 19771
rect 8125 19737 8159 19771
rect 8159 19737 8168 19771
rect 8116 19728 8168 19737
rect 9588 19728 9640 19780
rect 9864 19728 9916 19780
rect 2596 19660 2648 19712
rect 2780 19660 2832 19712
rect 2964 19660 3016 19712
rect 7748 19660 7800 19712
rect 8300 19660 8352 19712
rect 10416 19660 10468 19712
rect 13544 19660 13596 19712
rect 14648 19660 14700 19712
rect 17592 19864 17644 19916
rect 17776 19907 17828 19916
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 17960 19907 18012 19916
rect 17960 19873 17969 19907
rect 17969 19873 18003 19907
rect 18003 19873 18012 19907
rect 17960 19864 18012 19873
rect 18604 19864 18656 19916
rect 19156 19864 19208 19916
rect 16672 19660 16724 19712
rect 4947 19558 4999 19610
rect 5011 19558 5063 19610
rect 5075 19558 5127 19610
rect 5139 19558 5191 19610
rect 12878 19558 12930 19610
rect 12942 19558 12994 19610
rect 13006 19558 13058 19610
rect 13070 19558 13122 19610
rect 20808 19558 20860 19610
rect 20872 19558 20924 19610
rect 20936 19558 20988 19610
rect 21000 19558 21052 19610
rect 2596 19456 2648 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 5908 19456 5960 19508
rect 7748 19456 7800 19508
rect 2688 19388 2740 19440
rect 3056 19363 3108 19372
rect 3056 19329 3065 19363
rect 3065 19329 3099 19363
rect 3099 19329 3108 19363
rect 3056 19320 3108 19329
rect 3608 19320 3660 19372
rect 5448 19388 5500 19440
rect 6184 19388 6236 19440
rect 6552 19388 6604 19440
rect 8116 19456 8168 19508
rect 13360 19456 13412 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 18236 19456 18288 19508
rect 10876 19388 10928 19440
rect 10968 19388 11020 19440
rect 16120 19363 16172 19372
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2964 19252 3016 19304
rect 4344 19252 4396 19304
rect 4712 19252 4764 19304
rect 6184 19252 6236 19304
rect 7012 19252 7064 19304
rect 8300 19252 8352 19304
rect 10416 19252 10468 19304
rect 10968 19252 11020 19304
rect 2412 19184 2464 19236
rect 3424 19227 3476 19236
rect 3424 19193 3433 19227
rect 3433 19193 3467 19227
rect 3467 19193 3476 19227
rect 3424 19184 3476 19193
rect 4620 19184 4672 19236
rect 7748 19184 7800 19236
rect 10692 19227 10744 19236
rect 10692 19193 10701 19227
rect 10701 19193 10735 19227
rect 10735 19193 10744 19227
rect 10692 19184 10744 19193
rect 10876 19184 10928 19236
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 11152 19184 11204 19236
rect 13176 19184 13228 19236
rect 13728 19252 13780 19304
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 15476 19252 15528 19304
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 17132 19320 17184 19372
rect 18236 19363 18288 19372
rect 14188 19184 14240 19236
rect 16488 19295 16540 19304
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 18236 19329 18242 19363
rect 18242 19329 18288 19363
rect 18236 19320 18288 19329
rect 16488 19252 16540 19261
rect 17868 19252 17920 19304
rect 16580 19184 16632 19236
rect 17132 19184 17184 19236
rect 4344 19116 4396 19168
rect 7380 19116 7432 19168
rect 8208 19116 8260 19168
rect 9680 19116 9732 19168
rect 10048 19116 10100 19168
rect 15752 19116 15804 19168
rect 16304 19116 16356 19168
rect 18328 19116 18380 19168
rect 8912 19014 8964 19066
rect 8976 19014 9028 19066
rect 9040 19014 9092 19066
rect 9104 19014 9156 19066
rect 16843 19014 16895 19066
rect 16907 19014 16959 19066
rect 16971 19014 17023 19066
rect 17035 19014 17087 19066
rect 1492 18912 1544 18964
rect 2412 18912 2464 18964
rect 6460 18912 6512 18964
rect 4528 18844 4580 18896
rect 4620 18776 4672 18828
rect 7288 18819 7340 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 3884 18708 3936 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 5632 18708 5684 18760
rect 3516 18572 3568 18624
rect 7288 18785 7297 18819
rect 7297 18785 7331 18819
rect 7331 18785 7340 18819
rect 7288 18776 7340 18785
rect 7656 18912 7708 18964
rect 10140 18912 10192 18964
rect 10876 18912 10928 18964
rect 13728 18912 13780 18964
rect 18236 18912 18288 18964
rect 10416 18844 10468 18896
rect 7380 18708 7432 18760
rect 7472 18708 7524 18760
rect 10784 18819 10836 18828
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 11796 18776 11848 18828
rect 12624 18776 12676 18828
rect 13636 18776 13688 18828
rect 16028 18844 16080 18896
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 15200 18776 15252 18828
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 16672 18776 16724 18828
rect 17868 18776 17920 18828
rect 7656 18640 7708 18692
rect 9588 18708 9640 18760
rect 13912 18751 13964 18760
rect 10048 18640 10100 18692
rect 13912 18717 13921 18751
rect 13921 18717 13955 18751
rect 13955 18717 13964 18751
rect 13912 18708 13964 18717
rect 15476 18708 15528 18760
rect 9680 18572 9732 18624
rect 15752 18572 15804 18624
rect 19524 18640 19576 18692
rect 17868 18572 17920 18624
rect 4947 18470 4999 18522
rect 5011 18470 5063 18522
rect 5075 18470 5127 18522
rect 5139 18470 5191 18522
rect 12878 18470 12930 18522
rect 12942 18470 12994 18522
rect 13006 18470 13058 18522
rect 13070 18470 13122 18522
rect 20808 18470 20860 18522
rect 20872 18470 20924 18522
rect 20936 18470 20988 18522
rect 21000 18470 21052 18522
rect 8300 18368 8352 18420
rect 8576 18368 8628 18420
rect 10140 18368 10192 18420
rect 11152 18300 11204 18352
rect 2504 18232 2556 18284
rect 3516 18275 3568 18284
rect 2688 18164 2740 18216
rect 3056 18164 3108 18216
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 4160 18232 4212 18284
rect 4344 18232 4396 18284
rect 6828 18232 6880 18284
rect 8208 18232 8260 18284
rect 11244 18275 11296 18284
rect 1768 18096 1820 18148
rect 7472 18164 7524 18216
rect 8576 18207 8628 18216
rect 1400 18028 1452 18080
rect 4896 18096 4948 18148
rect 6368 18096 6420 18148
rect 7564 18096 7616 18148
rect 3608 18028 3660 18080
rect 4344 18028 4396 18080
rect 5540 18028 5592 18080
rect 5908 18028 5960 18080
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 10784 18207 10836 18216
rect 10784 18173 10793 18207
rect 10793 18173 10827 18207
rect 10827 18173 10836 18207
rect 10784 18164 10836 18173
rect 11244 18241 11253 18275
rect 11253 18241 11287 18275
rect 11287 18241 11296 18275
rect 11244 18232 11296 18241
rect 12716 18232 12768 18284
rect 13360 18300 13412 18352
rect 13728 18300 13780 18352
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 13912 18164 13964 18216
rect 15476 18207 15528 18216
rect 15476 18173 15485 18207
rect 15485 18173 15519 18207
rect 15519 18173 15528 18207
rect 15476 18164 15528 18173
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 17960 18164 18012 18216
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 13636 18096 13688 18148
rect 17868 18096 17920 18148
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 15292 18028 15344 18080
rect 16396 18028 16448 18080
rect 8912 17926 8964 17978
rect 8976 17926 9028 17978
rect 9040 17926 9092 17978
rect 9104 17926 9156 17978
rect 16843 17926 16895 17978
rect 16907 17926 16959 17978
rect 16971 17926 17023 17978
rect 17035 17926 17087 17978
rect 4620 17824 4672 17876
rect 7012 17867 7064 17876
rect 7012 17833 7021 17867
rect 7021 17833 7055 17867
rect 7055 17833 7064 17867
rect 7012 17824 7064 17833
rect 12440 17824 12492 17876
rect 14372 17824 14424 17876
rect 15752 17824 15804 17876
rect 1676 17756 1728 17808
rect 5540 17756 5592 17808
rect 13912 17756 13964 17808
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 2504 17688 2556 17740
rect 2688 17688 2740 17740
rect 2964 17688 3016 17740
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 6184 17688 6236 17740
rect 7380 17688 7432 17740
rect 8208 17731 8260 17740
rect 8208 17697 8217 17731
rect 8217 17697 8251 17731
rect 8251 17697 8260 17731
rect 8208 17688 8260 17697
rect 5724 17663 5776 17672
rect 4620 17552 4672 17604
rect 4896 17552 4948 17604
rect 3332 17484 3384 17536
rect 3516 17484 3568 17536
rect 3700 17527 3752 17536
rect 3700 17493 3709 17527
rect 3709 17493 3743 17527
rect 3743 17493 3752 17527
rect 3700 17484 3752 17493
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 11612 17620 11664 17672
rect 12164 17663 12216 17672
rect 7012 17552 7064 17604
rect 8668 17552 8720 17604
rect 11428 17552 11480 17604
rect 12164 17629 12180 17663
rect 12180 17629 12214 17663
rect 12214 17629 12216 17663
rect 12164 17620 12216 17629
rect 13820 17688 13872 17740
rect 15844 17688 15896 17740
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 16488 17688 16540 17740
rect 16580 17688 16632 17740
rect 13360 17620 13412 17672
rect 13176 17552 13228 17604
rect 5908 17484 5960 17536
rect 8024 17484 8076 17536
rect 10784 17484 10836 17536
rect 11704 17484 11756 17536
rect 13820 17484 13872 17536
rect 4947 17382 4999 17434
rect 5011 17382 5063 17434
rect 5075 17382 5127 17434
rect 5139 17382 5191 17434
rect 12878 17382 12930 17434
rect 12942 17382 12994 17434
rect 13006 17382 13058 17434
rect 13070 17382 13122 17434
rect 20808 17382 20860 17434
rect 20872 17382 20924 17434
rect 20936 17382 20988 17434
rect 21000 17382 21052 17434
rect 2228 17280 2280 17332
rect 2596 17212 2648 17264
rect 4344 17280 4396 17332
rect 10692 17280 10744 17332
rect 11612 17280 11664 17332
rect 16028 17280 16080 17332
rect 4712 17212 4764 17264
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 2136 17076 2188 17128
rect 2688 17076 2740 17128
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 7472 17212 7524 17264
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 7748 17187 7800 17196
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 7472 17076 7524 17128
rect 10140 17076 10192 17128
rect 10324 17076 10376 17128
rect 10600 17076 10652 17128
rect 12440 17144 12492 17196
rect 12532 17144 12584 17196
rect 17500 17144 17552 17196
rect 19064 17144 19116 17196
rect 12624 17119 12676 17128
rect 8024 17008 8076 17060
rect 9864 17051 9916 17060
rect 9864 17017 9873 17051
rect 9873 17017 9907 17051
rect 9907 17017 9916 17051
rect 9864 17008 9916 17017
rect 8300 16940 8352 16992
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 13728 17076 13780 17128
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 15568 17119 15620 17128
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 15568 17085 15577 17119
rect 15577 17085 15611 17119
rect 15611 17085 15620 17119
rect 15568 17076 15620 17085
rect 15844 17076 15896 17128
rect 12440 17008 12492 17017
rect 16028 17008 16080 17060
rect 18236 17076 18288 17128
rect 12164 16940 12216 16992
rect 15568 16940 15620 16992
rect 17132 16940 17184 16992
rect 18512 16940 18564 16992
rect 8912 16838 8964 16890
rect 8976 16838 9028 16890
rect 9040 16838 9092 16890
rect 9104 16838 9156 16890
rect 16843 16838 16895 16890
rect 16907 16838 16959 16890
rect 16971 16838 17023 16890
rect 17035 16838 17087 16890
rect 5540 16736 5592 16788
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 19064 16736 19116 16788
rect 3792 16668 3844 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 4160 16532 4212 16584
rect 4528 16668 4580 16720
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 11060 16668 11112 16720
rect 11704 16711 11756 16720
rect 6460 16600 6512 16652
rect 7472 16600 7524 16652
rect 9588 16600 9640 16652
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 8576 16575 8628 16584
rect 4344 16464 4396 16516
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 10048 16532 10100 16584
rect 10416 16600 10468 16652
rect 11152 16600 11204 16652
rect 11704 16677 11713 16711
rect 11713 16677 11747 16711
rect 11747 16677 11756 16711
rect 11704 16668 11756 16677
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 13728 16600 13780 16652
rect 13452 16532 13504 16584
rect 15476 16600 15528 16652
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 16120 16600 16172 16652
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 8300 16464 8352 16516
rect 15568 16532 15620 16584
rect 14648 16464 14700 16516
rect 15108 16464 15160 16516
rect 3976 16396 4028 16448
rect 8392 16396 8444 16448
rect 8576 16396 8628 16448
rect 10968 16396 11020 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14280 16396 14332 16448
rect 14556 16396 14608 16448
rect 16948 16396 17000 16448
rect 18420 16396 18472 16448
rect 4947 16294 4999 16346
rect 5011 16294 5063 16346
rect 5075 16294 5127 16346
rect 5139 16294 5191 16346
rect 12878 16294 12930 16346
rect 12942 16294 12994 16346
rect 13006 16294 13058 16346
rect 13070 16294 13122 16346
rect 20808 16294 20860 16346
rect 20872 16294 20924 16346
rect 20936 16294 20988 16346
rect 21000 16294 21052 16346
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 8208 16192 8260 16244
rect 12256 16192 12308 16244
rect 16120 16192 16172 16244
rect 17132 16192 17184 16244
rect 17592 16192 17644 16244
rect 19248 16192 19300 16244
rect 2596 16124 2648 16176
rect 3976 16099 4028 16108
rect 3976 16065 3985 16099
rect 3985 16065 4019 16099
rect 4019 16065 4028 16099
rect 3976 16056 4028 16065
rect 4160 16056 4212 16108
rect 6184 16056 6236 16108
rect 6828 16056 6880 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 9864 16056 9916 16108
rect 12164 16056 12216 16108
rect 15016 16099 15068 16108
rect 2320 16031 2372 16040
rect 2320 15997 2326 16031
rect 2326 15997 2372 16031
rect 2320 15988 2372 15997
rect 2504 16031 2556 16040
rect 2504 15997 2518 16031
rect 2518 15997 2556 16031
rect 2504 15988 2556 15997
rect 3056 15988 3108 16040
rect 3700 16031 3752 16040
rect 3700 15997 3709 16031
rect 3709 15997 3743 16031
rect 3743 15997 3752 16031
rect 3700 15988 3752 15997
rect 6368 16031 6420 16040
rect 6368 15997 6377 16031
rect 6377 15997 6411 16031
rect 6411 15997 6420 16031
rect 6368 15988 6420 15997
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7104 15988 7156 16040
rect 2044 15920 2096 15972
rect 2964 15920 3016 15972
rect 7380 15920 7432 15972
rect 9772 15988 9824 16040
rect 12256 15988 12308 16040
rect 13544 15988 13596 16040
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 15660 15988 15712 16040
rect 16212 16056 16264 16108
rect 17500 16056 17552 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 18696 15988 18748 16040
rect 13452 15920 13504 15972
rect 16580 15920 16632 15972
rect 13176 15852 13228 15904
rect 8912 15750 8964 15802
rect 8976 15750 9028 15802
rect 9040 15750 9092 15802
rect 9104 15750 9156 15802
rect 16843 15750 16895 15802
rect 16907 15750 16959 15802
rect 16971 15750 17023 15802
rect 17035 15750 17087 15802
rect 1676 15580 1728 15632
rect 14464 15648 14516 15700
rect 14648 15648 14700 15700
rect 15476 15648 15528 15700
rect 17960 15691 18012 15700
rect 17960 15657 17969 15691
rect 17969 15657 18003 15691
rect 18003 15657 18012 15691
rect 17960 15648 18012 15657
rect 5264 15580 5316 15632
rect 6644 15580 6696 15632
rect 2504 15512 2556 15564
rect 2688 15512 2740 15564
rect 3608 15512 3660 15564
rect 4068 15512 4120 15564
rect 2412 15444 2464 15496
rect 4160 15444 4212 15496
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 7196 15512 7248 15564
rect 7840 15512 7892 15564
rect 8392 15512 8444 15564
rect 9220 15512 9272 15564
rect 6644 15444 6696 15496
rect 8208 15444 8260 15496
rect 2964 15376 3016 15428
rect 9772 15512 9824 15564
rect 12164 15512 12216 15564
rect 12532 15444 12584 15496
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 14556 15580 14608 15632
rect 15384 15580 15436 15632
rect 15476 15512 15528 15564
rect 15660 15512 15712 15564
rect 16304 15555 16356 15564
rect 16304 15521 16313 15555
rect 16313 15521 16347 15555
rect 16347 15521 16356 15555
rect 16304 15512 16356 15521
rect 16672 15512 16724 15564
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 9220 15308 9272 15360
rect 12440 15308 12492 15360
rect 18144 15444 18196 15496
rect 18420 15444 18472 15496
rect 17500 15419 17552 15428
rect 17500 15385 17524 15419
rect 17524 15385 17552 15419
rect 17500 15376 17552 15385
rect 17592 15351 17644 15360
rect 17592 15317 17601 15351
rect 17601 15317 17635 15351
rect 17635 15317 17644 15351
rect 17592 15308 17644 15317
rect 4947 15206 4999 15258
rect 5011 15206 5063 15258
rect 5075 15206 5127 15258
rect 5139 15206 5191 15258
rect 12878 15206 12930 15258
rect 12942 15206 12994 15258
rect 13006 15206 13058 15258
rect 13070 15206 13122 15258
rect 20808 15206 20860 15258
rect 20872 15206 20924 15258
rect 20936 15206 20988 15258
rect 21000 15206 21052 15258
rect 5264 15104 5316 15156
rect 5448 15104 5500 15156
rect 8208 15104 8260 15156
rect 3608 15036 3660 15088
rect 2688 14968 2740 15020
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 8576 15036 8628 15088
rect 13544 15079 13596 15088
rect 13544 15045 13553 15079
rect 13553 15045 13587 15079
rect 13587 15045 13596 15079
rect 13544 15036 13596 15045
rect 2504 14900 2556 14952
rect 2780 14900 2832 14952
rect 1768 14832 1820 14884
rect 2596 14832 2648 14884
rect 3976 14900 4028 14952
rect 4344 14900 4396 14952
rect 4620 14900 4672 14952
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 5908 14900 5960 14952
rect 8576 14900 8628 14952
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 10048 14900 10100 14952
rect 10416 14900 10468 14952
rect 10876 14900 10928 14952
rect 12164 14900 12216 14952
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 13636 14968 13688 15020
rect 13268 14900 13320 14952
rect 15752 15036 15804 15088
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 15752 14900 15804 14952
rect 16580 14900 16632 14952
rect 17960 14900 18012 14952
rect 4068 14832 4120 14884
rect 9680 14832 9732 14884
rect 3240 14764 3292 14816
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 11428 14807 11480 14816
rect 11428 14773 11437 14807
rect 11437 14773 11471 14807
rect 11471 14773 11480 14807
rect 11428 14764 11480 14773
rect 11704 14764 11756 14816
rect 14648 14764 14700 14816
rect 15568 14764 15620 14816
rect 18052 14764 18104 14816
rect 8912 14662 8964 14714
rect 8976 14662 9028 14714
rect 9040 14662 9092 14714
rect 9104 14662 9156 14714
rect 16843 14662 16895 14714
rect 16907 14662 16959 14714
rect 16971 14662 17023 14714
rect 17035 14662 17087 14714
rect 11428 14560 11480 14612
rect 11888 14560 11940 14612
rect 2228 14492 2280 14544
rect 4068 14492 4120 14544
rect 8576 14535 8628 14544
rect 8576 14501 8585 14535
rect 8585 14501 8619 14535
rect 8619 14501 8628 14535
rect 8576 14492 8628 14501
rect 8852 14492 8904 14544
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 7932 14424 7984 14476
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 11244 14467 11296 14476
rect 2412 14356 2464 14408
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 2964 14356 3016 14408
rect 3700 14356 3752 14408
rect 5264 14356 5316 14408
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 5908 14288 5960 14340
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 11428 14424 11480 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 12164 14492 12216 14544
rect 12900 14492 12952 14544
rect 13728 14492 13780 14544
rect 15200 14560 15252 14612
rect 15752 14560 15804 14612
rect 15660 14492 15712 14544
rect 12256 14467 12308 14476
rect 12256 14433 12265 14467
rect 12265 14433 12299 14467
rect 12299 14433 12308 14467
rect 12256 14424 12308 14433
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 12900 14288 12952 14340
rect 16856 14424 16908 14476
rect 15292 14356 15344 14408
rect 15844 14356 15896 14408
rect 17132 14356 17184 14408
rect 1676 14220 1728 14272
rect 2688 14220 2740 14272
rect 5448 14220 5500 14272
rect 6828 14220 6880 14272
rect 7932 14220 7984 14272
rect 9956 14220 10008 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 13912 14220 13964 14272
rect 17868 14220 17920 14272
rect 17960 14220 18012 14272
rect 18144 14263 18196 14272
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 4947 14118 4999 14170
rect 5011 14118 5063 14170
rect 5075 14118 5127 14170
rect 5139 14118 5191 14170
rect 12878 14118 12930 14170
rect 12942 14118 12994 14170
rect 13006 14118 13058 14170
rect 13070 14118 13122 14170
rect 20808 14118 20860 14170
rect 20872 14118 20924 14170
rect 20936 14118 20988 14170
rect 21000 14118 21052 14170
rect 3976 14016 4028 14068
rect 7012 14016 7064 14068
rect 9956 14016 10008 14068
rect 11244 14016 11296 14068
rect 11704 14016 11756 14068
rect 11980 14016 12032 14068
rect 12348 14016 12400 14068
rect 7472 13948 7524 14000
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 4068 13880 4120 13932
rect 2780 13812 2832 13864
rect 3976 13812 4028 13864
rect 5908 13880 5960 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 7932 13880 7984 13932
rect 6552 13812 6604 13864
rect 7748 13812 7800 13864
rect 9220 13948 9272 14000
rect 12532 13948 12584 14000
rect 13360 13948 13412 14000
rect 17868 13948 17920 14000
rect 15568 13923 15620 13932
rect 9772 13812 9824 13864
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15660 13880 15712 13932
rect 11336 13812 11388 13864
rect 11428 13812 11480 13864
rect 8208 13744 8260 13796
rect 8852 13744 8904 13796
rect 9588 13787 9640 13796
rect 9588 13753 9597 13787
rect 9597 13753 9631 13787
rect 9631 13753 9640 13787
rect 9588 13744 9640 13753
rect 13176 13812 13228 13864
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 15384 13744 15436 13796
rect 11796 13676 11848 13728
rect 12164 13676 12216 13728
rect 13728 13676 13780 13728
rect 14372 13676 14424 13728
rect 16856 13812 16908 13864
rect 17868 13812 17920 13864
rect 8912 13574 8964 13626
rect 8976 13574 9028 13626
rect 9040 13574 9092 13626
rect 9104 13574 9156 13626
rect 16843 13574 16895 13626
rect 16907 13574 16959 13626
rect 16971 13574 17023 13626
rect 17035 13574 17087 13626
rect 2504 13472 2556 13524
rect 6092 13515 6144 13524
rect 5264 13404 5316 13456
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 13636 13472 13688 13524
rect 11888 13404 11940 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 5540 13336 5592 13388
rect 6644 13379 6696 13388
rect 6644 13345 6653 13379
rect 6653 13345 6687 13379
rect 6687 13345 6696 13379
rect 6644 13336 6696 13345
rect 7012 13379 7064 13388
rect 7012 13345 7026 13379
rect 7026 13345 7064 13379
rect 7012 13336 7064 13345
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 5816 13268 5868 13320
rect 6184 13268 6236 13320
rect 7472 13336 7524 13388
rect 9588 13336 9640 13388
rect 13636 13336 13688 13388
rect 7840 13268 7892 13320
rect 8116 13268 8168 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9220 13268 9272 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9864 13268 9916 13320
rect 18512 13472 18564 13524
rect 15292 13447 15344 13456
rect 15292 13413 15301 13447
rect 15301 13413 15335 13447
rect 15335 13413 15344 13447
rect 15292 13404 15344 13413
rect 16120 13404 16172 13456
rect 16488 13404 16540 13456
rect 17132 13404 17184 13456
rect 16212 13336 16264 13388
rect 18052 13404 18104 13456
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17960 13379 18012 13388
rect 17684 13336 17736 13345
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 18972 13336 19024 13388
rect 5540 13200 5592 13252
rect 4712 13132 4764 13184
rect 7840 13132 7892 13184
rect 8392 13132 8444 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 15752 13268 15804 13320
rect 13176 13200 13228 13252
rect 16304 13200 16356 13252
rect 13636 13132 13688 13184
rect 15384 13132 15436 13184
rect 15476 13132 15528 13184
rect 15660 13132 15712 13184
rect 4947 13030 4999 13082
rect 5011 13030 5063 13082
rect 5075 13030 5127 13082
rect 5139 13030 5191 13082
rect 12878 13030 12930 13082
rect 12942 13030 12994 13082
rect 13006 13030 13058 13082
rect 13070 13030 13122 13082
rect 20808 13030 20860 13082
rect 20872 13030 20924 13082
rect 20936 13030 20988 13082
rect 21000 13030 21052 13082
rect 6368 12928 6420 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 13452 12928 13504 12980
rect 13728 12928 13780 12980
rect 3332 12835 3384 12844
rect 3056 12724 3108 12776
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 9864 12860 9916 12912
rect 14372 12903 14424 12912
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 16488 12860 16540 12912
rect 4252 12792 4304 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5632 12792 5684 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 2504 12656 2556 12708
rect 2780 12699 2832 12708
rect 2780 12665 2789 12699
rect 2789 12665 2823 12699
rect 2823 12665 2832 12699
rect 2780 12656 2832 12665
rect 4160 12656 4212 12708
rect 5264 12656 5316 12708
rect 8944 12724 8996 12776
rect 10048 12792 10100 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 8852 12656 8904 12708
rect 10784 12724 10836 12776
rect 11336 12724 11388 12776
rect 12440 12724 12492 12776
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 10416 12656 10468 12708
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 16672 12724 16724 12776
rect 17132 12724 17184 12776
rect 8484 12588 8536 12640
rect 18328 12656 18380 12708
rect 8912 12486 8964 12538
rect 8976 12486 9028 12538
rect 9040 12486 9092 12538
rect 9104 12486 9156 12538
rect 16843 12486 16895 12538
rect 16907 12486 16959 12538
rect 16971 12486 17023 12538
rect 17035 12486 17087 12538
rect 2228 12384 2280 12436
rect 2320 12384 2372 12436
rect 2044 12316 2096 12368
rect 3424 12316 3476 12368
rect 4528 12316 4580 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 6644 12316 6696 12368
rect 6920 12316 6972 12368
rect 7012 12248 7064 12300
rect 7932 12248 7984 12300
rect 8484 12248 8536 12300
rect 8668 12248 8720 12300
rect 2780 12180 2832 12232
rect 5724 12180 5776 12232
rect 7656 12180 7708 12232
rect 7932 12112 7984 12164
rect 8484 12155 8536 12164
rect 8484 12121 8493 12155
rect 8493 12121 8527 12155
rect 8527 12121 8536 12155
rect 8484 12112 8536 12121
rect 1400 12044 1452 12096
rect 2596 12044 2648 12096
rect 5448 12044 5500 12096
rect 9588 12044 9640 12096
rect 10968 12316 11020 12368
rect 12532 12316 12584 12368
rect 13268 12384 13320 12436
rect 18328 12384 18380 12436
rect 11060 12248 11112 12300
rect 12348 12248 12400 12300
rect 13360 12248 13412 12300
rect 13912 12248 13964 12300
rect 17132 12248 17184 12300
rect 17868 12248 17920 12300
rect 18972 12291 19024 12300
rect 18972 12257 18981 12291
rect 18981 12257 19015 12291
rect 19015 12257 19024 12291
rect 18972 12248 19024 12257
rect 11520 12180 11572 12232
rect 16672 12180 16724 12232
rect 17684 12180 17736 12232
rect 13728 12112 13780 12164
rect 17592 12112 17644 12164
rect 17960 12112 18012 12164
rect 10876 12044 10928 12096
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 12256 12044 12308 12053
rect 18052 12044 18104 12096
rect 4947 11942 4999 11994
rect 5011 11942 5063 11994
rect 5075 11942 5127 11994
rect 5139 11942 5191 11994
rect 12878 11942 12930 11994
rect 12942 11942 12994 11994
rect 13006 11942 13058 11994
rect 13070 11942 13122 11994
rect 20808 11942 20860 11994
rect 20872 11942 20924 11994
rect 20936 11942 20988 11994
rect 21000 11942 21052 11994
rect 10876 11840 10928 11892
rect 11060 11840 11112 11892
rect 4068 11772 4120 11824
rect 6552 11772 6604 11824
rect 6828 11772 6880 11824
rect 9588 11772 9640 11824
rect 12348 11772 12400 11824
rect 17316 11840 17368 11892
rect 18972 11840 19024 11892
rect 16580 11772 16632 11824
rect 17224 11772 17276 11824
rect 17592 11772 17644 11824
rect 2044 11704 2096 11756
rect 6644 11704 6696 11756
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 10416 11704 10468 11756
rect 10968 11704 11020 11756
rect 11152 11704 11204 11756
rect 11888 11704 11940 11756
rect 17132 11704 17184 11756
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 1676 11568 1728 11620
rect 2320 11636 2372 11688
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 6368 11636 6420 11688
rect 2412 11568 2464 11620
rect 3608 11568 3660 11620
rect 4896 11568 4948 11620
rect 6092 11568 6144 11620
rect 7012 11636 7064 11688
rect 7840 11636 7892 11688
rect 12164 11636 12216 11688
rect 10784 11568 10836 11620
rect 12532 11636 12584 11688
rect 14004 11636 14056 11688
rect 14464 11636 14516 11688
rect 16580 11636 16632 11688
rect 17868 11636 17920 11688
rect 16856 11568 16908 11620
rect 17500 11568 17552 11620
rect 6552 11500 6604 11552
rect 7932 11500 7984 11552
rect 12440 11500 12492 11552
rect 12532 11500 12584 11552
rect 13360 11500 13412 11552
rect 16488 11500 16540 11552
rect 18972 11568 19024 11620
rect 8912 11398 8964 11450
rect 8976 11398 9028 11450
rect 9040 11398 9092 11450
rect 9104 11398 9156 11450
rect 16843 11398 16895 11450
rect 16907 11398 16959 11450
rect 16971 11398 17023 11450
rect 17035 11398 17087 11450
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 6736 11339 6788 11348
rect 2780 11296 2832 11305
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 6828 11296 6880 11348
rect 5448 11228 5500 11280
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 4252 11160 4304 11212
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 6920 11160 6972 11212
rect 1584 11092 1636 11144
rect 1860 11092 1912 11144
rect 4160 11092 4212 11144
rect 4804 11092 4856 11144
rect 8484 11160 8536 11212
rect 11520 11160 11572 11212
rect 13360 11160 13412 11212
rect 15568 11296 15620 11348
rect 17868 11296 17920 11348
rect 17132 11228 17184 11280
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 8116 11092 8168 11144
rect 9772 11092 9824 11144
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 12716 11092 12768 11144
rect 13636 11092 13688 11144
rect 14004 11092 14056 11144
rect 7840 11024 7892 11076
rect 12164 11067 12216 11076
rect 12164 11033 12173 11067
rect 12173 11033 12207 11067
rect 12207 11033 12216 11067
rect 12164 11024 12216 11033
rect 12440 11024 12492 11076
rect 6184 10956 6236 11008
rect 11244 10956 11296 11008
rect 11980 10956 12032 11008
rect 14096 11024 14148 11076
rect 14740 11024 14792 11076
rect 16028 10956 16080 11008
rect 16304 10956 16356 11008
rect 18420 10956 18472 11008
rect 4947 10854 4999 10906
rect 5011 10854 5063 10906
rect 5075 10854 5127 10906
rect 5139 10854 5191 10906
rect 12878 10854 12930 10906
rect 12942 10854 12994 10906
rect 13006 10854 13058 10906
rect 13070 10854 13122 10906
rect 20808 10854 20860 10906
rect 20872 10854 20924 10906
rect 20936 10854 20988 10906
rect 21000 10854 21052 10906
rect 3700 10752 3752 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 5540 10752 5592 10804
rect 11060 10752 11112 10804
rect 1860 10616 1912 10668
rect 4160 10659 4212 10668
rect 3148 10548 3200 10600
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 6552 10591 6604 10600
rect 3240 10480 3292 10532
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 7380 10684 7432 10736
rect 11244 10684 11296 10736
rect 11704 10616 11756 10668
rect 11796 10616 11848 10668
rect 14464 10684 14516 10736
rect 15568 10752 15620 10804
rect 16396 10752 16448 10804
rect 16672 10752 16724 10804
rect 17592 10752 17644 10804
rect 7656 10548 7708 10600
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 7932 10480 7984 10532
rect 10784 10548 10836 10600
rect 11520 10591 11572 10600
rect 7012 10412 7064 10464
rect 7380 10412 7432 10464
rect 9956 10412 10008 10464
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12532 10548 12584 10600
rect 13268 10548 13320 10600
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 15292 10548 15344 10600
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16396 10591 16448 10600
rect 16120 10548 16172 10557
rect 16396 10557 16405 10591
rect 16405 10557 16439 10591
rect 16439 10557 16448 10591
rect 16396 10548 16448 10557
rect 16488 10591 16540 10600
rect 16488 10557 16497 10591
rect 16497 10557 16531 10591
rect 16531 10557 16540 10591
rect 16488 10548 16540 10557
rect 18236 10548 18288 10600
rect 18420 10548 18472 10600
rect 13728 10412 13780 10464
rect 13912 10412 13964 10464
rect 8912 10310 8964 10362
rect 8976 10310 9028 10362
rect 9040 10310 9092 10362
rect 9104 10310 9156 10362
rect 16843 10310 16895 10362
rect 16907 10310 16959 10362
rect 16971 10310 17023 10362
rect 17035 10310 17087 10362
rect 2412 10208 2464 10260
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 3700 10004 3752 10056
rect 2044 9979 2096 9988
rect 2044 9945 2053 9979
rect 2053 9945 2087 9979
rect 2087 9945 2096 9979
rect 2044 9936 2096 9945
rect 11336 10208 11388 10260
rect 13636 10208 13688 10260
rect 13912 10208 13964 10260
rect 7012 10183 7064 10192
rect 7012 10149 7021 10183
rect 7021 10149 7055 10183
rect 7055 10149 7064 10183
rect 7012 10140 7064 10149
rect 7104 10140 7156 10192
rect 7472 10140 7524 10192
rect 16028 10208 16080 10260
rect 16304 10140 16356 10192
rect 16488 10183 16540 10192
rect 16488 10149 16497 10183
rect 16497 10149 16531 10183
rect 16531 10149 16540 10183
rect 16488 10140 16540 10149
rect 17960 10140 18012 10192
rect 6644 10072 6696 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 11060 10072 11112 10124
rect 12256 10072 12308 10124
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 7012 10004 7064 10056
rect 7932 10004 7984 10056
rect 11980 10004 12032 10056
rect 12440 10004 12492 10056
rect 15200 10072 15252 10124
rect 16672 10115 16724 10124
rect 16672 10081 16678 10115
rect 16678 10081 16724 10115
rect 16672 10072 16724 10081
rect 16212 10004 16264 10056
rect 16396 10004 16448 10056
rect 16488 10004 16540 10056
rect 18972 10072 19024 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 17224 10004 17276 10056
rect 7564 9868 7616 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 13268 9936 13320 9988
rect 10140 9868 10192 9920
rect 11520 9868 11572 9920
rect 12348 9868 12400 9920
rect 14004 9868 14056 9920
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 17316 9936 17368 9988
rect 18236 9936 18288 9988
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 21180 9868 21232 9920
rect 4947 9766 4999 9818
rect 5011 9766 5063 9818
rect 5075 9766 5127 9818
rect 5139 9766 5191 9818
rect 12878 9766 12930 9818
rect 12942 9766 12994 9818
rect 13006 9766 13058 9818
rect 13070 9766 13122 9818
rect 20808 9766 20860 9818
rect 20872 9766 20924 9818
rect 20936 9766 20988 9818
rect 21000 9766 21052 9818
rect 3056 9596 3108 9648
rect 5172 9596 5224 9648
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 5816 9528 5868 9580
rect 6276 9528 6328 9580
rect 10784 9664 10836 9716
rect 18144 9664 18196 9716
rect 10968 9596 11020 9648
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 4896 9460 4948 9512
rect 5080 9460 5132 9512
rect 6184 9460 6236 9512
rect 7564 9460 7616 9512
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 7472 9392 7524 9444
rect 8576 9460 8628 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 10416 9460 10468 9512
rect 3424 9324 3476 9376
rect 3884 9324 3936 9376
rect 5448 9324 5500 9376
rect 7840 9324 7892 9376
rect 10968 9324 11020 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 11888 9528 11940 9580
rect 13728 9528 13780 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 11980 9460 12032 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 16304 9528 16356 9580
rect 17224 9460 17276 9512
rect 18144 9460 18196 9512
rect 15476 9392 15528 9444
rect 16304 9324 16356 9376
rect 16580 9324 16632 9376
rect 18236 9392 18288 9444
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 8912 9222 8964 9274
rect 8976 9222 9028 9274
rect 9040 9222 9092 9274
rect 9104 9222 9156 9274
rect 16843 9222 16895 9274
rect 16907 9222 16959 9274
rect 16971 9222 17023 9274
rect 17035 9222 17087 9274
rect 2136 9120 2188 9172
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 3884 9052 3936 9104
rect 5356 9052 5408 9104
rect 4160 8984 4212 9036
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 5448 8984 5500 9036
rect 8116 9052 8168 9104
rect 8300 9052 8352 9104
rect 9220 9052 9272 9104
rect 12440 9052 12492 9104
rect 6920 8984 6972 9036
rect 8024 8984 8076 9036
rect 2872 8916 2924 8968
rect 4068 8848 4120 8900
rect 6736 8916 6788 8968
rect 11060 8984 11112 9036
rect 12348 8984 12400 9036
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 13820 8984 13872 9036
rect 14556 9052 14608 9104
rect 17316 9052 17368 9104
rect 11152 8916 11204 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12532 8916 12584 8968
rect 18144 8984 18196 9036
rect 14004 8916 14056 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 17224 8916 17276 8968
rect 6460 8848 6512 8900
rect 2964 8780 3016 8832
rect 10784 8848 10836 8900
rect 17500 8848 17552 8900
rect 9680 8780 9732 8832
rect 12440 8780 12492 8832
rect 13268 8780 13320 8832
rect 16396 8780 16448 8832
rect 4947 8678 4999 8730
rect 5011 8678 5063 8730
rect 5075 8678 5127 8730
rect 5139 8678 5191 8730
rect 12878 8678 12930 8730
rect 12942 8678 12994 8730
rect 13006 8678 13058 8730
rect 13070 8678 13122 8730
rect 20808 8678 20860 8730
rect 20872 8678 20924 8730
rect 20936 8678 20988 8730
rect 21000 8678 21052 8730
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 7472 8576 7524 8628
rect 2320 8508 2372 8560
rect 2688 8508 2740 8560
rect 2688 8372 2740 8424
rect 2964 8415 3016 8424
rect 1676 8304 1728 8356
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 5356 8508 5408 8560
rect 6920 8508 6972 8560
rect 7196 8508 7248 8560
rect 10968 8551 11020 8560
rect 4436 8440 4488 8492
rect 4252 8372 4304 8424
rect 5540 8372 5592 8424
rect 6368 8372 6420 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 11336 8440 11388 8492
rect 11980 8440 12032 8492
rect 4528 8304 4580 8356
rect 9772 8304 9824 8356
rect 11244 8372 11296 8424
rect 12348 8372 12400 8424
rect 12716 8347 12768 8356
rect 388 8236 440 8288
rect 6092 8236 6144 8288
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 10876 8236 10928 8288
rect 11060 8236 11112 8288
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 13268 8576 13320 8628
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 13820 8508 13872 8560
rect 14004 8508 14056 8560
rect 13268 8440 13320 8492
rect 13728 8440 13780 8492
rect 17224 8508 17276 8560
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14740 8440 14792 8492
rect 20168 8440 20220 8492
rect 13360 8372 13412 8424
rect 14004 8372 14056 8424
rect 14280 8372 14332 8424
rect 14924 8372 14976 8424
rect 17960 8372 18012 8424
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 13268 8236 13320 8288
rect 21180 8304 21232 8356
rect 18144 8279 18196 8288
rect 18144 8245 18153 8279
rect 18153 8245 18187 8279
rect 18187 8245 18196 8279
rect 18144 8236 18196 8245
rect 8912 8134 8964 8186
rect 8976 8134 9028 8186
rect 9040 8134 9092 8186
rect 9104 8134 9156 8186
rect 16843 8134 16895 8186
rect 16907 8134 16959 8186
rect 16971 8134 17023 8186
rect 17035 8134 17087 8186
rect 3976 8032 4028 8084
rect 7380 8032 7432 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 4344 7896 4396 7948
rect 5264 7896 5316 7948
rect 6920 7964 6972 8016
rect 10968 8032 11020 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 12256 8032 12308 8084
rect 12440 8032 12492 8084
rect 12716 8032 12768 8084
rect 13268 8032 13320 8084
rect 6552 7896 6604 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1860 7828 1912 7880
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 4068 7760 4120 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 6736 7692 6788 7744
rect 7104 7760 7156 7812
rect 11520 7964 11572 8016
rect 13636 7964 13688 8016
rect 7564 7896 7616 7948
rect 9220 7896 9272 7948
rect 9588 7896 9640 7948
rect 12716 7896 12768 7948
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13084 7896 13136 7948
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 14556 7964 14608 8016
rect 16304 8007 16356 8016
rect 16304 7973 16313 8007
rect 16313 7973 16347 8007
rect 16347 7973 16356 8007
rect 16304 7964 16356 7973
rect 14372 7896 14424 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 18144 7964 18196 8016
rect 17224 7896 17276 7948
rect 17500 7939 17552 7948
rect 17500 7905 17509 7939
rect 17509 7905 17543 7939
rect 17543 7905 17552 7939
rect 17500 7896 17552 7905
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 14464 7828 14516 7880
rect 16580 7828 16632 7880
rect 8300 7803 8352 7812
rect 8300 7769 8309 7803
rect 8309 7769 8343 7803
rect 8343 7769 8352 7803
rect 8300 7760 8352 7769
rect 11704 7760 11756 7812
rect 11980 7760 12032 7812
rect 12348 7760 12400 7812
rect 12808 7760 12860 7812
rect 16856 7760 16908 7812
rect 14924 7692 14976 7744
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 4947 7590 4999 7642
rect 5011 7590 5063 7642
rect 5075 7590 5127 7642
rect 5139 7590 5191 7642
rect 12878 7590 12930 7642
rect 12942 7590 12994 7642
rect 13006 7590 13058 7642
rect 13070 7590 13122 7642
rect 20808 7590 20860 7642
rect 20872 7590 20924 7642
rect 20936 7590 20988 7642
rect 21000 7590 21052 7642
rect 3792 7488 3844 7540
rect 3976 7488 4028 7540
rect 4528 7488 4580 7540
rect 9496 7488 9548 7540
rect 10048 7488 10100 7540
rect 10692 7488 10744 7540
rect 11704 7488 11756 7540
rect 18420 7488 18472 7540
rect 9680 7420 9732 7472
rect 10508 7420 10560 7472
rect 3700 7284 3752 7336
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 2688 7148 2740 7200
rect 5448 7352 5500 7404
rect 6736 7352 6788 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 11612 7352 11664 7404
rect 12532 7420 12584 7472
rect 13728 7420 13780 7472
rect 16856 7463 16908 7472
rect 16856 7429 16865 7463
rect 16865 7429 16899 7463
rect 16899 7429 16908 7463
rect 16856 7420 16908 7429
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13176 7352 13228 7404
rect 14188 7352 14240 7404
rect 4528 7284 4580 7336
rect 5264 7284 5316 7336
rect 5080 7259 5132 7268
rect 5080 7225 5089 7259
rect 5089 7225 5123 7259
rect 5123 7225 5132 7259
rect 5080 7216 5132 7225
rect 10968 7216 11020 7268
rect 6920 7148 6972 7200
rect 11060 7148 11112 7200
rect 14280 7327 14332 7336
rect 12440 7259 12492 7268
rect 12440 7225 12449 7259
rect 12449 7225 12483 7259
rect 12483 7225 12492 7259
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 19064 7352 19116 7404
rect 17500 7284 17552 7336
rect 12440 7216 12492 7225
rect 12808 7148 12860 7200
rect 13728 7148 13780 7200
rect 16580 7148 16632 7200
rect 17316 7216 17368 7268
rect 17132 7148 17184 7200
rect 8912 7046 8964 7098
rect 8976 7046 9028 7098
rect 9040 7046 9092 7098
rect 9104 7046 9156 7098
rect 16843 7046 16895 7098
rect 16907 7046 16959 7098
rect 16971 7046 17023 7098
rect 17035 7046 17087 7098
rect 4252 6944 4304 6996
rect 3700 6876 3752 6928
rect 4160 6876 4212 6928
rect 4436 6919 4488 6928
rect 4436 6885 4445 6919
rect 4445 6885 4479 6919
rect 4479 6885 4488 6919
rect 4436 6876 4488 6885
rect 1676 6740 1728 6792
rect 2688 6672 2740 6724
rect 2964 6808 3016 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4160 6740 4212 6792
rect 5448 6876 5500 6928
rect 5908 6876 5960 6928
rect 6828 6876 6880 6928
rect 5540 6808 5592 6860
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 6736 6808 6788 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 5908 6740 5960 6792
rect 7932 6740 7984 6792
rect 9956 6740 10008 6792
rect 2964 6672 3016 6724
rect 5080 6672 5132 6724
rect 12164 6944 12216 6996
rect 10416 6876 10468 6928
rect 11060 6808 11112 6860
rect 11612 6876 11664 6928
rect 12532 6944 12584 6996
rect 12808 6944 12860 6996
rect 14280 6944 14332 6996
rect 17500 6944 17552 6996
rect 12716 6876 12768 6928
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 3056 6604 3108 6656
rect 3516 6604 3568 6656
rect 5448 6604 5500 6656
rect 12532 6808 12584 6860
rect 13360 6808 13412 6860
rect 17132 6876 17184 6928
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 13176 6740 13228 6792
rect 13912 6740 13964 6792
rect 14188 6740 14240 6792
rect 16120 6740 16172 6792
rect 16580 6740 16632 6792
rect 17408 6808 17460 6860
rect 18972 6740 19024 6792
rect 11336 6672 11388 6724
rect 13912 6604 13964 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 4947 6502 4999 6554
rect 5011 6502 5063 6554
rect 5075 6502 5127 6554
rect 5139 6502 5191 6554
rect 12878 6502 12930 6554
rect 12942 6502 12994 6554
rect 13006 6502 13058 6554
rect 13070 6502 13122 6554
rect 20808 6502 20860 6554
rect 20872 6502 20924 6554
rect 20936 6502 20988 6554
rect 21000 6502 21052 6554
rect 9956 6400 10008 6452
rect 11612 6400 11664 6452
rect 11888 6400 11940 6452
rect 13176 6400 13228 6452
rect 13268 6400 13320 6452
rect 15200 6400 15252 6452
rect 16580 6443 16632 6452
rect 16580 6409 16589 6443
rect 16589 6409 16623 6443
rect 16623 6409 16632 6443
rect 16580 6400 16632 6409
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 4252 6332 4304 6384
rect 7932 6375 7984 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 4436 6264 4488 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 1768 6196 1820 6248
rect 4252 6196 4304 6248
rect 4988 6196 5040 6248
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 7932 6332 7984 6341
rect 10692 6332 10744 6384
rect 5632 6264 5684 6316
rect 6092 6264 6144 6316
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 7012 6239 7064 6248
rect 7012 6205 7021 6239
rect 7021 6205 7055 6239
rect 7055 6205 7064 6239
rect 7012 6196 7064 6205
rect 7104 6196 7156 6248
rect 2412 6128 2464 6180
rect 6920 6128 6972 6180
rect 9864 6196 9916 6248
rect 11152 6264 11204 6316
rect 13360 6264 13412 6316
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 14280 6264 14332 6316
rect 15384 6264 15436 6316
rect 10784 6239 10836 6248
rect 9956 6128 10008 6180
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 13912 6239 13964 6248
rect 13452 6128 13504 6180
rect 4436 6060 4488 6112
rect 4528 6060 4580 6112
rect 4988 6060 5040 6112
rect 7472 6060 7524 6112
rect 11060 6060 11112 6112
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 15108 6196 15160 6248
rect 15384 6060 15436 6112
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 8912 5958 8964 6010
rect 8976 5958 9028 6010
rect 9040 5958 9092 6010
rect 9104 5958 9156 6010
rect 16843 5958 16895 6010
rect 16907 5958 16959 6010
rect 16971 5958 17023 6010
rect 17035 5958 17087 6010
rect 3056 5899 3108 5908
rect 3056 5865 3065 5899
rect 3065 5865 3099 5899
rect 3099 5865 3108 5899
rect 3056 5856 3108 5865
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 9588 5856 9640 5908
rect 10968 5856 11020 5908
rect 11060 5856 11112 5908
rect 18144 5856 18196 5908
rect 4436 5831 4488 5840
rect 4436 5797 4445 5831
rect 4445 5797 4479 5831
rect 4479 5797 4488 5831
rect 4436 5788 4488 5797
rect 4804 5831 4856 5840
rect 4804 5797 4813 5831
rect 4813 5797 4847 5831
rect 4847 5797 4856 5831
rect 4804 5788 4856 5797
rect 5356 5788 5408 5840
rect 6368 5831 6420 5840
rect 6368 5797 6377 5831
rect 6377 5797 6411 5831
rect 6411 5797 6420 5831
rect 6368 5788 6420 5797
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 5908 5763 5960 5772
rect 4344 5720 4396 5729
rect 5908 5729 5917 5763
rect 5917 5729 5951 5763
rect 5951 5729 5960 5763
rect 11152 5788 11204 5840
rect 5908 5720 5960 5729
rect 4436 5652 4488 5704
rect 5448 5652 5500 5704
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 9956 5763 10008 5772
rect 9588 5652 9640 5704
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 13268 5720 13320 5772
rect 13360 5652 13412 5704
rect 5356 5584 5408 5636
rect 5540 5584 5592 5636
rect 15200 5720 15252 5772
rect 14464 5652 14516 5704
rect 14556 5652 14608 5704
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 10416 5516 10468 5568
rect 14004 5584 14056 5636
rect 13360 5516 13412 5568
rect 4947 5414 4999 5466
rect 5011 5414 5063 5466
rect 5075 5414 5127 5466
rect 5139 5414 5191 5466
rect 12878 5414 12930 5466
rect 12942 5414 12994 5466
rect 13006 5414 13058 5466
rect 13070 5414 13122 5466
rect 20808 5414 20860 5466
rect 20872 5414 20924 5466
rect 20936 5414 20988 5466
rect 21000 5414 21052 5466
rect 4344 5312 4396 5364
rect 6828 5312 6880 5364
rect 3700 5244 3752 5296
rect 2964 5176 3016 5228
rect 4160 5244 4212 5296
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 5172 5244 5224 5296
rect 5540 5244 5592 5296
rect 6000 5244 6052 5296
rect 13452 5312 13504 5364
rect 8760 5244 8812 5296
rect 14464 5287 14516 5296
rect 14464 5253 14473 5287
rect 14473 5253 14507 5287
rect 14507 5253 14516 5287
rect 14464 5244 14516 5253
rect 13360 5219 13412 5228
rect 5356 5151 5408 5160
rect 2596 5040 2648 5092
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5264 5040 5316 5092
rect 5540 5108 5592 5160
rect 5908 5040 5960 5092
rect 3884 4972 3936 5024
rect 4344 4972 4396 5024
rect 10140 5040 10192 5092
rect 10324 5108 10376 5160
rect 10692 5151 10744 5160
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 10692 5108 10744 5117
rect 11244 5108 11296 5160
rect 12348 5108 12400 5160
rect 12716 5108 12768 5160
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 11060 5040 11112 5092
rect 10784 4972 10836 5024
rect 12164 4972 12216 5024
rect 18604 5040 18656 5092
rect 8912 4870 8964 4922
rect 8976 4870 9028 4922
rect 9040 4870 9092 4922
rect 9104 4870 9156 4922
rect 16843 4870 16895 4922
rect 16907 4870 16959 4922
rect 16971 4870 17023 4922
rect 17035 4870 17087 4922
rect 9772 4768 9824 4820
rect 11980 4768 12032 4820
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 4160 4632 4212 4684
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 5540 4700 5592 4752
rect 7012 4700 7064 4752
rect 13176 4768 13228 4820
rect 14372 4768 14424 4820
rect 14832 4768 14884 4820
rect 15200 4768 15252 4820
rect 16028 4768 16080 4820
rect 4804 4632 4856 4641
rect 5356 4632 5408 4684
rect 6460 4632 6512 4684
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 6920 4632 6972 4684
rect 8484 4632 8536 4684
rect 13728 4700 13780 4752
rect 14188 4700 14240 4752
rect 13360 4632 13412 4684
rect 13820 4632 13872 4684
rect 23940 4632 23992 4684
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 3792 4564 3844 4616
rect 5632 4564 5684 4616
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 12164 4564 12216 4616
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 23572 4564 23624 4616
rect 24308 4496 24360 4548
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 23296 4471 23348 4480
rect 23296 4437 23305 4471
rect 23305 4437 23339 4471
rect 23339 4437 23348 4471
rect 23296 4428 23348 4437
rect 23388 4428 23440 4480
rect 4947 4326 4999 4378
rect 5011 4326 5063 4378
rect 5075 4326 5127 4378
rect 5139 4326 5191 4378
rect 12878 4326 12930 4378
rect 12942 4326 12994 4378
rect 13006 4326 13058 4378
rect 13070 4326 13122 4378
rect 20808 4326 20860 4378
rect 20872 4326 20924 4378
rect 20936 4326 20988 4378
rect 21000 4326 21052 4378
rect 4160 4224 4212 4276
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 3700 4156 3752 4208
rect 22284 4199 22336 4208
rect 756 4088 808 4140
rect 1492 4088 1544 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2228 4088 2280 4140
rect 3792 4088 3844 4140
rect 22284 4165 22293 4199
rect 22293 4165 22327 4199
rect 22327 4165 22336 4199
rect 22284 4156 22336 4165
rect 112 4020 164 4072
rect 1308 4020 1360 4072
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 6828 4088 6880 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 9864 4088 9916 4140
rect 10416 4088 10468 4140
rect 11244 4088 11296 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13268 4088 13320 4140
rect 14556 4088 14608 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 22192 4131 22244 4140
rect 22192 4097 22198 4131
rect 22198 4097 22244 4131
rect 22192 4088 22244 4097
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 5724 4020 5776 4072
rect 8668 4020 8720 4072
rect 6368 3952 6420 4004
rect 9772 3952 9824 4004
rect 11612 4020 11664 4072
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13360 4020 13412 4072
rect 13728 4020 13780 4072
rect 14924 4020 14976 4072
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 15016 3952 15068 4004
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 9956 3884 10008 3936
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 23388 3952 23440 4004
rect 18512 3884 18564 3936
rect 22192 3884 22244 3936
rect 23020 3884 23072 3936
rect 8912 3782 8964 3834
rect 8976 3782 9028 3834
rect 9040 3782 9092 3834
rect 9104 3782 9156 3834
rect 16843 3782 16895 3834
rect 16907 3782 16959 3834
rect 16971 3782 17023 3834
rect 17035 3782 17087 3834
rect 4804 3680 4856 3732
rect 8208 3680 8260 3732
rect 11152 3680 11204 3732
rect 13084 3680 13136 3732
rect 22376 3680 22428 3732
rect 2688 3587 2740 3596
rect 2688 3553 2697 3587
rect 2697 3553 2731 3587
rect 2731 3553 2740 3587
rect 2688 3544 2740 3553
rect 7288 3612 7340 3664
rect 4068 3544 4120 3596
rect 4528 3544 4580 3596
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 9772 3544 9824 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 16120 3612 16172 3664
rect 22560 3612 22612 3664
rect 12992 3544 13044 3596
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 6828 3476 6880 3528
rect 10876 3476 10928 3528
rect 10968 3476 11020 3528
rect 11336 3476 11388 3528
rect 13820 3544 13872 3596
rect 14004 3544 14056 3596
rect 14556 3544 14608 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 18236 3587 18288 3596
rect 18236 3553 18245 3587
rect 18245 3553 18279 3587
rect 18279 3553 18288 3587
rect 18236 3544 18288 3553
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 16488 3476 16540 3528
rect 18512 3476 18564 3528
rect 17224 3408 17276 3460
rect 17868 3408 17920 3460
rect 22100 3476 22152 3528
rect 21824 3408 21876 3460
rect 1400 3340 1452 3392
rect 3608 3340 3660 3392
rect 6460 3340 6512 3392
rect 10324 3340 10376 3392
rect 12716 3340 12768 3392
rect 15384 3383 15436 3392
rect 15384 3349 15393 3383
rect 15393 3349 15427 3383
rect 15427 3349 15436 3383
rect 15384 3340 15436 3349
rect 16120 3340 16172 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 17500 3340 17552 3392
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 22928 3340 22980 3392
rect 4947 3238 4999 3290
rect 5011 3238 5063 3290
rect 5075 3238 5127 3290
rect 5139 3238 5191 3290
rect 12878 3238 12930 3290
rect 12942 3238 12994 3290
rect 13006 3238 13058 3290
rect 13070 3238 13122 3290
rect 20808 3238 20860 3290
rect 20872 3238 20924 3290
rect 20936 3238 20988 3290
rect 21000 3238 21052 3290
rect 2964 3136 3016 3188
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 5264 3136 5316 3188
rect 7288 3136 7340 3188
rect 8484 3136 8536 3188
rect 10324 3136 10376 3188
rect 12440 3068 12492 3120
rect 13820 3111 13872 3120
rect 13820 3077 13829 3111
rect 13829 3077 13863 3111
rect 13863 3077 13872 3111
rect 13820 3068 13872 3077
rect 2136 3000 2188 3052
rect 4804 3000 4856 3052
rect 1124 2932 1176 2984
rect 1860 2932 1912 2984
rect 7932 3000 7984 3052
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 6828 2932 6880 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 9864 2932 9916 2984
rect 10968 2975 11020 2984
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 12348 2932 12400 2984
rect 15384 3136 15436 3188
rect 18972 3136 19024 3188
rect 22284 3136 22336 3188
rect 14648 3068 14700 3120
rect 14924 3068 14976 3120
rect 20076 3068 20128 3120
rect 20352 3068 20404 3120
rect 14832 3000 14884 3052
rect 15108 3000 15160 3052
rect 20720 3000 20772 3052
rect 19340 2932 19392 2984
rect 21456 2932 21508 2984
rect 24676 2932 24728 2984
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 15384 2864 15436 2916
rect 19616 2864 19668 2916
rect 21180 2864 21232 2916
rect 22376 2864 22428 2916
rect 25412 2864 25464 2916
rect 1952 2796 2004 2848
rect 8024 2796 8076 2848
rect 13912 2796 13964 2848
rect 15292 2796 15344 2848
rect 15752 2796 15804 2848
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 22744 2796 22796 2848
rect 23388 2796 23440 2848
rect 25780 2796 25832 2848
rect 8912 2694 8964 2746
rect 8976 2694 9028 2746
rect 9040 2694 9092 2746
rect 9104 2694 9156 2746
rect 16843 2694 16895 2746
rect 16907 2694 16959 2746
rect 16971 2694 17023 2746
rect 17035 2694 17087 2746
rect 7748 2592 7800 2644
rect 1584 2524 1636 2576
rect 5356 2524 5408 2576
rect 5632 2524 5684 2576
rect 11152 2592 11204 2644
rect 15016 2592 15068 2644
rect 18604 2592 18656 2644
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 18696 2524 18748 2576
rect 22376 2567 22428 2576
rect 22376 2533 22385 2567
rect 22385 2533 22419 2567
rect 22419 2533 22428 2567
rect 22376 2524 22428 2533
rect 1952 2456 2004 2508
rect 4252 2499 4304 2508
rect 1860 2388 1912 2440
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 6460 2456 6512 2508
rect 7012 2456 7064 2508
rect 8024 2456 8076 2508
rect 9772 2456 9824 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 12440 2456 12492 2508
rect 13912 2456 13964 2508
rect 15384 2456 15436 2508
rect 19708 2456 19760 2508
rect 2320 2388 2372 2440
rect 6368 2388 6420 2440
rect 15108 2388 15160 2440
rect 17316 2388 17368 2440
rect 2044 2320 2096 2372
rect 14648 2320 14700 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 4436 2252 4488 2304
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 23388 2456 23440 2508
rect 22744 2431 22796 2440
rect 22744 2397 22753 2431
rect 22753 2397 22787 2431
rect 22787 2397 22796 2431
rect 22744 2388 22796 2397
rect 25044 2252 25096 2304
rect 4947 2150 4999 2202
rect 5011 2150 5063 2202
rect 5075 2150 5127 2202
rect 5139 2150 5191 2202
rect 12878 2150 12930 2202
rect 12942 2150 12994 2202
rect 13006 2150 13058 2202
rect 13070 2150 13122 2202
rect 20808 2150 20860 2202
rect 20872 2150 20924 2202
rect 20936 2150 20988 2202
rect 21000 2150 21052 2202
rect 2872 2048 2924 2100
rect 14280 2048 14332 2100
rect 2504 1980 2556 2032
rect 18604 1980 18656 2032
rect 4620 1912 4672 1964
rect 5080 1912 5132 1964
rect 12716 1300 12768 1352
rect 13268 1300 13320 1352
rect 11152 960 11204 1012
rect 12072 960 12124 1012
<< metal2 >>
rect 386 49200 442 50000
rect 1122 49200 1178 50000
rect 1950 49200 2006 50000
rect 2686 49200 2742 50000
rect 3514 49200 3570 50000
rect 4250 49200 4306 50000
rect 5078 49200 5134 50000
rect 5906 49200 5962 50000
rect 6642 49200 6698 50000
rect 7470 49200 7526 50000
rect 8206 49200 8262 50000
rect 9034 49200 9090 50000
rect 9770 49200 9826 50000
rect 10598 49200 10654 50000
rect 11426 49200 11482 50000
rect 12162 49200 12218 50000
rect 12990 49200 13046 50000
rect 13726 49200 13782 50000
rect 14554 49200 14610 50000
rect 15290 49200 15346 50000
rect 16118 49200 16174 50000
rect 16946 49200 17002 50000
rect 17682 49200 17738 50000
rect 18510 49200 18566 50000
rect 19246 49200 19302 50000
rect 20074 49200 20130 50000
rect 20810 49200 20866 50000
rect 21638 49200 21694 50000
rect 22466 49200 22522 50000
rect 23202 49200 23258 50000
rect 24030 49200 24086 50000
rect 24766 49200 24822 50000
rect 25594 49200 25650 50000
rect 400 45966 428 49200
rect 1136 46646 1164 49200
rect 1964 46714 1992 49200
rect 2700 46918 2728 49200
rect 3054 47288 3110 47297
rect 3054 47223 3110 47232
rect 3068 46986 3096 47223
rect 3056 46980 3108 46986
rect 3056 46922 3108 46928
rect 2688 46912 2740 46918
rect 2688 46854 2740 46860
rect 3332 46912 3384 46918
rect 3332 46854 3384 46860
rect 1952 46708 2004 46714
rect 1952 46650 2004 46656
rect 1124 46640 1176 46646
rect 1124 46582 1176 46588
rect 388 45960 440 45966
rect 388 45902 440 45908
rect 2688 45960 2740 45966
rect 2688 45902 2740 45908
rect 2596 43172 2648 43178
rect 2596 43114 2648 43120
rect 2608 41682 2636 43114
rect 1952 41676 2004 41682
rect 1952 41618 2004 41624
rect 2596 41676 2648 41682
rect 2596 41618 2648 41624
rect 1964 40390 1992 41618
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1964 38486 1992 40326
rect 2504 39976 2556 39982
rect 2504 39918 2556 39924
rect 2516 39098 2544 39918
rect 2700 39574 2728 45902
rect 3344 43194 3372 46854
rect 3424 44260 3476 44266
rect 3424 44202 3476 44208
rect 3436 43926 3464 44202
rect 3424 43920 3476 43926
rect 3424 43862 3476 43868
rect 3528 43314 3556 49200
rect 4160 44804 4212 44810
rect 4160 44746 4212 44752
rect 4172 44334 4200 44746
rect 4160 44328 4212 44334
rect 4160 44270 4212 44276
rect 3516 43308 3568 43314
rect 3516 43250 3568 43256
rect 3700 43240 3752 43246
rect 3344 43166 3556 43194
rect 3700 43182 3752 43188
rect 3148 43104 3200 43110
rect 3148 43046 3200 43052
rect 3160 41070 3188 43046
rect 3424 42152 3476 42158
rect 3424 42094 3476 42100
rect 3330 41712 3386 41721
rect 3330 41647 3386 41656
rect 2964 41064 3016 41070
rect 2964 41006 3016 41012
rect 3148 41064 3200 41070
rect 3148 41006 3200 41012
rect 2688 39568 2740 39574
rect 2688 39510 2740 39516
rect 2504 39092 2556 39098
rect 2504 39034 2556 39040
rect 2410 38992 2466 39001
rect 2410 38927 2412 38936
rect 2464 38927 2466 38936
rect 2412 38898 2464 38904
rect 1952 38480 2004 38486
rect 1952 38422 2004 38428
rect 2424 37330 2452 38898
rect 2412 37324 2464 37330
rect 2412 37266 2464 37272
rect 2700 35698 2728 39510
rect 2976 39001 3004 41006
rect 3148 40588 3200 40594
rect 3148 40530 3200 40536
rect 2962 38992 3018 39001
rect 2962 38927 3018 38936
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 3068 36786 3096 37062
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 3160 36582 3188 40530
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3344 36530 3372 41647
rect 3436 41274 3464 42094
rect 3424 41268 3476 41274
rect 3424 41210 3476 41216
rect 3528 40050 3556 43166
rect 3712 42362 3740 43182
rect 3976 42560 4028 42566
rect 3976 42502 4028 42508
rect 3700 42356 3752 42362
rect 3700 42298 3752 42304
rect 3988 42158 4016 42502
rect 4172 42294 4200 44270
rect 4160 42288 4212 42294
rect 4160 42230 4212 42236
rect 3976 42152 4028 42158
rect 3976 42094 4028 42100
rect 4172 41614 4200 42230
rect 4264 41818 4292 49200
rect 5092 46900 5120 49200
rect 5092 46872 5304 46900
rect 4921 46812 5217 46832
rect 4977 46810 5001 46812
rect 5057 46810 5081 46812
rect 5137 46810 5161 46812
rect 4999 46758 5001 46810
rect 5063 46758 5075 46810
rect 5137 46758 5139 46810
rect 4977 46756 5001 46758
rect 5057 46756 5081 46758
rect 5137 46756 5161 46758
rect 4921 46736 5217 46756
rect 4344 46708 4396 46714
rect 4344 46650 4396 46656
rect 4252 41812 4304 41818
rect 4252 41754 4304 41760
rect 4068 41608 4120 41614
rect 4068 41550 4120 41556
rect 4160 41608 4212 41614
rect 4212 41568 4292 41596
rect 4160 41550 4212 41556
rect 3700 41064 3752 41070
rect 3700 41006 3752 41012
rect 3516 40044 3568 40050
rect 3516 39986 3568 39992
rect 3528 39386 3556 39986
rect 3528 39358 3648 39386
rect 3424 38888 3476 38894
rect 3424 38830 3476 38836
rect 3436 38010 3464 38830
rect 3516 38820 3568 38826
rect 3516 38762 3568 38768
rect 3528 38554 3556 38762
rect 3516 38548 3568 38554
rect 3516 38490 3568 38496
rect 3620 38486 3648 39358
rect 3712 39098 3740 41006
rect 4080 41002 4108 41550
rect 4160 41472 4212 41478
rect 4160 41414 4212 41420
rect 4068 40996 4120 41002
rect 4068 40938 4120 40944
rect 4172 40730 4200 41414
rect 4160 40724 4212 40730
rect 4160 40666 4212 40672
rect 4264 39846 4292 41568
rect 4252 39840 4304 39846
rect 4252 39782 4304 39788
rect 3700 39092 3752 39098
rect 3700 39034 3752 39040
rect 3700 38888 3752 38894
rect 3700 38830 3752 38836
rect 3608 38480 3660 38486
rect 3608 38422 3660 38428
rect 3424 38004 3476 38010
rect 3424 37946 3476 37952
rect 3160 36310 3188 36518
rect 3344 36502 3464 36530
rect 3148 36304 3200 36310
rect 3148 36246 3200 36252
rect 3330 36136 3386 36145
rect 3330 36071 3386 36080
rect 3240 36032 3292 36038
rect 3240 35974 3292 35980
rect 2044 35692 2096 35698
rect 2044 35634 2096 35640
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 2056 35086 2084 35634
rect 2688 35556 2740 35562
rect 2688 35498 2740 35504
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1492 33516 1544 33522
rect 1492 33458 1544 33464
rect 1504 31346 1532 33458
rect 1964 32978 1992 33798
rect 1952 32972 2004 32978
rect 1952 32914 2004 32920
rect 1584 32224 1636 32230
rect 1584 32166 1636 32172
rect 1492 31340 1544 31346
rect 1492 31282 1544 31288
rect 1504 29714 1532 31282
rect 1492 29708 1544 29714
rect 1492 29650 1544 29656
rect 1504 29102 1532 29650
rect 1492 29096 1544 29102
rect 1492 29038 1544 29044
rect 1504 28558 1532 29038
rect 1492 28552 1544 28558
rect 1492 28494 1544 28500
rect 1504 28014 1532 28494
rect 1492 28008 1544 28014
rect 1492 27950 1544 27956
rect 1492 26580 1544 26586
rect 1492 26522 1544 26528
rect 1308 23860 1360 23866
rect 1308 23802 1360 23808
rect 388 8288 440 8294
rect 388 8230 440 8236
rect 112 4072 164 4078
rect 112 4014 164 4020
rect 124 800 152 4014
rect 400 800 428 8230
rect 756 4140 808 4146
rect 756 4082 808 4088
rect 768 800 796 4082
rect 1320 4078 1348 23802
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 18766 1440 20878
rect 1504 19922 1532 26522
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 18970 1532 19858
rect 1596 19417 1624 32166
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1676 28008 1728 28014
rect 1676 27950 1728 27956
rect 1688 25430 1716 27950
rect 1780 26586 1808 31078
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 1768 26580 1820 26586
rect 1768 26522 1820 26528
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1872 25906 1900 26182
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1964 25702 1992 26726
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1676 25424 1728 25430
rect 1676 25366 1728 25372
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1780 24410 1808 25298
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 1768 23656 1820 23662
rect 1768 23598 1820 23604
rect 1676 23588 1728 23594
rect 1676 23530 1728 23536
rect 1688 23186 1716 23530
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1676 22568 1728 22574
rect 1674 22536 1676 22545
rect 1728 22536 1730 22545
rect 1674 22471 1730 22480
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1688 20602 1716 20878
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1780 19310 1808 23598
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1872 22778 1900 22918
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 2056 20618 2084 35022
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2608 34066 2636 34478
rect 2596 34060 2648 34066
rect 2596 34002 2648 34008
rect 2700 33998 2728 35498
rect 3056 34604 3108 34610
rect 3056 34546 3108 34552
rect 2964 34400 3016 34406
rect 2964 34342 3016 34348
rect 2976 34066 3004 34342
rect 2964 34060 3016 34066
rect 2964 34002 3016 34008
rect 2688 33992 2740 33998
rect 2688 33934 2740 33940
rect 2700 33114 2728 33934
rect 3068 33114 3096 34546
rect 3148 34060 3200 34066
rect 3148 34002 3200 34008
rect 2688 33108 2740 33114
rect 2688 33050 2740 33056
rect 3056 33108 3108 33114
rect 3056 33050 3108 33056
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2504 30184 2556 30190
rect 2504 30126 2556 30132
rect 2516 29510 2544 30126
rect 2504 29504 2556 29510
rect 2504 29446 2556 29452
rect 2412 27872 2464 27878
rect 2412 27814 2464 27820
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2240 25294 2268 26318
rect 2424 25362 2452 27814
rect 2516 25650 2544 29446
rect 2792 29322 2820 31894
rect 2964 31884 3016 31890
rect 2884 31844 2964 31872
rect 2884 30326 2912 31844
rect 2964 31826 3016 31832
rect 3068 31278 3096 32302
rect 3160 31385 3188 34002
rect 3146 31376 3202 31385
rect 3146 31311 3202 31320
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3068 30938 3096 31214
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 2964 30796 3016 30802
rect 2964 30738 3016 30744
rect 2872 30320 2924 30326
rect 2872 30262 2924 30268
rect 2792 29294 2912 29322
rect 2780 28960 2832 28966
rect 2780 28902 2832 28908
rect 2688 28620 2740 28626
rect 2792 28608 2820 28902
rect 2740 28580 2820 28608
rect 2688 28562 2740 28568
rect 2792 28218 2820 28580
rect 2780 28212 2832 28218
rect 2780 28154 2832 28160
rect 2792 27878 2820 28154
rect 2884 28014 2912 29294
rect 2976 28626 3004 30738
rect 3068 30190 3096 30874
rect 3056 30184 3108 30190
rect 3056 30126 3108 30132
rect 3160 29866 3188 31311
rect 3068 29838 3188 29866
rect 3068 29034 3096 29838
rect 3148 29776 3200 29782
rect 3148 29718 3200 29724
rect 3056 29028 3108 29034
rect 3056 28970 3108 28976
rect 2964 28620 3016 28626
rect 2964 28562 3016 28568
rect 2872 28008 2924 28014
rect 2872 27950 2924 27956
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2780 27328 2832 27334
rect 2780 27270 2832 27276
rect 2594 26480 2650 26489
rect 2792 26450 2820 27270
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2594 26415 2596 26424
rect 2648 26415 2650 26424
rect 2780 26444 2832 26450
rect 2596 26386 2648 26392
rect 2780 26386 2832 26392
rect 2688 26376 2740 26382
rect 2688 26318 2740 26324
rect 2516 25622 2636 25650
rect 2412 25356 2464 25362
rect 2332 25316 2412 25344
rect 2228 25288 2280 25294
rect 2228 25230 2280 25236
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2148 23798 2176 24142
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 2240 23662 2268 25230
rect 2332 24750 2360 25316
rect 2412 25298 2464 25304
rect 2412 25220 2464 25226
rect 2412 25162 2464 25168
rect 2424 24750 2452 25162
rect 2320 24744 2372 24750
rect 2320 24686 2372 24692
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2240 21894 2268 23598
rect 2332 22710 2360 24686
rect 2424 24070 2452 24686
rect 2608 24274 2636 25622
rect 2700 24818 2728 26318
rect 2884 25838 2912 26930
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2884 25362 2912 25774
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2700 24342 2728 24754
rect 2688 24336 2740 24342
rect 2688 24278 2740 24284
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2516 24154 2544 24210
rect 2688 24200 2740 24206
rect 2516 24126 2636 24154
rect 2688 24142 2740 24148
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 1964 20590 2084 20618
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1412 18086 1440 18702
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 16658 1440 18022
rect 1688 17814 1716 18702
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 1676 17808 1728 17814
rect 1676 17750 1728 17756
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 15638 1716 16526
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1780 14890 1808 18090
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 13394 1716 14214
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12186 1440 13262
rect 1412 12158 1624 12186
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 9042 1440 12038
rect 1596 11150 1624 12158
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1688 11218 1716 11562
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1872 10674 1900 11086
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 9518 1900 10610
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 7954 1716 8298
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1872 7886 1900 9454
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1412 6254 1440 7822
rect 1964 7562 1992 20590
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 2240 20482 2268 21830
rect 2332 21010 2360 22034
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2056 19922 2084 20470
rect 2240 20454 2360 20482
rect 2332 20398 2360 20454
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2056 15978 2084 19858
rect 2148 19786 2176 19926
rect 2136 19780 2188 19786
rect 2136 19722 2188 19728
rect 2148 17134 2176 19722
rect 2240 17338 2268 20334
rect 2332 17746 2360 20334
rect 2424 19242 2452 24006
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2516 23118 2544 23802
rect 2608 23662 2636 24126
rect 2700 23866 2728 24142
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2504 23112 2556 23118
rect 2504 23054 2556 23060
rect 2516 20942 2544 23054
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2504 20324 2556 20330
rect 2504 20266 2556 20272
rect 2412 19236 2464 19242
rect 2412 19178 2464 19184
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2320 17740 2372 17746
rect 2424 17728 2452 18906
rect 2516 18290 2544 20266
rect 2608 19990 2636 23598
rect 2700 23322 2728 23666
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2700 22778 2728 23258
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2872 22432 2924 22438
rect 2792 22392 2872 22420
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 19514 2636 19654
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2504 17740 2556 17746
rect 2424 17700 2504 17728
rect 2320 17682 2372 17688
rect 2504 17682 2556 17688
rect 2608 17626 2636 19450
rect 2700 19446 2728 19790
rect 2792 19718 2820 22392
rect 2872 22374 2924 22380
rect 2976 22250 3004 28562
rect 3056 28552 3108 28558
rect 3056 28494 3108 28500
rect 3068 27130 3096 28494
rect 3160 28218 3188 29718
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 3148 27328 3200 27334
rect 3148 27270 3200 27276
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 3160 26994 3188 27270
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 3160 26450 3188 26726
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 3068 25430 3096 26318
rect 3160 25770 3188 26386
rect 3148 25764 3200 25770
rect 3148 25706 3200 25712
rect 3056 25424 3108 25430
rect 3056 25366 3108 25372
rect 3160 22642 3188 25706
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 2884 22222 3004 22250
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 2688 19440 2740 19446
rect 2688 19382 2740 19388
rect 2700 18222 2728 19382
rect 2884 19258 2912 22222
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 3056 21072 3108 21078
rect 3056 21014 3108 21020
rect 3068 20466 3096 21014
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3068 19854 3096 20402
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19310 3004 19654
rect 3068 19378 3096 19790
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 2792 19230 2912 19258
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2332 17598 2636 17626
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2332 16046 2360 17598
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2608 16182 2636 17206
rect 2700 17134 2728 17682
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 2056 12374 2084 15914
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2240 12442 2268 14486
rect 2332 12442 2360 15982
rect 2516 15570 2544 15982
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2412 15496 2464 15502
rect 2608 15450 2636 16118
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2412 15438 2464 15444
rect 2424 14414 2452 15438
rect 2516 15422 2636 15450
rect 2516 14958 2544 15422
rect 2700 15026 2728 15506
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2792 14958 2820 19230
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 15978 3004 17682
rect 3068 17202 3096 18158
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3068 16046 3096 16526
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15434 3004 15914
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 3160 15026 3188 21422
rect 3252 17354 3280 35974
rect 3344 26586 3372 36071
rect 3436 29782 3464 36502
rect 3712 34202 3740 38830
rect 4068 38412 4120 38418
rect 4068 38354 4120 38360
rect 3884 37800 3936 37806
rect 3884 37742 3936 37748
rect 3700 34196 3752 34202
rect 3700 34138 3752 34144
rect 3700 33312 3752 33318
rect 3700 33254 3752 33260
rect 3712 32978 3740 33254
rect 3700 32972 3752 32978
rect 3700 32914 3752 32920
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3514 30560 3570 30569
rect 3514 30495 3570 30504
rect 3528 30394 3556 30495
rect 3516 30388 3568 30394
rect 3516 30330 3568 30336
rect 3516 30184 3568 30190
rect 3516 30126 3568 30132
rect 3528 29850 3556 30126
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 3424 29776 3476 29782
rect 3424 29718 3476 29724
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3436 22488 3464 29582
rect 3528 26246 3556 29786
rect 3620 29646 3648 30874
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3608 29028 3660 29034
rect 3608 28970 3660 28976
rect 3516 26240 3568 26246
rect 3516 26182 3568 26188
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3528 23526 3556 24686
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3344 22460 3464 22488
rect 3344 21486 3372 22460
rect 3424 21956 3476 21962
rect 3424 21898 3476 21904
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3344 17542 3372 21422
rect 3436 19417 3464 21898
rect 3620 20058 3648 28970
rect 3712 21078 3740 32914
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 3804 28694 3832 32302
rect 3792 28688 3844 28694
rect 3792 28630 3844 28636
rect 3792 27532 3844 27538
rect 3792 27474 3844 27480
rect 3804 26994 3832 27474
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3792 26512 3844 26518
rect 3790 26480 3792 26489
rect 3844 26480 3846 26489
rect 3790 26415 3846 26424
rect 3896 25906 3924 37742
rect 4080 36718 4108 38354
rect 4160 37324 4212 37330
rect 4160 37266 4212 37272
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 4172 34950 4200 37266
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 4264 36786 4292 37198
rect 4356 36922 4384 46650
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 4816 45506 4844 45902
rect 4921 45724 5217 45744
rect 4977 45722 5001 45724
rect 5057 45722 5081 45724
rect 5137 45722 5161 45724
rect 4999 45670 5001 45722
rect 5063 45670 5075 45722
rect 5137 45670 5139 45722
rect 4977 45668 5001 45670
rect 5057 45668 5081 45670
rect 5137 45668 5161 45670
rect 4921 45648 5217 45668
rect 5276 45506 5304 46872
rect 5724 46640 5776 46646
rect 5724 46582 5776 46588
rect 5448 46436 5500 46442
rect 5448 46378 5500 46384
rect 5356 45960 5408 45966
rect 5356 45902 5408 45908
rect 5368 45626 5396 45902
rect 5356 45620 5408 45626
rect 5356 45562 5408 45568
rect 4816 45478 4936 45506
rect 5276 45478 5396 45506
rect 4712 45416 4764 45422
rect 4712 45358 4764 45364
rect 4724 44946 4752 45358
rect 4804 45280 4856 45286
rect 4804 45222 4856 45228
rect 4816 45014 4844 45222
rect 4804 45008 4856 45014
rect 4804 44950 4856 44956
rect 4712 44940 4764 44946
rect 4632 44900 4712 44928
rect 4632 43722 4660 44900
rect 4712 44882 4764 44888
rect 4908 44810 4936 45478
rect 5264 45416 5316 45422
rect 5264 45358 5316 45364
rect 4896 44804 4948 44810
rect 4896 44746 4948 44752
rect 4921 44636 5217 44656
rect 4977 44634 5001 44636
rect 5057 44634 5081 44636
rect 5137 44634 5161 44636
rect 4999 44582 5001 44634
rect 5063 44582 5075 44634
rect 5137 44582 5139 44634
rect 4977 44580 5001 44582
rect 5057 44580 5081 44582
rect 5137 44580 5161 44582
rect 4921 44560 5217 44580
rect 4804 44328 4856 44334
rect 4804 44270 4856 44276
rect 4712 43852 4764 43858
rect 4712 43794 4764 43800
rect 4620 43716 4672 43722
rect 4620 43658 4672 43664
rect 4436 42832 4488 42838
rect 4436 42774 4488 42780
rect 4448 41478 4476 42774
rect 4632 42634 4660 43658
rect 4620 42628 4672 42634
rect 4620 42570 4672 42576
rect 4632 42362 4660 42570
rect 4620 42356 4672 42362
rect 4620 42298 4672 42304
rect 4528 41608 4580 41614
rect 4528 41550 4580 41556
rect 4436 41472 4488 41478
rect 4436 41414 4488 41420
rect 4540 41138 4568 41550
rect 4632 41274 4660 42298
rect 4620 41268 4672 41274
rect 4620 41210 4672 41216
rect 4528 41132 4580 41138
rect 4528 41074 4580 41080
rect 4436 40588 4488 40594
rect 4436 40530 4488 40536
rect 4344 36916 4396 36922
rect 4344 36858 4396 36864
rect 4252 36780 4304 36786
rect 4252 36722 4304 36728
rect 4448 35714 4476 40530
rect 4724 39506 4752 43794
rect 4816 43654 4844 44270
rect 4804 43648 4856 43654
rect 4804 43590 4856 43596
rect 4921 43548 5217 43568
rect 4977 43546 5001 43548
rect 5057 43546 5081 43548
rect 5137 43546 5161 43548
rect 4999 43494 5001 43546
rect 5063 43494 5075 43546
rect 5137 43494 5139 43546
rect 4977 43492 5001 43494
rect 5057 43492 5081 43494
rect 5137 43492 5161 43494
rect 4921 43472 5217 43492
rect 4804 42628 4856 42634
rect 4804 42570 4856 42576
rect 4816 42294 4844 42570
rect 4921 42460 5217 42480
rect 4977 42458 5001 42460
rect 5057 42458 5081 42460
rect 5137 42458 5161 42460
rect 4999 42406 5001 42458
rect 5063 42406 5075 42458
rect 5137 42406 5139 42458
rect 4977 42404 5001 42406
rect 5057 42404 5081 42406
rect 5137 42404 5161 42406
rect 4921 42384 5217 42404
rect 4804 42288 4856 42294
rect 4804 42230 4856 42236
rect 4921 41372 5217 41392
rect 4977 41370 5001 41372
rect 5057 41370 5081 41372
rect 5137 41370 5161 41372
rect 4999 41318 5001 41370
rect 5063 41318 5075 41370
rect 5137 41318 5139 41370
rect 4977 41316 5001 41318
rect 5057 41316 5081 41318
rect 5137 41316 5161 41318
rect 4921 41296 5217 41316
rect 4804 41064 4856 41070
rect 4804 41006 4856 41012
rect 4816 40594 4844 41006
rect 4804 40588 4856 40594
rect 4804 40530 4856 40536
rect 4921 40284 5217 40304
rect 4977 40282 5001 40284
rect 5057 40282 5081 40284
rect 5137 40282 5161 40284
rect 4999 40230 5001 40282
rect 5063 40230 5075 40282
rect 5137 40230 5139 40282
rect 4977 40228 5001 40230
rect 5057 40228 5081 40230
rect 5137 40228 5161 40230
rect 4921 40208 5217 40228
rect 5276 40186 5304 45358
rect 5368 44538 5396 45478
rect 5460 45422 5488 46378
rect 5632 46368 5684 46374
rect 5632 46310 5684 46316
rect 5448 45416 5500 45422
rect 5448 45358 5500 45364
rect 5460 44962 5488 45358
rect 5644 45354 5672 46310
rect 5632 45348 5684 45354
rect 5632 45290 5684 45296
rect 5460 44934 5580 44962
rect 5448 44872 5500 44878
rect 5448 44814 5500 44820
rect 5356 44532 5408 44538
rect 5356 44474 5408 44480
rect 5356 44328 5408 44334
rect 5356 44270 5408 44276
rect 5368 44198 5396 44270
rect 5356 44192 5408 44198
rect 5356 44134 5408 44140
rect 5368 43246 5396 44134
rect 5356 43240 5408 43246
rect 5356 43182 5408 43188
rect 5368 42838 5396 43182
rect 5356 42832 5408 42838
rect 5356 42774 5408 42780
rect 5356 42696 5408 42702
rect 5356 42638 5408 42644
rect 5368 42158 5396 42638
rect 5356 42152 5408 42158
rect 5356 42094 5408 42100
rect 5356 40588 5408 40594
rect 5356 40530 5408 40536
rect 5264 40180 5316 40186
rect 5264 40122 5316 40128
rect 5368 39982 5396 40530
rect 4804 39976 4856 39982
rect 4804 39918 4856 39924
rect 5356 39976 5408 39982
rect 5356 39918 5408 39924
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 4712 39500 4764 39506
rect 4712 39442 4764 39448
rect 4528 39296 4580 39302
rect 4528 39238 4580 39244
rect 4540 38962 4568 39238
rect 4528 38956 4580 38962
rect 4528 38898 4580 38904
rect 4540 37806 4568 38898
rect 4528 37800 4580 37806
rect 4528 37742 4580 37748
rect 4356 35686 4476 35714
rect 4252 35148 4304 35154
rect 4252 35090 4304 35096
rect 4160 34944 4212 34950
rect 4160 34886 4212 34892
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 3988 32502 4016 33390
rect 4080 33114 4108 34478
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3976 32496 4028 32502
rect 3976 32438 4028 32444
rect 4080 32366 4108 33050
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 3976 30660 4028 30666
rect 3976 30602 4028 30608
rect 3988 28422 4016 30602
rect 4172 30190 4200 33390
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4080 29102 4108 30126
rect 4160 30048 4212 30054
rect 4160 29990 4212 29996
rect 4172 29714 4200 29990
rect 4160 29708 4212 29714
rect 4160 29650 4212 29656
rect 4160 29164 4212 29170
rect 4160 29106 4212 29112
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4080 28762 4108 29038
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 4080 27606 4108 28698
rect 4172 28665 4200 29106
rect 4158 28656 4214 28665
rect 4158 28591 4214 28600
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 3988 27062 4016 27406
rect 4172 27130 4200 27406
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4080 26858 4108 26930
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 3976 26580 4028 26586
rect 3976 26522 4028 26528
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3422 19408 3478 19417
rect 3620 19378 3648 19994
rect 3422 19343 3478 19352
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3252 17326 3372 17354
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2516 14482 2544 14894
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11762 2084 12310
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2332 11694 2360 12378
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2042 10024 2098 10033
rect 2042 9959 2044 9968
rect 2096 9959 2098 9968
rect 2044 9930 2096 9936
rect 2148 9178 2176 11630
rect 2424 11626 2452 14350
rect 2516 13530 2544 14418
rect 2608 14414 2636 14826
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 10266 2452 11562
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 1964 7534 2084 7562
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6322 1716 6734
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1768 6248 1820 6254
rect 1820 6196 1900 6202
rect 1768 6190 1900 6196
rect 1780 6174 1900 6190
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1504 4146 1532 5714
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1124 2984 1176 2990
rect 1124 2926 1176 2932
rect 1136 800 1164 2926
rect 1412 1306 1440 3334
rect 1596 2582 1624 5510
rect 1872 4078 1900 6174
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1872 2990 1900 4014
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 1964 2514 1992 2790
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1412 1278 1532 1306
rect 1504 800 1532 1278
rect 1872 800 1900 2382
rect 2056 2378 2084 7534
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2148 4146 2176 4558
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2148 3058 2176 3470
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 2240 800 2268 4082
rect 2332 2446 2360 8502
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 6186 2452 7142
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2516 4026 2544 12650
rect 2608 12102 2636 14350
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10130 2636 10406
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2700 8566 2728 14214
rect 2792 13870 2820 14894
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 13938 3004 14350
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12322 2820 12650
rect 2792 12294 2912 12322
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2792 11354 2820 12174
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2884 8974 2912 12294
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 7206 2728 8366
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 6730 2728 7142
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2424 3998 2544 4026
rect 2424 2825 2452 3998
rect 2410 2816 2466 2825
rect 2410 2751 2466 2760
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2038 2544 2246
rect 2504 2032 2556 2038
rect 2504 1974 2556 1980
rect 2608 800 2636 5034
rect 2700 4622 2728 6666
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 3602 2728 4558
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2884 2106 2912 8910
rect 2976 8838 3004 10066
rect 3068 9654 3096 12718
rect 3160 12458 3188 14962
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 13938 3280 14758
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3344 12850 3372 17326
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3160 12430 3280 12458
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10130 3188 10542
rect 3252 10538 3280 12430
rect 3436 12374 3464 19178
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 18290 3556 18566
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3608 18080 3660 18086
rect 3660 18028 3740 18034
rect 3608 18022 3740 18028
rect 3620 18006 3740 18022
rect 3712 17542 3740 18006
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3160 9110 3188 10066
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 7750 3004 8366
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 6866 3004 7686
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6390 3004 6666
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3068 5914 3096 6598
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2976 5001 3004 5170
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 2976 4690 3004 4927
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2976 800 3004 3130
rect 3252 800 3280 10474
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 3210 3464 9318
rect 3528 6662 3556 17478
rect 3712 16046 3740 17478
rect 3804 16726 3832 23462
rect 3884 23180 3936 23186
rect 3884 23122 3936 23128
rect 3896 21486 3924 23122
rect 3988 21690 4016 26522
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 4080 26314 4108 26386
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4066 24984 4122 24993
rect 4066 24919 4122 24928
rect 4080 24886 4108 24919
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 4080 23322 4108 24686
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4172 23202 4200 26930
rect 4264 23730 4292 35090
rect 4356 34746 4384 35686
rect 4436 35624 4488 35630
rect 4436 35566 4488 35572
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 4448 31482 4476 35566
rect 4528 34536 4580 34542
rect 4528 34478 4580 34484
rect 4540 32910 4568 34478
rect 4632 33522 4660 39442
rect 4712 35624 4764 35630
rect 4712 35566 4764 35572
rect 4724 35494 4752 35566
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4724 34542 4752 35430
rect 4712 34536 4764 34542
rect 4712 34478 4764 34484
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 4816 33266 4844 39918
rect 5264 39840 5316 39846
rect 5264 39782 5316 39788
rect 4921 39196 5217 39216
rect 4977 39194 5001 39196
rect 5057 39194 5081 39196
rect 5137 39194 5161 39196
rect 4999 39142 5001 39194
rect 5063 39142 5075 39194
rect 5137 39142 5139 39194
rect 4977 39140 5001 39142
rect 5057 39140 5081 39142
rect 5137 39140 5161 39142
rect 4921 39120 5217 39140
rect 5276 38162 5304 39782
rect 5368 39506 5396 39918
rect 5356 39500 5408 39506
rect 5356 39442 5408 39448
rect 5368 38962 5396 39442
rect 5356 38956 5408 38962
rect 5356 38898 5408 38904
rect 5460 38282 5488 44814
rect 5552 44334 5580 44934
rect 5540 44328 5592 44334
rect 5540 44270 5592 44276
rect 5540 42152 5592 42158
rect 5540 42094 5592 42100
rect 5552 38962 5580 42094
rect 5540 38956 5592 38962
rect 5540 38898 5592 38904
rect 5540 38752 5592 38758
rect 5540 38694 5592 38700
rect 5448 38276 5500 38282
rect 5448 38218 5500 38224
rect 5276 38134 5488 38162
rect 4921 38108 5217 38128
rect 4977 38106 5001 38108
rect 5057 38106 5081 38108
rect 5137 38106 5161 38108
rect 4999 38054 5001 38106
rect 5063 38054 5075 38106
rect 5137 38054 5139 38106
rect 4977 38052 5001 38054
rect 5057 38052 5081 38054
rect 5137 38052 5161 38054
rect 4921 38032 5217 38052
rect 5460 37262 5488 38134
rect 5552 37806 5580 38694
rect 5540 37800 5592 37806
rect 5540 37742 5592 37748
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 4921 37020 5217 37040
rect 4977 37018 5001 37020
rect 5057 37018 5081 37020
rect 5137 37018 5161 37020
rect 4999 36966 5001 37018
rect 5063 36966 5075 37018
rect 5137 36966 5139 37018
rect 4977 36964 5001 36966
rect 5057 36964 5081 36966
rect 5137 36964 5161 36966
rect 4921 36944 5217 36964
rect 5356 36712 5408 36718
rect 5356 36654 5408 36660
rect 5368 36242 5396 36654
rect 5460 36258 5488 37198
rect 5552 36582 5580 37742
rect 5736 37466 5764 46582
rect 5920 46510 5948 49200
rect 6276 46980 6328 46986
rect 6276 46922 6328 46928
rect 5908 46504 5960 46510
rect 5908 46446 5960 46452
rect 5920 46170 5948 46446
rect 5908 46164 5960 46170
rect 5908 46106 5960 46112
rect 5908 43172 5960 43178
rect 5908 43114 5960 43120
rect 5816 42696 5868 42702
rect 5816 42638 5868 42644
rect 5828 42362 5856 42638
rect 5816 42356 5868 42362
rect 5816 42298 5868 42304
rect 5920 40662 5948 43114
rect 5908 40656 5960 40662
rect 5908 40598 5960 40604
rect 5908 38888 5960 38894
rect 5908 38830 5960 38836
rect 5816 38820 5868 38826
rect 5816 38762 5868 38768
rect 5632 37460 5684 37466
rect 5632 37402 5684 37408
rect 5724 37460 5776 37466
rect 5724 37402 5776 37408
rect 5644 36922 5672 37402
rect 5632 36916 5684 36922
rect 5632 36858 5684 36864
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 5552 36394 5580 36518
rect 5552 36366 5672 36394
rect 5172 36236 5224 36242
rect 5172 36178 5224 36184
rect 5356 36236 5408 36242
rect 5460 36230 5580 36258
rect 5356 36178 5408 36184
rect 5184 36020 5212 36178
rect 5552 36174 5580 36230
rect 5540 36168 5592 36174
rect 5540 36110 5592 36116
rect 5184 35992 5488 36020
rect 4921 35932 5217 35952
rect 4977 35930 5001 35932
rect 5057 35930 5081 35932
rect 5137 35930 5161 35932
rect 4999 35878 5001 35930
rect 5063 35878 5075 35930
rect 5137 35878 5139 35930
rect 4977 35876 5001 35878
rect 5057 35876 5081 35878
rect 5137 35876 5161 35878
rect 4921 35856 5217 35876
rect 5356 35284 5408 35290
rect 5356 35226 5408 35232
rect 4921 34844 5217 34864
rect 4977 34842 5001 34844
rect 5057 34842 5081 34844
rect 5137 34842 5161 34844
rect 4999 34790 5001 34842
rect 5063 34790 5075 34842
rect 5137 34790 5139 34842
rect 4977 34788 5001 34790
rect 5057 34788 5081 34790
rect 5137 34788 5161 34790
rect 4921 34768 5217 34788
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 4921 33756 5217 33776
rect 4977 33754 5001 33756
rect 5057 33754 5081 33756
rect 5137 33754 5161 33756
rect 4999 33702 5001 33754
rect 5063 33702 5075 33754
rect 5137 33702 5139 33754
rect 4977 33700 5001 33702
rect 5057 33700 5081 33702
rect 5137 33700 5161 33702
rect 4921 33680 5217 33700
rect 4632 33238 4844 33266
rect 4528 32904 4580 32910
rect 4528 32846 4580 32852
rect 4528 31748 4580 31754
rect 4528 31690 4580 31696
rect 4436 31476 4488 31482
rect 4436 31418 4488 31424
rect 4436 30728 4488 30734
rect 4436 30670 4488 30676
rect 4344 30116 4396 30122
rect 4344 30058 4396 30064
rect 4356 28694 4384 30058
rect 4448 29850 4476 30670
rect 4436 29844 4488 29850
rect 4436 29786 4488 29792
rect 4540 29186 4568 31690
rect 4448 29158 4568 29186
rect 4344 28688 4396 28694
rect 4344 28630 4396 28636
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4356 25906 4384 28358
rect 4448 26790 4476 29158
rect 4528 29096 4580 29102
rect 4528 29038 4580 29044
rect 4540 28490 4568 29038
rect 4528 28484 4580 28490
rect 4528 28426 4580 28432
rect 4526 28384 4582 28393
rect 4526 28319 4582 28328
rect 4540 26994 4568 28319
rect 4632 28082 4660 33238
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 4724 32230 4752 32846
rect 4921 32668 5217 32688
rect 4977 32666 5001 32668
rect 5057 32666 5081 32668
rect 5137 32666 5161 32668
rect 4999 32614 5001 32666
rect 5063 32614 5075 32666
rect 5137 32614 5139 32666
rect 4977 32612 5001 32614
rect 5057 32612 5081 32614
rect 5137 32612 5161 32614
rect 4921 32592 5217 32612
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4620 28076 4672 28082
rect 4620 28018 4672 28024
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4724 26874 4752 32166
rect 4816 31890 4844 32302
rect 5276 32230 5304 34478
rect 5368 34241 5396 35226
rect 5354 34232 5410 34241
rect 5354 34167 5410 34176
rect 5356 33312 5408 33318
rect 5356 33254 5408 33260
rect 5264 32224 5316 32230
rect 5264 32166 5316 32172
rect 4804 31884 4856 31890
rect 4804 31826 4856 31832
rect 4816 30938 4844 31826
rect 4921 31580 5217 31600
rect 4977 31578 5001 31580
rect 5057 31578 5081 31580
rect 5137 31578 5161 31580
rect 4999 31526 5001 31578
rect 5063 31526 5075 31578
rect 5137 31526 5139 31578
rect 4977 31524 5001 31526
rect 5057 31524 5081 31526
rect 5137 31524 5161 31526
rect 4921 31504 5217 31524
rect 5172 31408 5224 31414
rect 4894 31376 4950 31385
rect 5172 31350 5224 31356
rect 4894 31311 4950 31320
rect 4908 31278 4936 31311
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4804 30932 4856 30938
rect 4804 30874 4856 30880
rect 5184 30580 5212 31350
rect 5276 30802 5304 32166
rect 5368 31686 5396 33254
rect 5460 31754 5488 35992
rect 5644 35630 5672 36366
rect 5736 36242 5764 37402
rect 5724 36236 5776 36242
rect 5724 36178 5776 36184
rect 5632 35624 5684 35630
rect 5632 35566 5684 35572
rect 5724 35148 5776 35154
rect 5724 35090 5776 35096
rect 5632 34672 5684 34678
rect 5632 34614 5684 34620
rect 5540 34400 5592 34406
rect 5540 34342 5592 34348
rect 5552 33454 5580 34342
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5644 33386 5672 34614
rect 5736 33998 5764 35090
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 5736 33590 5764 33934
rect 5724 33584 5776 33590
rect 5724 33526 5776 33532
rect 5828 33538 5856 38762
rect 5920 38350 5948 38830
rect 6000 38412 6052 38418
rect 6000 38354 6052 38360
rect 5908 38344 5960 38350
rect 5908 38286 5960 38292
rect 5908 34060 5960 34066
rect 5908 34002 5960 34008
rect 5920 33658 5948 34002
rect 6012 33946 6040 38354
rect 6288 37942 6316 46922
rect 6368 43852 6420 43858
rect 6368 43794 6420 43800
rect 6380 40050 6408 43794
rect 6656 42702 6684 49200
rect 7484 45422 7512 49200
rect 8220 47274 8248 49200
rect 9048 47546 9076 49200
rect 9048 47518 9352 47546
rect 8886 47356 9182 47376
rect 8942 47354 8966 47356
rect 9022 47354 9046 47356
rect 9102 47354 9126 47356
rect 8964 47302 8966 47354
rect 9028 47302 9040 47354
rect 9102 47302 9104 47354
rect 8942 47300 8966 47302
rect 9022 47300 9046 47302
rect 9102 47300 9126 47302
rect 8886 47280 9182 47300
rect 8128 47246 8248 47274
rect 7656 46504 7708 46510
rect 7656 46446 7708 46452
rect 7472 45416 7524 45422
rect 7472 45358 7524 45364
rect 7484 45082 7512 45358
rect 7472 45076 7524 45082
rect 7472 45018 7524 45024
rect 7668 44402 7696 46446
rect 7748 45416 7800 45422
rect 7748 45358 7800 45364
rect 7656 44396 7708 44402
rect 7656 44338 7708 44344
rect 7668 44010 7696 44338
rect 7484 43982 7696 44010
rect 7380 43920 7432 43926
rect 7380 43862 7432 43868
rect 6920 43648 6972 43654
rect 6920 43590 6972 43596
rect 6644 42696 6696 42702
rect 6644 42638 6696 42644
rect 6828 42560 6880 42566
rect 6828 42502 6880 42508
rect 6840 41138 6868 42502
rect 6932 42226 6960 43590
rect 7392 43246 7420 43862
rect 7380 43240 7432 43246
rect 7380 43182 7432 43188
rect 6920 42220 6972 42226
rect 6920 42162 6972 42168
rect 7012 42220 7064 42226
rect 7012 42162 7064 42168
rect 6932 41614 6960 42162
rect 6920 41608 6972 41614
rect 6920 41550 6972 41556
rect 6828 41132 6880 41138
rect 6828 41074 6880 41080
rect 6736 40588 6788 40594
rect 6736 40530 6788 40536
rect 6368 40044 6420 40050
rect 6368 39986 6420 39992
rect 6380 39370 6408 39986
rect 6552 39432 6604 39438
rect 6552 39374 6604 39380
rect 6368 39364 6420 39370
rect 6368 39306 6420 39312
rect 6380 38010 6408 39306
rect 6368 38004 6420 38010
rect 6368 37946 6420 37952
rect 6276 37936 6328 37942
rect 6276 37878 6328 37884
rect 6368 37800 6420 37806
rect 6368 37742 6420 37748
rect 6092 35556 6144 35562
rect 6092 35498 6144 35504
rect 6104 34066 6132 35498
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6012 33918 6132 33946
rect 5908 33652 5960 33658
rect 5908 33594 5960 33600
rect 5632 33380 5684 33386
rect 5632 33322 5684 33328
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5448 31748 5500 31754
rect 5448 31690 5500 31696
rect 5356 31680 5408 31686
rect 5552 31668 5580 33254
rect 5644 32212 5672 33322
rect 5736 32858 5764 33526
rect 5828 33510 6040 33538
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 5920 32978 5948 33254
rect 5908 32972 5960 32978
rect 5908 32914 5960 32920
rect 5736 32830 5856 32858
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5736 32366 5764 32710
rect 5828 32502 5856 32830
rect 5816 32496 5868 32502
rect 5816 32438 5868 32444
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 5644 32184 5948 32212
rect 5724 32020 5776 32026
rect 5724 31962 5776 31968
rect 5356 31622 5408 31628
rect 5446 31648 5502 31657
rect 5368 30802 5396 31622
rect 5552 31640 5672 31668
rect 5446 31583 5502 31592
rect 5264 30796 5316 30802
rect 5264 30738 5316 30744
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 5356 30660 5408 30666
rect 5356 30602 5408 30608
rect 5184 30552 5304 30580
rect 4921 30492 5217 30512
rect 4977 30490 5001 30492
rect 5057 30490 5081 30492
rect 5137 30490 5161 30492
rect 4999 30438 5001 30490
rect 5063 30438 5075 30490
rect 5137 30438 5139 30490
rect 4977 30436 5001 30438
rect 5057 30436 5081 30438
rect 5137 30436 5161 30438
rect 4921 30416 5217 30436
rect 4921 29404 5217 29424
rect 4977 29402 5001 29404
rect 5057 29402 5081 29404
rect 5137 29402 5161 29404
rect 4999 29350 5001 29402
rect 5063 29350 5075 29402
rect 5137 29350 5139 29402
rect 4977 29348 5001 29350
rect 5057 29348 5081 29350
rect 5137 29348 5161 29350
rect 4921 29328 5217 29348
rect 5276 29288 5304 30552
rect 5368 29850 5396 30602
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5092 29260 5304 29288
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4816 28665 4844 28970
rect 4802 28656 4858 28665
rect 4802 28591 4858 28600
rect 4804 28552 4856 28558
rect 4802 28520 4804 28529
rect 5092 28529 5120 29260
rect 4856 28520 4858 28529
rect 4802 28455 4858 28464
rect 5078 28520 5134 28529
rect 5078 28455 5134 28464
rect 5264 28484 5316 28490
rect 5264 28426 5316 28432
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4540 26846 4752 26874
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 4436 26240 4488 26246
rect 4436 26182 4488 26188
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 4356 24750 4384 25842
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 4080 23174 4200 23202
rect 4080 22710 4108 23174
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 4080 21486 4108 21966
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 4080 21146 4108 21422
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4172 18766 4200 23054
rect 4356 22930 4384 23666
rect 4264 22902 4384 22930
rect 4264 21593 4292 22902
rect 4448 22794 4476 26182
rect 4356 22766 4476 22794
rect 4250 21584 4306 21593
rect 4250 21519 4306 21528
rect 4356 21434 4384 22766
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4264 21406 4384 21434
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 3620 15094 3648 15506
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 3712 14414 3740 15982
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3620 3398 3648 11562
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3712 10062 3740 10746
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 7342 3740 9998
rect 3804 7546 3832 16662
rect 3896 9382 3924 18702
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4172 17218 4200 18226
rect 4080 17190 4200 17218
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16114 4016 16390
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4080 15570 4108 17190
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16590 4200 17070
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 16114 4200 16526
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14074 4016 14894
rect 4080 14890 4108 15506
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 14550 4108 14826
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3712 5302 3740 6870
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3712 4214 3740 5238
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4622 3832 5102
rect 3896 5030 3924 9046
rect 3988 8090 4016 13806
rect 4080 12306 4108 13874
rect 4172 12714 4200 15438
rect 4264 14464 4292 21406
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4356 21010 4384 21286
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4342 20904 4398 20913
rect 4342 20839 4398 20848
rect 4356 19310 4384 20839
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4356 18290 4384 19110
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4356 17746 4384 18022
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4356 17338 4384 17682
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4356 14958 4384 16458
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4264 14436 4384 14464
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4080 8906 4108 11766
rect 4264 11218 4292 12786
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10674 4200 11086
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4080 7818 4108 8191
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3804 4146 3832 4558
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3436 3182 3648 3210
rect 3620 800 3648 3182
rect 3988 800 4016 7482
rect 4172 6934 4200 8978
rect 4356 8786 4384 14436
rect 4448 9081 4476 22646
rect 4540 19394 4568 26846
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4632 21962 4660 26726
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4724 24954 4752 25230
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4724 22710 4752 23598
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21350 4752 21830
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4816 20398 4844 28358
rect 4921 28316 5217 28336
rect 4977 28314 5001 28316
rect 5057 28314 5081 28316
rect 5137 28314 5161 28316
rect 4999 28262 5001 28314
rect 5063 28262 5075 28314
rect 5137 28262 5139 28314
rect 4977 28260 5001 28262
rect 5057 28260 5081 28262
rect 5137 28260 5161 28262
rect 4921 28240 5217 28260
rect 4894 28112 4950 28121
rect 5276 28082 5304 28426
rect 4894 28047 4950 28056
rect 5264 28076 5316 28082
rect 4908 27674 4936 28047
rect 5264 28018 5316 28024
rect 5368 28014 5396 29786
rect 5356 28008 5408 28014
rect 5356 27950 5408 27956
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 4908 27538 4936 27610
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 4921 27228 5217 27248
rect 4977 27226 5001 27228
rect 5057 27226 5081 27228
rect 5137 27226 5161 27228
rect 4999 27174 5001 27226
rect 5063 27174 5075 27226
rect 5137 27174 5139 27226
rect 4977 27172 5001 27174
rect 5057 27172 5081 27174
rect 5137 27172 5161 27174
rect 4921 27152 5217 27172
rect 5276 26314 5304 27474
rect 5264 26308 5316 26314
rect 5264 26250 5316 26256
rect 4921 26140 5217 26160
rect 4977 26138 5001 26140
rect 5057 26138 5081 26140
rect 5137 26138 5161 26140
rect 4999 26086 5001 26138
rect 5063 26086 5075 26138
rect 5137 26086 5139 26138
rect 4977 26084 5001 26086
rect 5057 26084 5081 26086
rect 5137 26084 5161 26086
rect 4921 26064 5217 26084
rect 5368 25906 5396 27950
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5264 25832 5316 25838
rect 5264 25774 5316 25780
rect 4921 25052 5217 25072
rect 4977 25050 5001 25052
rect 5057 25050 5081 25052
rect 5137 25050 5161 25052
rect 4999 24998 5001 25050
rect 5063 24998 5075 25050
rect 5137 24998 5139 25050
rect 4977 24996 5001 24998
rect 5057 24996 5081 24998
rect 5137 24996 5161 24998
rect 4921 24976 5217 24996
rect 4921 23964 5217 23984
rect 4977 23962 5001 23964
rect 5057 23962 5081 23964
rect 5137 23962 5161 23964
rect 4999 23910 5001 23962
rect 5063 23910 5075 23962
rect 5137 23910 5139 23962
rect 4977 23908 5001 23910
rect 5057 23908 5081 23910
rect 5137 23908 5161 23910
rect 4921 23888 5217 23908
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 5000 23186 5028 23530
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 4921 22876 5217 22896
rect 4977 22874 5001 22876
rect 5057 22874 5081 22876
rect 5137 22874 5161 22876
rect 4999 22822 5001 22874
rect 5063 22822 5075 22874
rect 5137 22822 5139 22874
rect 4977 22820 5001 22822
rect 5057 22820 5081 22822
rect 5137 22820 5161 22822
rect 4921 22800 5217 22820
rect 5276 22760 5304 25774
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5368 23254 5396 24142
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5354 23080 5410 23089
rect 5354 23015 5410 23024
rect 5092 22732 5304 22760
rect 4988 22704 5040 22710
rect 4988 22646 5040 22652
rect 5000 22098 5028 22646
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 5092 22030 5120 22732
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 4921 21788 5217 21808
rect 4977 21786 5001 21788
rect 5057 21786 5081 21788
rect 5137 21786 5161 21788
rect 4999 21734 5001 21786
rect 5063 21734 5075 21786
rect 5137 21734 5139 21786
rect 4977 21732 5001 21734
rect 5057 21732 5081 21734
rect 5137 21732 5161 21734
rect 4921 21712 5217 21732
rect 4921 20700 5217 20720
rect 4977 20698 5001 20700
rect 5057 20698 5081 20700
rect 5137 20698 5161 20700
rect 4999 20646 5001 20698
rect 5063 20646 5075 20698
rect 5137 20646 5139 20698
rect 4977 20644 5001 20646
rect 5057 20644 5081 20646
rect 5137 20644 5161 20646
rect 4921 20624 5217 20644
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4724 19514 4752 20334
rect 4921 19612 5217 19632
rect 4977 19610 5001 19612
rect 5057 19610 5081 19612
rect 5137 19610 5161 19612
rect 4999 19558 5001 19610
rect 5063 19558 5075 19610
rect 5137 19558 5139 19610
rect 4977 19556 5001 19558
rect 5057 19556 5081 19558
rect 5137 19556 5161 19558
rect 4921 19536 5217 19556
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4986 19408 5042 19417
rect 4540 19366 4844 19394
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4540 16726 4568 18838
rect 4632 18834 4660 19178
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4632 17882 4660 18770
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4632 16538 4660 17546
rect 4724 17270 4752 19246
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4724 16658 4752 17206
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4540 16510 4660 16538
rect 4540 12374 4568 16510
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4632 11694 4660 14894
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12850 4752 13126
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4816 12730 4844 19366
rect 4986 19343 5042 19352
rect 5000 18737 5028 19343
rect 4986 18728 5042 18737
rect 4986 18663 5042 18672
rect 4921 18524 5217 18544
rect 4977 18522 5001 18524
rect 5057 18522 5081 18524
rect 5137 18522 5161 18524
rect 4999 18470 5001 18522
rect 5063 18470 5075 18522
rect 5137 18470 5139 18522
rect 4977 18468 5001 18470
rect 5057 18468 5081 18470
rect 5137 18468 5161 18470
rect 4921 18448 5217 18468
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4908 17610 4936 18090
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4921 17436 5217 17456
rect 4977 17434 5001 17436
rect 5057 17434 5081 17436
rect 5137 17434 5161 17436
rect 4999 17382 5001 17434
rect 5063 17382 5075 17434
rect 5137 17382 5139 17434
rect 4977 17380 5001 17382
rect 5057 17380 5081 17382
rect 5137 17380 5161 17382
rect 4921 17360 5217 17380
rect 4921 16348 5217 16368
rect 4977 16346 5001 16348
rect 5057 16346 5081 16348
rect 5137 16346 5161 16348
rect 4999 16294 5001 16346
rect 5063 16294 5075 16346
rect 5137 16294 5139 16346
rect 4977 16292 5001 16294
rect 5057 16292 5081 16294
rect 5137 16292 5161 16294
rect 4921 16272 5217 16292
rect 5276 15638 5304 22034
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 4921 15260 5217 15280
rect 4977 15258 5001 15260
rect 5057 15258 5081 15260
rect 5137 15258 5161 15260
rect 4999 15206 5001 15258
rect 5063 15206 5075 15258
rect 5137 15206 5139 15258
rect 4977 15204 5001 15206
rect 5057 15204 5081 15206
rect 5137 15204 5161 15206
rect 4921 15184 5217 15204
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5276 14958 5304 15098
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 4921 14172 5217 14192
rect 4977 14170 5001 14172
rect 5057 14170 5081 14172
rect 5137 14170 5161 14172
rect 4999 14118 5001 14170
rect 5063 14118 5075 14170
rect 5137 14118 5139 14170
rect 4977 14116 5001 14118
rect 5057 14116 5081 14118
rect 5137 14116 5161 14118
rect 4921 14096 5217 14116
rect 5276 13462 5304 14350
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 4921 13084 5217 13104
rect 4977 13082 5001 13084
rect 5057 13082 5081 13084
rect 5137 13082 5161 13084
rect 4999 13030 5001 13082
rect 5063 13030 5075 13082
rect 5137 13030 5139 13082
rect 4977 13028 5001 13030
rect 5057 13028 5081 13030
rect 5137 13028 5161 13030
rect 4921 13008 5217 13028
rect 5170 12880 5226 12889
rect 5170 12815 5172 12824
rect 5224 12815 5226 12824
rect 5172 12786 5224 12792
rect 4724 12702 4844 12730
rect 5264 12708 5316 12714
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4434 9072 4490 9081
rect 4434 9007 4490 9016
rect 4356 8758 4660 8786
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4264 7002 4292 8366
rect 4356 7954 4384 8570
rect 4434 8528 4490 8537
rect 4434 8463 4436 8472
rect 4488 8463 4490 8472
rect 4436 8434 4488 8440
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4448 7018 4476 8434
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4540 7546 4568 8298
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4356 6990 4476 7018
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4080 5234 4108 6734
rect 4172 5302 4200 6734
rect 4264 6390 4292 6802
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4252 6248 4304 6254
rect 4356 6236 4384 6990
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4448 6322 4476 6870
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4304 6208 4384 6236
rect 4252 6190 4304 6196
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 3602 4108 5170
rect 4172 4690 4200 5238
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4282 4200 4626
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3194 4108 3538
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4264 2514 4292 6190
rect 4540 6118 4568 7278
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4448 5846 4476 6054
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5370 4384 5714
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4356 800 4384 4966
rect 4448 2310 4476 5646
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4540 2514 4568 3538
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4632 1970 4660 8758
rect 4620 1964 4672 1970
rect 4620 1906 4672 1912
rect 4724 800 4752 12702
rect 5264 12650 5316 12656
rect 4921 11996 5217 12016
rect 4977 11994 5001 11996
rect 5057 11994 5081 11996
rect 5137 11994 5161 11996
rect 4999 11942 5001 11994
rect 5063 11942 5075 11994
rect 5137 11942 5139 11994
rect 4977 11940 5001 11942
rect 5057 11940 5081 11942
rect 5137 11940 5161 11942
rect 4921 11920 5217 11940
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4908 11218 4936 11562
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 5846 4844 11086
rect 4921 10908 5217 10928
rect 4977 10906 5001 10908
rect 5057 10906 5081 10908
rect 5137 10906 5161 10908
rect 4999 10854 5001 10906
rect 5063 10854 5075 10906
rect 5137 10854 5139 10906
rect 4977 10852 5001 10854
rect 5057 10852 5081 10854
rect 5137 10852 5161 10854
rect 4921 10832 5217 10852
rect 4921 9820 5217 9840
rect 4977 9818 5001 9820
rect 5057 9818 5081 9820
rect 5137 9818 5161 9820
rect 4999 9766 5001 9818
rect 5063 9766 5075 9818
rect 5137 9766 5139 9818
rect 4977 9764 5001 9766
rect 5057 9764 5081 9766
rect 5137 9764 5161 9766
rect 4921 9744 5217 9764
rect 5172 9648 5224 9654
rect 4894 9616 4950 9625
rect 5172 9590 5224 9596
rect 4894 9551 4950 9560
rect 4908 9518 4936 9551
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5080 9512 5132 9518
rect 5184 9489 5212 9590
rect 5080 9454 5132 9460
rect 5170 9480 5226 9489
rect 5092 9042 5120 9454
rect 5170 9415 5226 9424
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4921 8732 5217 8752
rect 4977 8730 5001 8732
rect 5057 8730 5081 8732
rect 5137 8730 5161 8732
rect 4999 8678 5001 8730
rect 5063 8678 5075 8730
rect 5137 8678 5139 8730
rect 4977 8676 5001 8678
rect 5057 8676 5081 8678
rect 5137 8676 5161 8678
rect 4921 8656 5217 8676
rect 5276 8650 5304 12650
rect 5368 9110 5396 23015
rect 5460 22556 5488 31583
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 5552 27334 5580 30330
rect 5644 28014 5672 31640
rect 5736 30802 5764 31962
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5828 31686 5856 31826
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5816 30864 5868 30870
rect 5816 30806 5868 30812
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 5724 30116 5776 30122
rect 5724 30058 5776 30064
rect 5736 29850 5764 30058
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 5828 28914 5856 30806
rect 5920 30666 5948 32184
rect 5908 30660 5960 30666
rect 5908 30602 5960 30608
rect 5908 30116 5960 30122
rect 5908 30058 5960 30064
rect 5736 28886 5856 28914
rect 5632 28008 5684 28014
rect 5632 27950 5684 27956
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5644 25770 5672 27950
rect 5632 25764 5684 25770
rect 5632 25706 5684 25712
rect 5736 25498 5764 28886
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5828 26450 5856 28698
rect 5920 27946 5948 30058
rect 5908 27940 5960 27946
rect 5908 27882 5960 27888
rect 6012 26586 6040 33510
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 6000 26444 6052 26450
rect 6000 26386 6052 26392
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 5736 24886 5764 25434
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 5816 24880 5868 24886
rect 5816 24822 5868 24828
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5552 23662 5580 24346
rect 5828 23798 5856 24822
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5552 22658 5580 23598
rect 5552 22630 5672 22658
rect 5644 22574 5672 22630
rect 5632 22568 5684 22574
rect 5460 22528 5580 22556
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5460 19446 5488 21966
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5552 19258 5580 22528
rect 5632 22510 5684 22516
rect 5828 21554 5856 23598
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5724 21412 5776 21418
rect 5724 21354 5776 21360
rect 5736 19922 5764 21354
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5460 19230 5580 19258
rect 5460 15162 5488 19230
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17814 5580 18022
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5644 17134 5672 18702
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5736 17202 5764 17614
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5552 15570 5580 16730
rect 5540 15564 5592 15570
rect 5592 15524 5672 15552
rect 5540 15506 5592 15512
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14278 5488 14894
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5446 13832 5502 13841
rect 5446 13767 5502 13776
rect 5460 12102 5488 13767
rect 5552 13394 5580 14758
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5460 10810 5488 11222
rect 5552 10810 5580 13194
rect 5644 12850 5672 15524
rect 5828 13326 5856 21490
rect 5920 19854 5948 23054
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 19514 5948 19790
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5920 18086 5948 19450
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5920 17542 5948 18022
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 14958 5948 17478
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 13938 5948 14282
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5460 9466 5488 10746
rect 5736 10146 5764 12174
rect 5552 10118 5764 10146
rect 5552 9602 5580 10118
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5644 9738 5672 9998
rect 5644 9722 5764 9738
rect 5644 9716 5776 9722
rect 5644 9710 5724 9716
rect 5724 9658 5776 9664
rect 5920 9625 5948 13874
rect 5906 9616 5962 9625
rect 5552 9574 5764 9602
rect 5630 9480 5686 9489
rect 5460 9438 5580 9466
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5460 9042 5488 9318
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5276 8622 5488 8650
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4921 7644 5217 7664
rect 4977 7642 5001 7644
rect 5057 7642 5081 7644
rect 5137 7642 5161 7644
rect 4999 7590 5001 7642
rect 5063 7590 5075 7642
rect 5137 7590 5139 7642
rect 4977 7588 5001 7590
rect 5057 7588 5081 7590
rect 5137 7588 5161 7590
rect 4921 7568 5217 7588
rect 5276 7342 5304 7890
rect 5368 7886 5396 8502
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5092 6730 5120 7210
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4921 6556 5217 6576
rect 4977 6554 5001 6556
rect 5057 6554 5081 6556
rect 5137 6554 5161 6556
rect 4999 6502 5001 6554
rect 5063 6502 5075 6554
rect 5137 6502 5139 6554
rect 4977 6500 5001 6502
rect 5057 6500 5081 6502
rect 5137 6500 5161 6502
rect 4921 6480 5217 6500
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 6118 5028 6190
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4908 5658 4936 5850
rect 5000 5794 5028 6054
rect 5276 5914 5304 7278
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5846 5396 7822
rect 5460 7410 5488 8622
rect 5552 8430 5580 9438
rect 5630 9415 5686 9424
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6934 5488 7346
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5552 6866 5580 8366
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 5840 5408 5846
rect 5000 5766 5304 5794
rect 5356 5782 5408 5788
rect 4816 5630 4936 5658
rect 4816 4690 4844 5630
rect 4921 5468 5217 5488
rect 4977 5466 5001 5468
rect 5057 5466 5081 5468
rect 5137 5466 5161 5468
rect 4999 5414 5001 5466
rect 5063 5414 5075 5466
rect 5137 5414 5139 5466
rect 4977 5412 5001 5414
rect 5057 5412 5081 5414
rect 5137 5412 5161 5414
rect 4921 5392 5217 5412
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 3738 4844 4626
rect 5184 4570 5212 5238
rect 5276 5098 5304 5766
rect 5368 5642 5396 5782
rect 5460 5710 5488 6598
rect 5644 6322 5672 9415
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5166 5396 5578
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5460 4978 5488 5646
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5552 5302 5580 5578
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5368 4950 5488 4978
rect 5368 4690 5396 4950
rect 5552 4758 5580 5102
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5184 4542 5304 4570
rect 4921 4380 5217 4400
rect 4977 4378 5001 4380
rect 5057 4378 5081 4380
rect 5137 4378 5161 4380
rect 4999 4326 5001 4378
rect 5063 4326 5075 4378
rect 5137 4326 5139 4378
rect 4977 4324 5001 4326
rect 5057 4324 5081 4326
rect 5137 4324 5161 4326
rect 4921 4304 5217 4324
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4816 3058 4844 3674
rect 4921 3292 5217 3312
rect 4977 3290 5001 3292
rect 5057 3290 5081 3292
rect 5137 3290 5161 3292
rect 4999 3238 5001 3290
rect 5063 3238 5075 3290
rect 5137 3238 5139 3290
rect 4977 3236 5001 3238
rect 5057 3236 5081 3238
rect 5137 3236 5161 3238
rect 4921 3216 5217 3236
rect 5276 3194 5304 4542
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5368 2922 5396 4626
rect 5644 4622 5672 5510
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5736 4078 5764 9574
rect 5816 9580 5868 9586
rect 5906 9551 5962 9560
rect 5816 9522 5868 9528
rect 5724 4072 5776 4078
rect 5644 4020 5724 4026
rect 5644 4014 5776 4020
rect 5644 3998 5764 4014
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5368 2582 5396 2858
rect 5644 2582 5672 3998
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3602 5764 3878
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 4921 2204 5217 2224
rect 4977 2202 5001 2204
rect 5057 2202 5081 2204
rect 5137 2202 5161 2204
rect 4999 2150 5001 2202
rect 5063 2150 5075 2202
rect 5137 2150 5139 2202
rect 4977 2148 5001 2150
rect 5057 2148 5081 2150
rect 5137 2148 5161 2150
rect 4921 2128 5217 2148
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 5092 800 5120 1906
rect 5446 1864 5502 1873
rect 5446 1799 5502 1808
rect 5460 800 5488 1799
rect 5828 800 5856 9522
rect 5920 6934 5948 9551
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 5778 5948 6734
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5098 5948 5714
rect 6012 5302 6040 26386
rect 6104 13530 6132 33918
rect 6184 33448 6236 33454
rect 6184 33390 6236 33396
rect 6196 32910 6224 33390
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6196 31906 6224 32846
rect 6196 31890 6316 31906
rect 6196 31884 6328 31890
rect 6196 31878 6276 31884
rect 6276 31826 6328 31832
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 6196 30938 6224 31758
rect 6184 30932 6236 30938
rect 6184 30874 6236 30880
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 28626 6224 29446
rect 6184 28620 6236 28626
rect 6184 28562 6236 28568
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 6288 27130 6316 27406
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 19446 6224 22510
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6196 17746 6224 19246
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6196 16250 6224 17682
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6196 13410 6224 16050
rect 6104 13382 6224 13410
rect 6104 11626 6132 13382
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6104 9625 6132 11562
rect 6196 11014 6224 13262
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6090 9616 6146 9625
rect 6090 9551 6146 9560
rect 6104 8294 6132 9551
rect 6196 9518 6224 10950
rect 6288 9586 6316 27066
rect 6380 18154 6408 37742
rect 6460 36372 6512 36378
rect 6460 36314 6512 36320
rect 6472 36242 6500 36314
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 6472 34746 6500 36178
rect 6460 34740 6512 34746
rect 6460 34682 6512 34688
rect 6460 34604 6512 34610
rect 6460 34546 6512 34552
rect 6472 32910 6500 34546
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6460 32360 6512 32366
rect 6460 32302 6512 32308
rect 6472 30802 6500 32302
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6460 30184 6512 30190
rect 6460 30126 6512 30132
rect 6472 28422 6500 30126
rect 6460 28416 6512 28422
rect 6460 28358 6512 28364
rect 6472 26858 6500 28358
rect 6460 26852 6512 26858
rect 6460 26794 6512 26800
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 6472 18970 6500 26182
rect 6564 21593 6592 39374
rect 6644 38412 6696 38418
rect 6644 38354 6696 38360
rect 6550 21584 6606 21593
rect 6550 21519 6606 21528
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6564 21078 6592 21422
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6552 19440 6604 19446
rect 6552 19382 6604 19388
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6472 16794 6500 18906
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6380 12986 6408 15982
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6380 11694 6408 12922
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6472 9058 6500 16594
rect 6564 13870 6592 19382
rect 6656 15638 6684 38354
rect 6748 38010 6776 40530
rect 6840 39574 6868 41074
rect 7024 41070 7052 42162
rect 7196 41608 7248 41614
rect 7196 41550 7248 41556
rect 7012 41064 7064 41070
rect 7012 41006 7064 41012
rect 6828 39568 6880 39574
rect 6828 39510 6880 39516
rect 7024 39302 7052 41006
rect 7208 40526 7236 41550
rect 7392 41274 7420 43182
rect 7484 42226 7512 43982
rect 7656 43852 7708 43858
rect 7656 43794 7708 43800
rect 7564 43784 7616 43790
rect 7564 43726 7616 43732
rect 7472 42220 7524 42226
rect 7472 42162 7524 42168
rect 7472 41676 7524 41682
rect 7472 41618 7524 41624
rect 7380 41268 7432 41274
rect 7380 41210 7432 41216
rect 7288 41064 7340 41070
rect 7288 41006 7340 41012
rect 7300 40662 7328 41006
rect 7288 40656 7340 40662
rect 7288 40598 7340 40604
rect 7196 40520 7248 40526
rect 7196 40462 7248 40468
rect 7012 39296 7064 39302
rect 7012 39238 7064 39244
rect 7484 38962 7512 41618
rect 7472 38956 7524 38962
rect 7472 38898 7524 38904
rect 6828 38888 6880 38894
rect 6828 38830 6880 38836
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6840 35306 6868 38830
rect 7576 38418 7604 43726
rect 7668 42566 7696 43794
rect 7760 43654 7788 45358
rect 7932 44328 7984 44334
rect 7932 44270 7984 44276
rect 7944 43654 7972 44270
rect 8128 43926 8156 47246
rect 8208 47116 8260 47122
rect 8208 47058 8260 47064
rect 8220 46102 8248 47058
rect 8760 46504 8812 46510
rect 8760 46446 8812 46452
rect 8208 46096 8260 46102
rect 8208 46038 8260 46044
rect 8220 43994 8248 46038
rect 8484 45824 8536 45830
rect 8484 45766 8536 45772
rect 8496 45422 8524 45766
rect 8772 45626 8800 46446
rect 8886 46268 9182 46288
rect 8942 46266 8966 46268
rect 9022 46266 9046 46268
rect 9102 46266 9126 46268
rect 8964 46214 8966 46266
rect 9028 46214 9040 46266
rect 9102 46214 9104 46266
rect 8942 46212 8966 46214
rect 9022 46212 9046 46214
rect 9102 46212 9126 46214
rect 8886 46192 9182 46212
rect 8760 45620 8812 45626
rect 8760 45562 8812 45568
rect 8484 45416 8536 45422
rect 8484 45358 8536 45364
rect 8392 45348 8444 45354
rect 8392 45290 8444 45296
rect 8208 43988 8260 43994
rect 8208 43930 8260 43936
rect 8116 43920 8168 43926
rect 8116 43862 8168 43868
rect 7748 43648 7800 43654
rect 7748 43590 7800 43596
rect 7932 43648 7984 43654
rect 7932 43590 7984 43596
rect 8220 43246 8248 43930
rect 8208 43240 8260 43246
rect 8208 43182 8260 43188
rect 7748 43104 7800 43110
rect 7748 43046 7800 43052
rect 7656 42560 7708 42566
rect 7656 42502 7708 42508
rect 7760 41750 7788 43046
rect 8220 42838 8248 43182
rect 8208 42832 8260 42838
rect 8208 42774 8260 42780
rect 7840 42152 7892 42158
rect 7840 42094 7892 42100
rect 7748 41744 7800 41750
rect 7748 41686 7800 41692
rect 7852 41478 7880 42094
rect 7840 41472 7892 41478
rect 7840 41414 7892 41420
rect 8208 40588 8260 40594
rect 8208 40530 8260 40536
rect 7748 39908 7800 39914
rect 7748 39850 7800 39856
rect 7760 39506 7788 39850
rect 7748 39500 7800 39506
rect 7748 39442 7800 39448
rect 7656 38888 7708 38894
rect 7656 38830 7708 38836
rect 7668 38418 7696 38830
rect 7760 38554 7788 39442
rect 7840 39296 7892 39302
rect 7840 39238 7892 39244
rect 7748 38548 7800 38554
rect 7748 38490 7800 38496
rect 7564 38412 7616 38418
rect 7564 38354 7616 38360
rect 7656 38412 7708 38418
rect 7656 38354 7708 38360
rect 7668 37806 7696 38354
rect 7852 37874 7880 39238
rect 7930 38992 7986 39001
rect 7930 38927 7986 38936
rect 7840 37868 7892 37874
rect 7840 37810 7892 37816
rect 7656 37800 7708 37806
rect 7656 37742 7708 37748
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 7564 37324 7616 37330
rect 7564 37266 7616 37272
rect 7116 36922 7144 37266
rect 7104 36916 7156 36922
rect 7104 36858 7156 36864
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 6932 36310 6960 36654
rect 6920 36304 6972 36310
rect 6920 36246 6972 36252
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7392 35766 7420 36110
rect 7380 35760 7432 35766
rect 7380 35702 7432 35708
rect 7012 35488 7064 35494
rect 7012 35430 7064 35436
rect 6748 35278 6868 35306
rect 7024 35290 7052 35430
rect 7012 35284 7064 35290
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6564 11830 6592 13806
rect 6656 13394 6684 15438
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12374 6684 13330
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 10606 6592 11494
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6196 9030 6500 9058
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 6104 800 6132 6258
rect 6196 4570 6224 9030
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 5846 6408 8366
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6472 4690 6500 8842
rect 6564 7954 6592 10542
rect 6656 10130 6684 11698
rect 6748 11354 6776 35278
rect 7012 35226 7064 35232
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 6840 28762 6868 34682
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6840 27606 6868 28494
rect 6828 27600 6880 27606
rect 6828 27542 6880 27548
rect 6932 27538 6960 29990
rect 7024 29102 7052 30670
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 7024 27674 7052 29038
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 7024 27538 7052 27610
rect 6920 27532 6972 27538
rect 6920 27474 6972 27480
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6840 27130 6868 27270
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 26246 6868 26862
rect 6932 26586 6960 27474
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 7024 26466 7052 26726
rect 6932 26438 7052 26466
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6932 24410 6960 26438
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 7024 24750 7052 26318
rect 7116 25702 7144 32234
rect 7208 30870 7236 33798
rect 7300 31804 7328 35022
rect 7576 34542 7604 37266
rect 7944 36718 7972 38927
rect 8024 37732 8076 37738
rect 8024 37674 8076 37680
rect 8036 37466 8064 37674
rect 8024 37460 8076 37466
rect 8024 37402 8076 37408
rect 8036 37330 8064 37402
rect 8024 37324 8076 37330
rect 8024 37266 8076 37272
rect 8116 37120 8168 37126
rect 8116 37062 8168 37068
rect 8128 36922 8156 37062
rect 8116 36916 8168 36922
rect 8116 36858 8168 36864
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 8128 35222 8156 36858
rect 8116 35216 8168 35222
rect 8116 35158 8168 35164
rect 7472 34536 7524 34542
rect 7472 34478 7524 34484
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 7484 34202 7512 34478
rect 7748 34400 7800 34406
rect 7748 34342 7800 34348
rect 7472 34196 7524 34202
rect 7472 34138 7524 34144
rect 7380 33108 7432 33114
rect 7380 33050 7432 33056
rect 7392 31958 7420 33050
rect 7484 32434 7512 34138
rect 7760 33522 7788 34342
rect 7748 33516 7800 33522
rect 7748 33458 7800 33464
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 8024 32428 8076 32434
rect 8024 32370 8076 32376
rect 7932 32292 7984 32298
rect 7932 32234 7984 32240
rect 7944 32026 7972 32234
rect 7932 32020 7984 32026
rect 7932 31962 7984 31968
rect 7380 31952 7432 31958
rect 7380 31894 7432 31900
rect 7300 31776 7512 31804
rect 7196 30864 7248 30870
rect 7196 30806 7248 30812
rect 7196 30592 7248 30598
rect 7196 30534 7248 30540
rect 7208 29714 7236 30534
rect 7380 30116 7432 30122
rect 7380 30058 7432 30064
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 7196 29096 7248 29102
rect 7196 29038 7248 29044
rect 7208 28150 7236 29038
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7196 28144 7248 28150
rect 7196 28086 7248 28092
rect 7300 26518 7328 28358
rect 7288 26512 7340 26518
rect 7288 26454 7340 26460
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 22574 6868 24142
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22409 6868 22510
rect 6826 22400 6882 22409
rect 6826 22335 6882 22344
rect 6932 22114 6960 24210
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 7024 23662 7052 24006
rect 7116 23866 7144 25298
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6840 22086 6960 22114
rect 6840 21962 6868 22086
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 6840 20942 6868 21898
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20806 6868 20837
rect 6828 20800 6880 20806
rect 6826 20768 6828 20777
rect 6880 20768 6882 20777
rect 6826 20703 6882 20712
rect 6840 18290 6868 20703
rect 6932 20330 6960 21422
rect 7024 20346 7052 23462
rect 7116 22778 7144 23598
rect 7208 23066 7236 24686
rect 7300 23526 7328 26454
rect 7392 25158 7420 30058
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 7392 24274 7420 25094
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7392 23186 7420 23530
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7208 23038 7420 23066
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7194 22400 7250 22409
rect 7116 21010 7144 22374
rect 7194 22335 7250 22344
rect 7208 22166 7236 22335
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7116 20534 7144 20810
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7208 20466 7236 22102
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 21010 7328 21966
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 6920 20324 6972 20330
rect 7024 20318 7236 20346
rect 6920 20266 6972 20272
rect 6932 20058 6960 20266
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6918 19952 6974 19961
rect 6918 19887 6974 19896
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6840 16114 6868 18226
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6932 15722 6960 19887
rect 7024 19310 7052 20198
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 17882 7052 19246
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 7024 16046 7052 17546
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 6932 15694 7052 15722
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13938 6868 14214
rect 7024 14074 7052 15694
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12986 7052 13330
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6840 11354 6868 11766
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6932 11218 6960 12310
rect 7024 12306 7052 12922
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7024 11098 7052 11630
rect 6932 11070 7052 11098
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 8956 6684 10066
rect 6932 9042 6960 11070
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10198 7052 10406
rect 7116 10305 7144 15982
rect 7208 15570 7236 20318
rect 7300 18834 7328 20946
rect 7392 19174 7420 23038
rect 7484 22001 7512 31776
rect 8036 31686 8064 32370
rect 8116 32360 8168 32366
rect 8116 32302 8168 32308
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 8036 31278 8064 31622
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 8036 30666 8064 31214
rect 8024 30660 8076 30666
rect 8024 30602 8076 30608
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7564 28008 7616 28014
rect 7564 27950 7616 27956
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7576 26790 7604 27950
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26926 7696 27270
rect 7760 26994 7788 27950
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7564 26784 7616 26790
rect 7564 26726 7616 26732
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 7576 24274 7604 26386
rect 7668 25430 7696 26386
rect 7852 25838 7880 30534
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 8036 29782 8064 30126
rect 8024 29776 8076 29782
rect 8024 29718 8076 29724
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 8036 29306 8064 29582
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8024 28076 8076 28082
rect 8024 28018 8076 28024
rect 8036 26926 8064 28018
rect 8024 26920 8076 26926
rect 7944 26880 8024 26908
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7656 25424 7708 25430
rect 7656 25366 7708 25372
rect 7760 24818 7788 25706
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7852 24614 7880 24754
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7944 24392 7972 26880
rect 8024 26862 8076 26868
rect 8024 26308 8076 26314
rect 8024 26250 8076 26256
rect 8036 26042 8064 26250
rect 8024 26036 8076 26042
rect 8024 25978 8076 25984
rect 8024 25696 8076 25702
rect 8024 25638 8076 25644
rect 7760 24364 7972 24392
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7576 22817 7604 22918
rect 7562 22808 7618 22817
rect 7562 22743 7618 22752
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7470 21992 7526 22001
rect 7470 21927 7526 21936
rect 7576 21894 7604 22442
rect 7564 21888 7616 21894
rect 7470 21856 7526 21865
rect 7564 21830 7616 21836
rect 7470 21791 7526 21800
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7378 19000 7434 19009
rect 7378 18935 7434 18944
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7392 18766 7420 18935
rect 7484 18766 7512 21791
rect 7576 21729 7604 21830
rect 7562 21720 7618 21729
rect 7562 21655 7618 21664
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7576 20788 7604 21558
rect 7668 21350 7696 22510
rect 7760 21593 7788 24364
rect 8036 24290 8064 25638
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 7944 24262 8064 24290
rect 7746 21584 7802 21593
rect 7746 21519 7748 21528
rect 7800 21519 7802 21528
rect 7748 21490 7800 21496
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7668 20942 7696 21286
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7576 20760 7696 20788
rect 7564 20324 7616 20330
rect 7564 20266 7616 20272
rect 7380 18760 7432 18766
rect 7300 18708 7380 18714
rect 7300 18702 7432 18708
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7300 18686 7420 18702
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7300 15450 7328 18686
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 16114 7420 17682
rect 7484 17270 7512 18158
rect 7576 18154 7604 20266
rect 7668 18970 7696 20760
rect 7760 20058 7788 20878
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19514 7788 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16658 7512 17070
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7208 15422 7328 15450
rect 7102 10296 7158 10305
rect 7102 10231 7158 10240
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6736 8968 6788 8974
rect 6656 8928 6736 8956
rect 6736 8910 6788 8916
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6748 7750 6776 8910
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6932 8022 6960 8502
rect 7024 8294 7052 9998
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7410 6776 7686
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6866 6776 7346
rect 6920 7200 6972 7206
rect 7024 7188 7052 8230
rect 7116 7818 7144 10134
rect 7208 8566 7236 15422
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7300 7970 7328 14350
rect 7392 10742 7420 15914
rect 7484 14006 7512 16594
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7392 10470 7420 10678
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7484 10198 7512 13330
rect 7668 12322 7696 18634
rect 7760 17202 7788 19178
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7852 15570 7880 24210
rect 7944 22817 7972 24262
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7930 22808 7986 22817
rect 7930 22743 7986 22752
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7944 21010 7972 22578
rect 8036 22098 8064 24142
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 8036 20074 8064 22034
rect 8128 21622 8156 32302
rect 8220 27674 8248 40530
rect 8404 39506 8432 45290
rect 8886 45180 9182 45200
rect 8942 45178 8966 45180
rect 9022 45178 9046 45180
rect 9102 45178 9126 45180
rect 8964 45126 8966 45178
rect 9028 45126 9040 45178
rect 9102 45126 9104 45178
rect 8942 45124 8966 45126
rect 9022 45124 9046 45126
rect 9102 45124 9126 45126
rect 8886 45104 9182 45124
rect 9220 44940 9272 44946
rect 9220 44882 9272 44888
rect 8886 44092 9182 44112
rect 8942 44090 8966 44092
rect 9022 44090 9046 44092
rect 9102 44090 9126 44092
rect 8964 44038 8966 44090
rect 9028 44038 9040 44090
rect 9102 44038 9104 44090
rect 8942 44036 8966 44038
rect 9022 44036 9046 44038
rect 9102 44036 9126 44038
rect 8886 44016 9182 44036
rect 8886 43004 9182 43024
rect 8942 43002 8966 43004
rect 9022 43002 9046 43004
rect 9102 43002 9126 43004
rect 8964 42950 8966 43002
rect 9028 42950 9040 43002
rect 9102 42950 9104 43002
rect 8942 42948 8966 42950
rect 9022 42948 9046 42950
rect 9102 42948 9126 42950
rect 8886 42928 9182 42948
rect 8886 41916 9182 41936
rect 8942 41914 8966 41916
rect 9022 41914 9046 41916
rect 9102 41914 9126 41916
rect 8964 41862 8966 41914
rect 9028 41862 9040 41914
rect 9102 41862 9104 41914
rect 8942 41860 8966 41862
rect 9022 41860 9046 41862
rect 9102 41860 9126 41862
rect 8886 41840 9182 41860
rect 8886 40828 9182 40848
rect 8942 40826 8966 40828
rect 9022 40826 9046 40828
rect 9102 40826 9126 40828
rect 8964 40774 8966 40826
rect 9028 40774 9040 40826
rect 9102 40774 9104 40826
rect 8942 40772 8966 40774
rect 9022 40772 9046 40774
rect 9102 40772 9126 40774
rect 8886 40752 9182 40772
rect 8760 40588 8812 40594
rect 8760 40530 8812 40536
rect 8772 39982 8800 40530
rect 9232 40186 9260 44882
rect 9324 43314 9352 47518
rect 9784 44538 9812 49200
rect 10048 46912 10100 46918
rect 10048 46854 10100 46860
rect 10060 45014 10088 46854
rect 10612 46714 10640 49200
rect 11244 47252 11296 47258
rect 11244 47194 11296 47200
rect 10600 46708 10652 46714
rect 10600 46650 10652 46656
rect 10612 46034 10640 46650
rect 11152 46504 11204 46510
rect 11152 46446 11204 46452
rect 10600 46028 10652 46034
rect 10600 45970 10652 45976
rect 10784 46028 10836 46034
rect 10784 45970 10836 45976
rect 10796 45490 10824 45970
rect 10968 45960 11020 45966
rect 10968 45902 11020 45908
rect 10784 45484 10836 45490
rect 10784 45426 10836 45432
rect 10140 45416 10192 45422
rect 10140 45358 10192 45364
rect 10048 45008 10100 45014
rect 10048 44950 10100 44956
rect 10152 44742 10180 45358
rect 10140 44736 10192 44742
rect 10140 44678 10192 44684
rect 10980 44538 11008 45902
rect 9772 44532 9824 44538
rect 9772 44474 9824 44480
rect 10968 44532 11020 44538
rect 10968 44474 11020 44480
rect 9312 43308 9364 43314
rect 9312 43250 9364 43256
rect 9324 42362 9352 43250
rect 9496 43172 9548 43178
rect 9496 43114 9548 43120
rect 9312 42356 9364 42362
rect 9312 42298 9364 42304
rect 9508 41750 9536 43114
rect 9588 42764 9640 42770
rect 9784 42752 9812 44474
rect 10416 44328 10468 44334
rect 10416 44270 10468 44276
rect 9640 42724 9812 42752
rect 9588 42706 9640 42712
rect 9956 42696 10008 42702
rect 9956 42638 10008 42644
rect 9496 41744 9548 41750
rect 9496 41686 9548 41692
rect 9680 41676 9732 41682
rect 9680 41618 9732 41624
rect 9692 40526 9720 41618
rect 9968 41478 9996 42638
rect 9956 41472 10008 41478
rect 9956 41414 10008 41420
rect 9864 41064 9916 41070
rect 9864 41006 9916 41012
rect 9876 40594 9904 41006
rect 9864 40588 9916 40594
rect 9864 40530 9916 40536
rect 9680 40520 9732 40526
rect 9680 40462 9732 40468
rect 10048 40384 10100 40390
rect 10048 40326 10100 40332
rect 9220 40180 9272 40186
rect 9220 40122 9272 40128
rect 8760 39976 8812 39982
rect 8760 39918 8812 39924
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 9864 39976 9916 39982
rect 9864 39918 9916 39924
rect 8772 39506 8800 39918
rect 8886 39740 9182 39760
rect 8942 39738 8966 39740
rect 9022 39738 9046 39740
rect 9102 39738 9126 39740
rect 8964 39686 8966 39738
rect 9028 39686 9040 39738
rect 9102 39686 9104 39738
rect 8942 39684 8966 39686
rect 9022 39684 9046 39686
rect 9102 39684 9126 39686
rect 8886 39664 9182 39684
rect 8392 39500 8444 39506
rect 8392 39442 8444 39448
rect 8760 39500 8812 39506
rect 8760 39442 8812 39448
rect 8392 39364 8444 39370
rect 8392 39306 8444 39312
rect 8300 34672 8352 34678
rect 8300 34614 8352 34620
rect 8312 34066 8340 34614
rect 8300 34060 8352 34066
rect 8300 34002 8352 34008
rect 8312 31890 8340 34002
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8312 28529 8340 28562
rect 8298 28520 8354 28529
rect 8298 28455 8354 28464
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8208 27668 8260 27674
rect 8208 27610 8260 27616
rect 8312 27316 8340 27814
rect 8404 27470 8432 39306
rect 8760 38752 8812 38758
rect 8760 38694 8812 38700
rect 8772 38486 8800 38694
rect 8886 38652 9182 38672
rect 8942 38650 8966 38652
rect 9022 38650 9046 38652
rect 9102 38650 9126 38652
rect 8964 38598 8966 38650
rect 9028 38598 9040 38650
rect 9102 38598 9104 38650
rect 8942 38596 8966 38598
rect 9022 38596 9046 38598
rect 9102 38596 9126 38598
rect 8886 38576 9182 38596
rect 8760 38480 8812 38486
rect 8760 38422 8812 38428
rect 8668 38412 8720 38418
rect 8668 38354 8720 38360
rect 8680 36564 8708 38354
rect 8772 38214 8800 38422
rect 8760 38208 8812 38214
rect 8760 38150 8812 38156
rect 8760 37800 8812 37806
rect 8760 37742 8812 37748
rect 8772 37398 8800 37742
rect 8886 37564 9182 37584
rect 8942 37562 8966 37564
rect 9022 37562 9046 37564
rect 9102 37562 9126 37564
rect 8964 37510 8966 37562
rect 9028 37510 9040 37562
rect 9102 37510 9104 37562
rect 8942 37508 8966 37510
rect 9022 37508 9046 37510
rect 9102 37508 9126 37510
rect 8886 37488 9182 37508
rect 8760 37392 8812 37398
rect 8760 37334 8812 37340
rect 8760 36576 8812 36582
rect 8680 36536 8760 36564
rect 8760 36518 8812 36524
rect 8668 36168 8720 36174
rect 8668 36110 8720 36116
rect 8680 35630 8708 36110
rect 8668 35624 8720 35630
rect 8668 35566 8720 35572
rect 8484 35556 8536 35562
rect 8484 35498 8536 35504
rect 8496 34542 8524 35498
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8496 34202 8524 34478
rect 8484 34196 8536 34202
rect 8484 34138 8536 34144
rect 8772 33318 8800 36518
rect 8886 36476 9182 36496
rect 8942 36474 8966 36476
rect 9022 36474 9046 36476
rect 9102 36474 9126 36476
rect 8964 36422 8966 36474
rect 9028 36422 9040 36474
rect 9102 36422 9104 36474
rect 8942 36420 8966 36422
rect 9022 36420 9046 36422
rect 9102 36420 9126 36422
rect 8886 36400 9182 36420
rect 8852 36032 8904 36038
rect 8852 35974 8904 35980
rect 8864 35834 8892 35974
rect 8852 35828 8904 35834
rect 8852 35770 8904 35776
rect 8864 35562 8892 35770
rect 8852 35556 8904 35562
rect 8852 35498 8904 35504
rect 8886 35388 9182 35408
rect 8942 35386 8966 35388
rect 9022 35386 9046 35388
rect 9102 35386 9126 35388
rect 8964 35334 8966 35386
rect 9028 35334 9040 35386
rect 9102 35334 9104 35386
rect 8942 35332 8966 35334
rect 9022 35332 9046 35334
rect 9102 35332 9126 35334
rect 8886 35312 9182 35332
rect 8886 34300 9182 34320
rect 8942 34298 8966 34300
rect 9022 34298 9046 34300
rect 9102 34298 9126 34300
rect 8964 34246 8966 34298
rect 9028 34246 9040 34298
rect 9102 34246 9104 34298
rect 8942 34244 8966 34246
rect 9022 34244 9046 34246
rect 9102 34244 9126 34246
rect 8886 34224 9182 34244
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8886 33212 9182 33232
rect 8942 33210 8966 33212
rect 9022 33210 9046 33212
rect 9102 33210 9126 33212
rect 8964 33158 8966 33210
rect 9028 33158 9040 33210
rect 9102 33158 9104 33210
rect 8942 33156 8966 33158
rect 9022 33156 9046 33158
rect 9102 33156 9126 33158
rect 8886 33136 9182 33156
rect 9232 32230 9260 39918
rect 9876 39506 9904 39918
rect 9864 39500 9916 39506
rect 9864 39442 9916 39448
rect 9588 39024 9640 39030
rect 9586 38992 9588 39001
rect 9640 38992 9642 39001
rect 9586 38927 9642 38936
rect 9876 38894 9904 39442
rect 10060 39030 10088 40326
rect 10428 40186 10456 44270
rect 10508 43648 10560 43654
rect 10508 43590 10560 43596
rect 10520 43178 10548 43590
rect 10600 43240 10652 43246
rect 10600 43182 10652 43188
rect 10508 43172 10560 43178
rect 10508 43114 10560 43120
rect 10416 40180 10468 40186
rect 10416 40122 10468 40128
rect 10232 39908 10284 39914
rect 10232 39850 10284 39856
rect 10048 39024 10100 39030
rect 10048 38966 10100 38972
rect 9864 38888 9916 38894
rect 9864 38830 9916 38836
rect 9876 38554 9904 38830
rect 9864 38548 9916 38554
rect 9864 38490 9916 38496
rect 10048 37664 10100 37670
rect 10048 37606 10100 37612
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9692 35494 9720 36722
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9784 36582 9812 36654
rect 9772 36576 9824 36582
rect 9772 36518 9824 36524
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 9312 34740 9364 34746
rect 9312 34682 9364 34688
rect 9324 34542 9352 34682
rect 9692 34626 9720 35430
rect 9600 34598 9720 34626
rect 9312 34536 9364 34542
rect 9312 34478 9364 34484
rect 9220 32224 9272 32230
rect 9220 32166 9272 32172
rect 8886 32124 9182 32144
rect 8942 32122 8966 32124
rect 9022 32122 9046 32124
rect 9102 32122 9126 32124
rect 8964 32070 8966 32122
rect 9028 32070 9040 32122
rect 9102 32070 9104 32122
rect 8942 32068 8966 32070
rect 9022 32068 9046 32070
rect 9102 32068 9126 32070
rect 8886 32048 9182 32068
rect 8760 31816 8812 31822
rect 8760 31758 8812 31764
rect 8772 30258 8800 31758
rect 9220 31204 9272 31210
rect 9220 31146 9272 31152
rect 8886 31036 9182 31056
rect 8942 31034 8966 31036
rect 9022 31034 9046 31036
rect 9102 31034 9126 31036
rect 8964 30982 8966 31034
rect 9028 30982 9040 31034
rect 9102 30982 9104 31034
rect 8942 30980 8966 30982
rect 9022 30980 9046 30982
rect 9102 30980 9126 30982
rect 8886 30960 9182 30980
rect 8760 30252 8812 30258
rect 8760 30194 8812 30200
rect 9232 30190 9260 31146
rect 9220 30184 9272 30190
rect 9220 30126 9272 30132
rect 8668 30116 8720 30122
rect 8668 30058 8720 30064
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8312 27288 8432 27316
rect 8496 27305 8524 27610
rect 8404 27112 8432 27288
rect 8482 27296 8538 27305
rect 8482 27231 8538 27240
rect 8404 27084 8524 27112
rect 8300 27056 8352 27062
rect 8298 27024 8300 27033
rect 8352 27024 8354 27033
rect 8298 26959 8354 26968
rect 8300 26920 8352 26926
rect 8496 26908 8524 27084
rect 8352 26880 8524 26908
rect 8300 26862 8352 26868
rect 8208 26852 8260 26858
rect 8208 26794 8260 26800
rect 8220 26586 8248 26794
rect 8300 26784 8352 26790
rect 8298 26752 8300 26761
rect 8392 26784 8444 26790
rect 8352 26752 8354 26761
rect 8392 26726 8444 26732
rect 8298 26687 8354 26696
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 8220 24206 8248 25162
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8312 23526 8340 24210
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8312 23322 8340 23462
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8206 22128 8262 22137
rect 8206 22063 8262 22072
rect 8116 21616 8168 21622
rect 8116 21558 8168 21564
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 7944 20046 8064 20074
rect 8128 20058 8156 21354
rect 8220 20534 8248 22063
rect 8404 20924 8432 26726
rect 8588 25770 8616 29446
rect 8680 28150 8708 30058
rect 8886 29948 9182 29968
rect 8942 29946 8966 29948
rect 9022 29946 9046 29948
rect 9102 29946 9126 29948
rect 8964 29894 8966 29946
rect 9028 29894 9040 29946
rect 9102 29894 9104 29946
rect 8942 29892 8966 29894
rect 9022 29892 9046 29894
rect 9102 29892 9126 29894
rect 8886 29872 9182 29892
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 8680 27033 8708 27270
rect 8666 27024 8722 27033
rect 8666 26959 8722 26968
rect 8666 26752 8722 26761
rect 8666 26687 8722 26696
rect 8680 26586 8708 26687
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8588 24750 8616 25298
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8588 24410 8616 24686
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8482 22672 8538 22681
rect 8482 22607 8538 22616
rect 8496 22574 8524 22607
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8496 22234 8524 22510
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8496 21078 8524 21558
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8404 20896 8524 20924
rect 8390 20768 8446 20777
rect 8390 20703 8446 20712
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8116 20052 8168 20058
rect 7944 17678 7972 20046
rect 8116 19994 8168 20000
rect 8404 19990 8432 20703
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 8036 17542 8064 19858
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8128 19514 8156 19722
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8220 19174 8248 19858
rect 8390 19816 8446 19825
rect 8390 19751 8446 19760
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19310 8340 19654
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18290 8248 19110
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7576 12294 7696 12322
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7576 10010 7604 12294
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 10606 7696 12174
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7392 9982 7604 10010
rect 7392 8090 7420 9982
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9518 7604 9862
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 8634 7512 9386
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7208 7942 7328 7970
rect 7576 7954 7604 9454
rect 7564 7948 7616 7954
rect 7208 7886 7236 7942
rect 7564 7890 7616 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7286 7848 7342 7857
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6972 7160 7052 7188
rect 6920 7142 6972 7148
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 4842 6776 6802
rect 6840 5370 6868 6870
rect 7024 6254 7052 7160
rect 7116 6254 7144 7754
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6840 5001 6868 5306
rect 6826 4992 6882 5001
rect 6826 4927 6882 4936
rect 6748 4814 6868 4842
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6196 4542 6500 4570
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6380 2446 6408 3946
rect 6472 3398 6500 4542
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 2514 6500 3334
rect 6656 2666 6684 4626
rect 6840 4146 6868 4814
rect 6932 4690 6960 6122
rect 7024 4758 7052 6190
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 3534 6868 4082
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 2990 6868 3470
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6656 2638 6868 2666
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6380 1714 6408 2382
rect 6380 1686 6500 1714
rect 6472 800 6500 1686
rect 6840 800 6868 2638
rect 6932 2496 6960 4626
rect 7012 2508 7064 2514
rect 6932 2468 7012 2496
rect 7012 2450 7064 2456
rect 7208 800 7236 7822
rect 7286 7783 7342 7792
rect 7300 3670 7328 7783
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5778 7512 6054
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7668 4842 7696 10542
rect 7760 9518 7788 13806
rect 7852 13326 7880 15506
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7944 14278 7972 14418
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 13938 7972 14214
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12186 7880 13126
rect 7944 12306 7972 13874
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7852 12170 7972 12186
rect 7852 12164 7984 12170
rect 7852 12158 7932 12164
rect 7852 11694 7880 12158
rect 7932 12106 7984 12112
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7576 4814 7696 4842
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7300 3194 7328 3606
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7576 800 7604 4814
rect 7760 4026 7788 9454
rect 7852 9382 7880 11018
rect 7944 10538 7972 11494
rect 8036 10690 8064 17002
rect 8220 16250 8248 17682
rect 8312 16998 8340 18362
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15162 8248 15438
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 14482 8248 15098
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 11150 8156 13262
rect 8220 12481 8248 13738
rect 8206 12472 8262 12481
rect 8206 12407 8262 12416
rect 8206 12336 8262 12345
rect 8206 12271 8262 12280
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8036 10662 8156 10690
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7944 10062 7972 10474
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8036 9926 8064 10542
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 8128 9110 8156 10662
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7944 6390 7972 6734
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4146 7880 4422
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7760 3998 7880 4026
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7852 2938 7880 3998
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7944 3058 7972 3538
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7760 2650 7788 2926
rect 7852 2910 7972 2938
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7944 800 7972 2910
rect 8036 2854 8064 8978
rect 8220 3738 8248 12271
rect 8312 9194 8340 16458
rect 8404 16454 8432 19751
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8404 13326 8432 15506
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 11234 8432 13126
rect 8496 12850 8524 20896
rect 8588 18426 8616 24346
rect 8680 24274 8708 25774
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8588 16590 8616 18158
rect 8680 17610 8708 23598
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 15094 8616 16390
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8588 14550 8616 14894
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8680 14396 8708 17138
rect 8588 14368 8708 14396
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12306 8524 12582
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11762 8524 12106
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8404 11218 8524 11234
rect 8404 11212 8536 11218
rect 8404 11206 8484 11212
rect 8484 11154 8536 11160
rect 8312 9166 8432 9194
rect 8300 9104 8352 9110
rect 8298 9072 8300 9081
rect 8352 9072 8354 9081
rect 8298 9007 8354 9016
rect 8404 8430 8432 9166
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8312 7410 8340 7754
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8404 6780 8432 8366
rect 8312 6752 8432 6780
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2514 8064 2790
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8312 800 8340 6752
rect 8496 4690 8524 11154
rect 8588 9602 8616 14368
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12306 8708 13126
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8588 9574 8708 9602
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 8430 8616 9454
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8496 3194 8524 4626
rect 8680 4078 8708 9574
rect 8772 5302 8800 29038
rect 8886 28860 9182 28880
rect 8942 28858 8966 28860
rect 9022 28858 9046 28860
rect 9102 28858 9126 28860
rect 8964 28806 8966 28858
rect 9028 28806 9040 28858
rect 9102 28806 9104 28858
rect 8942 28804 8966 28806
rect 9022 28804 9046 28806
rect 9102 28804 9126 28806
rect 8886 28784 9182 28804
rect 8886 27772 9182 27792
rect 8942 27770 8966 27772
rect 9022 27770 9046 27772
rect 9102 27770 9126 27772
rect 8964 27718 8966 27770
rect 9028 27718 9040 27770
rect 9102 27718 9104 27770
rect 8942 27716 8966 27718
rect 9022 27716 9046 27718
rect 9102 27716 9126 27718
rect 8886 27696 9182 27716
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 8864 26926 8892 27066
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 8956 26858 8984 27406
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 8944 26852 8996 26858
rect 8944 26794 8996 26800
rect 8886 26684 9182 26704
rect 8942 26682 8966 26684
rect 9022 26682 9046 26684
rect 9102 26682 9126 26684
rect 8964 26630 8966 26682
rect 9028 26630 9040 26682
rect 9102 26630 9104 26682
rect 8942 26628 8966 26630
rect 9022 26628 9046 26630
rect 9102 26628 9126 26630
rect 8886 26608 9182 26628
rect 9232 26586 9260 26862
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 8886 25596 9182 25616
rect 8942 25594 8966 25596
rect 9022 25594 9046 25596
rect 9102 25594 9126 25596
rect 8964 25542 8966 25594
rect 9028 25542 9040 25594
rect 9102 25542 9104 25594
rect 8942 25540 8966 25542
rect 9022 25540 9046 25542
rect 9102 25540 9126 25542
rect 8886 25520 9182 25540
rect 9232 24857 9260 25638
rect 9218 24848 9274 24857
rect 9218 24783 9274 24792
rect 9220 24676 9272 24682
rect 9220 24618 9272 24624
rect 8886 24508 9182 24528
rect 8942 24506 8966 24508
rect 9022 24506 9046 24508
rect 9102 24506 9126 24508
rect 8964 24454 8966 24506
rect 9028 24454 9040 24506
rect 9102 24454 9104 24506
rect 8942 24452 8966 24454
rect 9022 24452 9046 24454
rect 9102 24452 9126 24454
rect 8886 24432 9182 24452
rect 9232 24410 9260 24618
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9220 23588 9272 23594
rect 9220 23530 9272 23536
rect 8886 23420 9182 23440
rect 8942 23418 8966 23420
rect 9022 23418 9046 23420
rect 9102 23418 9126 23420
rect 8964 23366 8966 23418
rect 9028 23366 9040 23418
rect 9102 23366 9104 23418
rect 8942 23364 8966 23366
rect 9022 23364 9046 23366
rect 9102 23364 9126 23366
rect 8886 23344 9182 23364
rect 8886 22332 9182 22352
rect 8942 22330 8966 22332
rect 9022 22330 9046 22332
rect 9102 22330 9126 22332
rect 8964 22278 8966 22330
rect 9028 22278 9040 22330
rect 9102 22278 9104 22330
rect 8942 22276 8966 22278
rect 9022 22276 9046 22278
rect 9102 22276 9126 22278
rect 8886 22256 9182 22276
rect 9232 21622 9260 23530
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9218 21448 9274 21457
rect 9218 21383 9274 21392
rect 8886 21244 9182 21264
rect 8942 21242 8966 21244
rect 9022 21242 9046 21244
rect 9102 21242 9126 21244
rect 8964 21190 8966 21242
rect 9028 21190 9040 21242
rect 9102 21190 9104 21242
rect 8942 21188 8966 21190
rect 9022 21188 9046 21190
rect 9102 21188 9126 21190
rect 8886 21168 9182 21188
rect 9126 21040 9182 21049
rect 9126 20975 9128 20984
rect 9180 20975 9182 20984
rect 9128 20946 9180 20952
rect 9140 20874 9168 20946
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 8850 20496 8906 20505
rect 8850 20431 8906 20440
rect 8864 20398 8892 20431
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8886 20156 9182 20176
rect 8942 20154 8966 20156
rect 9022 20154 9046 20156
rect 9102 20154 9126 20156
rect 8964 20102 8966 20154
rect 9028 20102 9040 20154
rect 9102 20102 9104 20154
rect 8942 20100 8966 20102
rect 9022 20100 9046 20102
rect 9102 20100 9126 20102
rect 8886 20080 9182 20100
rect 8886 19068 9182 19088
rect 8942 19066 8966 19068
rect 9022 19066 9046 19068
rect 9102 19066 9126 19068
rect 8964 19014 8966 19066
rect 9028 19014 9040 19066
rect 9102 19014 9104 19066
rect 8942 19012 8966 19014
rect 9022 19012 9046 19014
rect 9102 19012 9126 19014
rect 8886 18992 9182 19012
rect 8886 17980 9182 18000
rect 8942 17978 8966 17980
rect 9022 17978 9046 17980
rect 9102 17978 9126 17980
rect 8964 17926 8966 17978
rect 9028 17926 9040 17978
rect 9102 17926 9104 17978
rect 8942 17924 8966 17926
rect 9022 17924 9046 17926
rect 9102 17924 9126 17926
rect 8886 17904 9182 17924
rect 8886 16892 9182 16912
rect 8942 16890 8966 16892
rect 9022 16890 9046 16892
rect 9102 16890 9126 16892
rect 8964 16838 8966 16890
rect 9028 16838 9040 16890
rect 9102 16838 9104 16890
rect 8942 16836 8966 16838
rect 9022 16836 9046 16838
rect 9102 16836 9126 16838
rect 8886 16816 9182 16836
rect 8886 15804 9182 15824
rect 8942 15802 8966 15804
rect 9022 15802 9046 15804
rect 9102 15802 9126 15804
rect 8964 15750 8966 15802
rect 9028 15750 9040 15802
rect 9102 15750 9104 15802
rect 8942 15748 8966 15750
rect 9022 15748 9046 15750
rect 9102 15748 9126 15750
rect 8886 15728 9182 15748
rect 9232 15570 9260 21383
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8886 14716 9182 14736
rect 8942 14714 8966 14716
rect 9022 14714 9046 14716
rect 9102 14714 9126 14716
rect 8964 14662 8966 14714
rect 9028 14662 9040 14714
rect 9102 14662 9104 14714
rect 8942 14660 8966 14662
rect 9022 14660 9046 14662
rect 9102 14660 9126 14662
rect 8886 14640 9182 14660
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8864 13802 8892 14486
rect 9232 14006 9260 15302
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8886 13628 9182 13648
rect 8942 13626 8966 13628
rect 9022 13626 9046 13628
rect 9102 13626 9126 13628
rect 8964 13574 8966 13626
rect 9028 13574 9040 13626
rect 9102 13574 9104 13626
rect 8942 13572 8966 13574
rect 9022 13572 9046 13574
rect 9102 13572 9126 13574
rect 8886 13552 9182 13572
rect 9232 13512 9260 13942
rect 8956 13484 9260 13512
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12714 8892 12786
rect 8956 12782 8984 13484
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8886 12540 9182 12560
rect 8942 12538 8966 12540
rect 9022 12538 9046 12540
rect 9102 12538 9126 12540
rect 8964 12486 8966 12538
rect 9028 12486 9040 12538
rect 9102 12486 9104 12538
rect 8942 12484 8966 12486
rect 9022 12484 9046 12486
rect 9102 12484 9126 12486
rect 8886 12464 9182 12484
rect 8886 11452 9182 11472
rect 8942 11450 8966 11452
rect 9022 11450 9046 11452
rect 9102 11450 9126 11452
rect 8964 11398 8966 11450
rect 9028 11398 9040 11450
rect 9102 11398 9104 11450
rect 8942 11396 8966 11398
rect 9022 11396 9046 11398
rect 9102 11396 9126 11398
rect 8886 11376 9182 11396
rect 8886 10364 9182 10384
rect 8942 10362 8966 10364
rect 9022 10362 9046 10364
rect 9102 10362 9126 10364
rect 8964 10310 8966 10362
rect 9028 10310 9040 10362
rect 9102 10310 9104 10362
rect 8942 10308 8966 10310
rect 9022 10308 9046 10310
rect 9102 10308 9126 10310
rect 8886 10288 9182 10308
rect 8886 9276 9182 9296
rect 8942 9274 8966 9276
rect 9022 9274 9046 9276
rect 9102 9274 9126 9276
rect 8964 9222 8966 9274
rect 9028 9222 9040 9274
rect 9102 9222 9104 9274
rect 8942 9220 8966 9222
rect 9022 9220 9046 9222
rect 9102 9220 9126 9222
rect 8886 9200 9182 9220
rect 9232 9110 9260 13262
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 8886 8188 9182 8208
rect 8942 8186 8966 8188
rect 9022 8186 9046 8188
rect 9102 8186 9126 8188
rect 8964 8134 8966 8186
rect 9028 8134 9040 8186
rect 9102 8134 9104 8186
rect 8942 8132 8966 8134
rect 9022 8132 9046 8134
rect 9102 8132 9126 8134
rect 8886 8112 9182 8132
rect 9232 7954 9260 9046
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 8886 7100 9182 7120
rect 8942 7098 8966 7100
rect 9022 7098 9046 7100
rect 9102 7098 9126 7100
rect 8964 7046 8966 7098
rect 9028 7046 9040 7098
rect 9102 7046 9104 7098
rect 8942 7044 8966 7046
rect 9022 7044 9046 7046
rect 9102 7044 9126 7046
rect 8886 7024 9182 7044
rect 8886 6012 9182 6032
rect 8942 6010 8966 6012
rect 9022 6010 9046 6012
rect 9102 6010 9126 6012
rect 8964 5958 8966 6010
rect 9028 5958 9040 6010
rect 9102 5958 9104 6010
rect 8942 5956 8966 5958
rect 9022 5956 9046 5958
rect 9102 5956 9126 5958
rect 8886 5936 9182 5956
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8886 4924 9182 4944
rect 8942 4922 8966 4924
rect 9022 4922 9046 4924
rect 9102 4922 9126 4924
rect 8964 4870 8966 4922
rect 9028 4870 9040 4922
rect 9102 4870 9104 4922
rect 8942 4868 8966 4870
rect 9022 4868 9046 4870
rect 9102 4868 9126 4870
rect 8886 4848 9182 4868
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8680 800 8708 4014
rect 8886 3836 9182 3856
rect 8942 3834 8966 3836
rect 9022 3834 9046 3836
rect 9102 3834 9126 3836
rect 8964 3782 8966 3834
rect 9028 3782 9040 3834
rect 9102 3782 9104 3834
rect 8942 3780 8966 3782
rect 9022 3780 9046 3782
rect 9102 3780 9126 3782
rect 8886 3760 9182 3780
rect 9324 3380 9352 34478
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9416 30870 9444 31078
rect 9404 30864 9456 30870
rect 9404 30806 9456 30812
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9416 25838 9444 29650
rect 9508 26081 9536 31690
rect 9494 26072 9550 26081
rect 9494 26007 9496 26016
rect 9548 26007 9550 26016
rect 9496 25978 9548 25984
rect 9508 25947 9536 25978
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9496 25764 9548 25770
rect 9496 25706 9548 25712
rect 9508 24721 9536 25706
rect 9494 24712 9550 24721
rect 9494 24647 9550 24656
rect 9508 23662 9536 24647
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 13161 9444 22374
rect 9508 22080 9536 23190
rect 9600 22438 9628 34598
rect 9784 34542 9812 36518
rect 9864 34672 9916 34678
rect 9864 34614 9916 34620
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9876 34066 9904 34614
rect 9956 34536 10008 34542
rect 9956 34478 10008 34484
rect 9968 34202 9996 34478
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9864 34060 9916 34066
rect 9864 34002 9916 34008
rect 10060 33930 10088 37606
rect 10244 35170 10272 39850
rect 10612 38962 10640 43182
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 10600 38956 10652 38962
rect 10600 38898 10652 38904
rect 10600 38820 10652 38826
rect 10600 38762 10652 38768
rect 10416 37392 10468 37398
rect 10468 37340 10548 37346
rect 10416 37334 10548 37340
rect 10324 37324 10376 37330
rect 10428 37318 10548 37334
rect 10324 37266 10376 37272
rect 10336 36718 10364 37266
rect 10324 36712 10376 36718
rect 10324 36654 10376 36660
rect 10336 36582 10364 36654
rect 10324 36576 10376 36582
rect 10324 36518 10376 36524
rect 10244 35142 10364 35170
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10244 34746 10272 35022
rect 10232 34740 10284 34746
rect 10232 34682 10284 34688
rect 10140 34468 10192 34474
rect 10140 34410 10192 34416
rect 10048 33924 10100 33930
rect 10048 33866 10100 33872
rect 10048 33448 10100 33454
rect 10048 33390 10100 33396
rect 9680 33312 9732 33318
rect 9680 33254 9732 33260
rect 9692 32434 9720 33254
rect 9772 32972 9824 32978
rect 9772 32914 9824 32920
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9692 29238 9720 31418
rect 9784 31346 9812 32914
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9772 31340 9824 31346
rect 9772 31282 9824 31288
rect 9876 29782 9904 32710
rect 9968 32434 9996 32846
rect 9956 32428 10008 32434
rect 9956 32370 10008 32376
rect 10060 32026 10088 33390
rect 10152 32366 10180 34410
rect 10232 33448 10284 33454
rect 10232 33390 10284 33396
rect 10244 32978 10272 33390
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10336 32552 10364 35142
rect 10416 34060 10468 34066
rect 10416 34002 10468 34008
rect 10244 32524 10364 32552
rect 10140 32360 10192 32366
rect 10140 32302 10192 32308
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 10060 31872 10088 31962
rect 9968 31844 10088 31872
rect 9968 30802 9996 31844
rect 10244 31804 10272 32524
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10336 31822 10364 32370
rect 10428 32366 10456 34002
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10060 31776 10272 31804
rect 10324 31816 10376 31822
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9956 30660 10008 30666
rect 9956 30602 10008 30608
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9692 28150 9720 29174
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9784 27538 9812 29446
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9692 27130 9720 27474
rect 9876 27470 9904 27950
rect 9864 27464 9916 27470
rect 9864 27406 9916 27412
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9692 26897 9720 26930
rect 9772 26920 9824 26926
rect 9678 26888 9734 26897
rect 9772 26862 9824 26868
rect 9678 26823 9734 26832
rect 9784 26586 9812 26862
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9692 24342 9720 25298
rect 9680 24336 9732 24342
rect 9680 24278 9732 24284
rect 9784 24177 9812 26386
rect 9876 26246 9904 27406
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9770 24168 9826 24177
rect 9770 24103 9826 24112
rect 9680 24064 9732 24070
rect 9678 24032 9680 24041
rect 9732 24032 9734 24041
rect 9678 23967 9734 23976
rect 9678 23760 9734 23769
rect 9678 23695 9734 23704
rect 9692 22506 9720 23695
rect 9876 23254 9904 24822
rect 9968 24614 9996 30602
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9680 22500 9732 22506
rect 9680 22442 9732 22448
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9680 22092 9732 22098
rect 9508 22052 9628 22080
rect 9494 21992 9550 22001
rect 9494 21927 9550 21936
rect 9402 13152 9458 13161
rect 9402 13087 9458 13096
rect 9508 9704 9536 21927
rect 9600 21593 9628 22052
rect 9680 22034 9732 22040
rect 9586 21584 9642 21593
rect 9586 21519 9642 21528
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9600 20602 9628 21422
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9600 19990 9628 20334
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 18986 9628 19722
rect 9692 19174 9720 22034
rect 9784 21962 9812 22374
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 20924 9812 21422
rect 9876 21078 9904 21966
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9784 20896 9904 20924
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9600 18958 9720 18986
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 16658 9628 18702
rect 9692 18630 9720 18958
rect 9784 18884 9812 19858
rect 9876 19786 9904 20896
rect 9968 20398 9996 22918
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 10060 19292 10088 31776
rect 10324 31758 10376 31764
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10152 29102 10180 29582
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10152 24698 10180 29038
rect 10244 27538 10272 31622
rect 10428 31482 10456 32302
rect 10416 31476 10468 31482
rect 10416 31418 10468 31424
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10336 30938 10364 31282
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10428 30938 10456 31214
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10416 30932 10468 30938
rect 10416 30874 10468 30880
rect 10324 30796 10376 30802
rect 10324 30738 10376 30744
rect 10336 29102 10364 30738
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10416 27940 10468 27946
rect 10416 27882 10468 27888
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10428 26518 10456 27882
rect 10416 26512 10468 26518
rect 10416 26454 10468 26460
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10428 24818 10456 26182
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10152 24670 10364 24698
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10138 24440 10194 24449
rect 10138 24375 10194 24384
rect 10152 24342 10180 24375
rect 10140 24336 10192 24342
rect 10140 24278 10192 24284
rect 10138 24168 10194 24177
rect 10138 24103 10194 24112
rect 10152 24070 10180 24103
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10152 22710 10180 23122
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22098 10180 22374
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10060 19264 10180 19292
rect 10048 19168 10100 19174
rect 9954 19136 10010 19145
rect 10048 19110 10100 19116
rect 9954 19071 10010 19080
rect 9784 18856 9904 18884
rect 9876 18748 9904 18856
rect 9784 18720 9904 18748
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9784 16402 9812 18720
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9692 16374 9812 16402
rect 9692 14890 9720 16374
rect 9876 16114 9904 17002
rect 9968 16794 9996 19071
rect 10060 18850 10088 19110
rect 10152 18970 10180 19264
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10060 18822 10180 18850
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 16590 10088 18634
rect 10152 18426 10180 18822
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10152 16697 10180 17070
rect 10138 16688 10194 16697
rect 10138 16623 10140 16632
rect 10192 16623 10194 16632
rect 10140 16594 10192 16600
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9784 15570 9812 15982
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 10060 14958 10088 16526
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9784 13870 9812 14894
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 14074 9996 14214
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13394 9628 13738
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11830 9628 12038
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9692 11132 9720 13262
rect 9876 12918 9904 13262
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 10060 12850 10088 14894
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9772 11144 9824 11150
rect 9692 11104 9772 11132
rect 9692 10130 9720 11104
rect 9772 11086 9824 11092
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9508 9676 9628 9704
rect 9600 9568 9628 9676
rect 9508 9540 9628 9568
rect 9508 7546 9536 9540
rect 9692 9518 9720 10066
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 8838 9720 9454
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7954 9628 8230
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9692 7886 9720 8774
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 7562 9720 7822
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9600 7534 9720 7562
rect 9600 5914 9628 7534
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5710 9628 5850
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9232 3352 9352 3380
rect 8886 2748 9182 2768
rect 8942 2746 8966 2748
rect 9022 2746 9046 2748
rect 9102 2746 9126 2748
rect 8964 2694 8966 2746
rect 9028 2694 9040 2746
rect 9102 2694 9104 2746
rect 8942 2692 8966 2694
rect 9022 2692 9046 2694
rect 9102 2692 9126 2694
rect 8886 2672 9182 2692
rect 9232 2632 9260 3352
rect 9310 3224 9366 3233
rect 9310 3159 9366 3168
rect 8956 2604 9260 2632
rect 8956 800 8984 2604
rect 9324 800 9352 3159
rect 9692 800 9720 7414
rect 9784 4826 9812 8298
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6254 9904 6802
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 6458 9996 6734
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9968 5778 9996 6122
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9784 4010 9812 4762
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 2514 9812 3538
rect 9876 2990 9904 4082
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3602 9996 3878
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10060 800 10088 7482
rect 10152 6322 10180 9862
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 2514 10180 5034
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10244 1442 10272 24550
rect 10336 17134 10364 24670
rect 10428 22506 10456 24754
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10428 21078 10456 21354
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 19310 10456 19654
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10428 16658 10456 18838
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 14958 10456 16594
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10428 12714 10456 14894
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 9518 10456 11698
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 8401 10456 9454
rect 10414 8392 10470 8401
rect 10414 8327 10470 8336
rect 10520 7478 10548 37318
rect 10612 35306 10640 38762
rect 10704 36378 10732 42094
rect 11060 41064 11112 41070
rect 11060 41006 11112 41012
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 10876 39500 10928 39506
rect 10876 39442 10928 39448
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 10796 36922 10824 39374
rect 10888 38418 10916 39442
rect 10876 38412 10928 38418
rect 10876 38354 10928 38360
rect 10980 38298 11008 39918
rect 10888 38270 11008 38298
rect 10888 37874 10916 38270
rect 10968 38208 11020 38214
rect 10968 38150 11020 38156
rect 10980 38010 11008 38150
rect 10968 38004 11020 38010
rect 10968 37946 11020 37952
rect 10876 37868 10928 37874
rect 10876 37810 10928 37816
rect 10784 36916 10836 36922
rect 10784 36858 10836 36864
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10980 35630 11008 36858
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10612 35278 10824 35306
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 10612 33454 10640 33934
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10612 33114 10640 33390
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10692 32972 10744 32978
rect 10692 32914 10744 32920
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10612 31278 10640 32166
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 10704 26874 10732 32914
rect 10796 27033 10824 35278
rect 11072 34202 11100 41006
rect 11164 41002 11192 46446
rect 11256 45558 11284 47194
rect 11440 47002 11468 49200
rect 12176 47258 12204 49200
rect 13004 47410 13032 49200
rect 13004 47382 13492 47410
rect 12164 47252 12216 47258
rect 12164 47194 12216 47200
rect 12532 47116 12584 47122
rect 12532 47058 12584 47064
rect 12440 47048 12492 47054
rect 11440 46974 11652 47002
rect 12440 46990 12492 46996
rect 11428 46912 11480 46918
rect 11428 46854 11480 46860
rect 11336 46368 11388 46374
rect 11336 46310 11388 46316
rect 11244 45552 11296 45558
rect 11244 45494 11296 45500
rect 11348 44946 11376 46310
rect 11336 44940 11388 44946
rect 11336 44882 11388 44888
rect 11348 44470 11376 44882
rect 11336 44464 11388 44470
rect 11336 44406 11388 44412
rect 11348 43790 11376 44406
rect 11440 44266 11468 46854
rect 11520 44940 11572 44946
rect 11520 44882 11572 44888
rect 11428 44260 11480 44266
rect 11428 44202 11480 44208
rect 11428 43852 11480 43858
rect 11428 43794 11480 43800
rect 11336 43784 11388 43790
rect 11336 43726 11388 43732
rect 11348 43450 11376 43726
rect 11336 43444 11388 43450
rect 11336 43386 11388 43392
rect 11336 42152 11388 42158
rect 11336 42094 11388 42100
rect 11348 41750 11376 42094
rect 11336 41744 11388 41750
rect 11336 41686 11388 41692
rect 11348 41070 11376 41686
rect 11336 41064 11388 41070
rect 11336 41006 11388 41012
rect 11152 40996 11204 41002
rect 11152 40938 11204 40944
rect 11152 40588 11204 40594
rect 11152 40530 11204 40536
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 10980 32026 11008 32846
rect 10968 32020 11020 32026
rect 10968 31962 11020 31968
rect 11072 31872 11100 33866
rect 10980 31844 11100 31872
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 10888 27606 10916 27950
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10782 27024 10838 27033
rect 10782 26959 10838 26968
rect 10980 26874 11008 31844
rect 11060 31748 11112 31754
rect 11060 31690 11112 31696
rect 11072 30666 11100 31690
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 11164 30326 11192 40530
rect 11440 40118 11468 43794
rect 11532 42226 11560 44882
rect 11624 43314 11652 46974
rect 12348 46912 12400 46918
rect 12348 46854 12400 46860
rect 12360 46102 12388 46854
rect 12348 46096 12400 46102
rect 12348 46038 12400 46044
rect 12452 45082 12480 46990
rect 12544 46442 12572 47058
rect 12852 46812 13148 46832
rect 12908 46810 12932 46812
rect 12988 46810 13012 46812
rect 13068 46810 13092 46812
rect 12930 46758 12932 46810
rect 12994 46758 13006 46810
rect 13068 46758 13070 46810
rect 12908 46756 12932 46758
rect 12988 46756 13012 46758
rect 13068 46756 13092 46758
rect 12852 46736 13148 46756
rect 12532 46436 12584 46442
rect 12532 46378 12584 46384
rect 13176 46436 13228 46442
rect 13176 46378 13228 46384
rect 12716 46368 12768 46374
rect 12716 46310 12768 46316
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 12440 45076 12492 45082
rect 12440 45018 12492 45024
rect 12544 45014 12572 45358
rect 12728 45014 12756 46310
rect 12852 45724 13148 45744
rect 12908 45722 12932 45724
rect 12988 45722 13012 45724
rect 13068 45722 13092 45724
rect 12930 45670 12932 45722
rect 12994 45670 13006 45722
rect 13068 45670 13070 45722
rect 12908 45668 12932 45670
rect 12988 45668 13012 45670
rect 13068 45668 13092 45670
rect 12852 45648 13148 45668
rect 12532 45008 12584 45014
rect 12532 44950 12584 44956
rect 12716 45008 12768 45014
rect 12716 44950 12768 44956
rect 12624 44940 12676 44946
rect 12624 44882 12676 44888
rect 12440 44260 12492 44266
rect 12440 44202 12492 44208
rect 12256 43784 12308 43790
rect 12256 43726 12308 43732
rect 12268 43314 12296 43726
rect 12452 43722 12480 44202
rect 12532 43784 12584 43790
rect 12532 43726 12584 43732
rect 12440 43716 12492 43722
rect 12440 43658 12492 43664
rect 11612 43308 11664 43314
rect 11612 43250 11664 43256
rect 12256 43308 12308 43314
rect 12256 43250 12308 43256
rect 11624 42702 11652 43250
rect 12440 43104 12492 43110
rect 12440 43046 12492 43052
rect 12452 42770 12480 43046
rect 12440 42764 12492 42770
rect 12440 42706 12492 42712
rect 11612 42696 11664 42702
rect 11612 42638 11664 42644
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 11520 42220 11572 42226
rect 11520 42162 11572 42168
rect 11796 41676 11848 41682
rect 11796 41618 11848 41624
rect 11520 41064 11572 41070
rect 11520 41006 11572 41012
rect 11532 40594 11560 41006
rect 11520 40588 11572 40594
rect 11520 40530 11572 40536
rect 11428 40112 11480 40118
rect 11428 40054 11480 40060
rect 11428 39976 11480 39982
rect 11532 39964 11560 40530
rect 11480 39936 11560 39964
rect 11612 39976 11664 39982
rect 11428 39918 11480 39924
rect 11612 39918 11664 39924
rect 11336 38888 11388 38894
rect 11334 38856 11336 38865
rect 11388 38856 11390 38865
rect 11334 38791 11390 38800
rect 11336 38412 11388 38418
rect 11336 38354 11388 38360
rect 11244 38344 11296 38350
rect 11244 38286 11296 38292
rect 11256 37398 11284 38286
rect 11348 37806 11376 38354
rect 11440 38010 11468 39918
rect 11624 39098 11652 39918
rect 11612 39092 11664 39098
rect 11612 39034 11664 39040
rect 11428 38004 11480 38010
rect 11428 37946 11480 37952
rect 11336 37800 11388 37806
rect 11336 37742 11388 37748
rect 11612 37732 11664 37738
rect 11612 37674 11664 37680
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11244 37392 11296 37398
rect 11244 37334 11296 37340
rect 11532 37330 11560 37606
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 11256 36310 11284 37198
rect 11336 36712 11388 36718
rect 11336 36654 11388 36660
rect 11244 36304 11296 36310
rect 11244 36246 11296 36252
rect 11256 34066 11284 36246
rect 11348 36106 11376 36654
rect 11624 36582 11652 37674
rect 11704 37392 11756 37398
rect 11704 37334 11756 37340
rect 11612 36576 11664 36582
rect 11612 36518 11664 36524
rect 11716 36394 11744 37334
rect 11532 36366 11744 36394
rect 11532 36310 11560 36366
rect 11520 36304 11572 36310
rect 11520 36246 11572 36252
rect 11428 36236 11480 36242
rect 11428 36178 11480 36184
rect 11336 36100 11388 36106
rect 11336 36042 11388 36048
rect 11348 35714 11376 36042
rect 11440 35834 11468 36178
rect 11428 35828 11480 35834
rect 11428 35770 11480 35776
rect 11348 35686 11468 35714
rect 11440 35494 11468 35686
rect 11428 35488 11480 35494
rect 11428 35430 11480 35436
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 11348 34542 11376 34886
rect 11440 34746 11468 35430
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 11532 34626 11560 36246
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11612 35556 11664 35562
rect 11612 35498 11664 35504
rect 11440 34598 11560 34626
rect 11336 34536 11388 34542
rect 11336 34478 11388 34484
rect 11440 34134 11468 34598
rect 11428 34128 11480 34134
rect 11428 34070 11480 34076
rect 11244 34060 11296 34066
rect 11244 34002 11296 34008
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 11348 31890 11376 32914
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11440 30938 11468 34070
rect 11520 33584 11572 33590
rect 11520 33526 11572 33532
rect 11428 30932 11480 30938
rect 11428 30874 11480 30880
rect 11152 30320 11204 30326
rect 11152 30262 11204 30268
rect 11440 30190 11468 30874
rect 11532 30666 11560 33526
rect 11520 30660 11572 30666
rect 11520 30602 11572 30608
rect 11428 30184 11480 30190
rect 11428 30126 11480 30132
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29102 11100 29990
rect 11060 29096 11112 29102
rect 11060 29038 11112 29044
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 10704 26846 10824 26874
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10612 26042 10640 26250
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10692 25764 10744 25770
rect 10692 25706 10744 25712
rect 10704 24818 10732 25706
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10690 24304 10746 24313
rect 10690 24239 10692 24248
rect 10744 24239 10746 24248
rect 10692 24210 10744 24216
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10612 21010 10640 24006
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10704 22574 10732 23802
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10796 19394 10824 26846
rect 10888 26846 11008 26874
rect 10888 24750 10916 26846
rect 11072 25838 11100 27270
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 11072 24206 11100 25094
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11164 23730 11192 25842
rect 11256 25362 11284 28970
rect 11336 28960 11388 28966
rect 11336 28902 11388 28908
rect 11348 28626 11376 28902
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11256 24274 11284 25298
rect 11348 24750 11376 27474
rect 11440 27130 11468 30126
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11532 26466 11560 29786
rect 11624 27470 11652 35498
rect 11716 35290 11744 35770
rect 11704 35284 11756 35290
rect 11704 35226 11756 35232
rect 11704 32224 11756 32230
rect 11704 32166 11756 32172
rect 11716 31890 11744 32166
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11716 29714 11744 31826
rect 11808 30870 11836 41618
rect 12452 40594 12480 42502
rect 12544 41614 12572 43726
rect 12532 41608 12584 41614
rect 12532 41550 12584 41556
rect 12636 41138 12664 44882
rect 12716 44736 12768 44742
rect 12716 44678 12768 44684
rect 12728 43654 12756 44678
rect 12852 44636 13148 44656
rect 12908 44634 12932 44636
rect 12988 44634 13012 44636
rect 13068 44634 13092 44636
rect 12930 44582 12932 44634
rect 12994 44582 13006 44634
rect 13068 44582 13070 44634
rect 12908 44580 12932 44582
rect 12988 44580 13012 44582
rect 13068 44580 13092 44582
rect 12852 44560 13148 44580
rect 13188 44266 13216 46378
rect 13360 45484 13412 45490
rect 13360 45426 13412 45432
rect 13176 44260 13228 44266
rect 13176 44202 13228 44208
rect 12808 44192 12860 44198
rect 12808 44134 12860 44140
rect 12820 43926 12848 44134
rect 12808 43920 12860 43926
rect 12808 43862 12860 43868
rect 12716 43648 12768 43654
rect 12716 43590 12768 43596
rect 12728 41274 12756 43590
rect 12852 43548 13148 43568
rect 12908 43546 12932 43548
rect 12988 43546 13012 43548
rect 13068 43546 13092 43548
rect 12930 43494 12932 43546
rect 12994 43494 13006 43546
rect 13068 43494 13070 43546
rect 12908 43492 12932 43494
rect 12988 43492 13012 43494
rect 13068 43492 13092 43494
rect 12852 43472 13148 43492
rect 13372 43246 13400 45426
rect 13464 44010 13492 47382
rect 13740 46918 13768 49200
rect 14568 47190 14596 49200
rect 13820 47184 13872 47190
rect 13820 47126 13872 47132
rect 14556 47184 14608 47190
rect 14556 47126 14608 47132
rect 13728 46912 13780 46918
rect 13728 46854 13780 46860
rect 13636 45824 13688 45830
rect 13636 45766 13688 45772
rect 13648 44742 13676 45766
rect 13832 45626 13860 47126
rect 14004 47116 14056 47122
rect 14004 47058 14056 47064
rect 14188 47116 14240 47122
rect 14188 47058 14240 47064
rect 13912 46028 13964 46034
rect 13912 45970 13964 45976
rect 13820 45620 13872 45626
rect 13820 45562 13872 45568
rect 13636 44736 13688 44742
rect 13636 44678 13688 44684
rect 13924 44418 13952 45970
rect 13832 44390 13952 44418
rect 13464 43994 13584 44010
rect 13464 43988 13596 43994
rect 13464 43982 13544 43988
rect 12808 43240 12860 43246
rect 12808 43182 12860 43188
rect 13360 43240 13412 43246
rect 13360 43182 13412 43188
rect 12820 42702 12848 43182
rect 13464 42906 13492 43982
rect 13544 43930 13596 43936
rect 13544 43852 13596 43858
rect 13544 43794 13596 43800
rect 13452 42900 13504 42906
rect 13452 42842 13504 42848
rect 12808 42696 12860 42702
rect 12808 42638 12860 42644
rect 12852 42460 13148 42480
rect 12908 42458 12932 42460
rect 12988 42458 13012 42460
rect 13068 42458 13092 42460
rect 12930 42406 12932 42458
rect 12994 42406 13006 42458
rect 13068 42406 13070 42458
rect 12908 42404 12932 42406
rect 12988 42404 13012 42406
rect 13068 42404 13092 42406
rect 12852 42384 13148 42404
rect 13556 42226 13584 43794
rect 13544 42220 13596 42226
rect 13544 42162 13596 42168
rect 13176 41676 13228 41682
rect 13176 41618 13228 41624
rect 12852 41372 13148 41392
rect 12908 41370 12932 41372
rect 12988 41370 13012 41372
rect 13068 41370 13092 41372
rect 12930 41318 12932 41370
rect 12994 41318 13006 41370
rect 13068 41318 13070 41370
rect 12908 41316 12932 41318
rect 12988 41316 13012 41318
rect 13068 41316 13092 41318
rect 12852 41296 13148 41316
rect 12716 41268 12768 41274
rect 12716 41210 12768 41216
rect 12624 41132 12676 41138
rect 12624 41074 12676 41080
rect 12440 40588 12492 40594
rect 12440 40530 12492 40536
rect 12452 39506 12480 40530
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12728 40186 12756 40462
rect 12852 40284 13148 40304
rect 12908 40282 12932 40284
rect 12988 40282 13012 40284
rect 13068 40282 13092 40284
rect 12930 40230 12932 40282
rect 12994 40230 13006 40282
rect 13068 40230 13070 40282
rect 12908 40228 12932 40230
rect 12988 40228 13012 40230
rect 13068 40228 13092 40230
rect 12852 40208 13148 40228
rect 12716 40180 12768 40186
rect 12716 40122 12768 40128
rect 13188 39506 13216 41618
rect 13268 41064 13320 41070
rect 13268 41006 13320 41012
rect 12440 39500 12492 39506
rect 12440 39442 12492 39448
rect 13176 39500 13228 39506
rect 13176 39442 13228 39448
rect 12624 39364 12676 39370
rect 12624 39306 12676 39312
rect 12072 39024 12124 39030
rect 12070 38992 12072 39001
rect 12124 38992 12126 39001
rect 12636 38962 12664 39306
rect 12852 39196 13148 39216
rect 12908 39194 12932 39196
rect 12988 39194 13012 39196
rect 13068 39194 13092 39196
rect 12930 39142 12932 39194
rect 12994 39142 13006 39194
rect 13068 39142 13070 39194
rect 12908 39140 12932 39142
rect 12988 39140 13012 39142
rect 13068 39140 13092 39142
rect 12852 39120 13148 39140
rect 12070 38927 12126 38936
rect 12624 38956 12676 38962
rect 12624 38898 12676 38904
rect 12716 38888 12768 38894
rect 12716 38830 12768 38836
rect 12728 38010 12756 38830
rect 13188 38214 13216 39442
rect 13176 38208 13228 38214
rect 13176 38150 13228 38156
rect 12852 38108 13148 38128
rect 12908 38106 12932 38108
rect 12988 38106 13012 38108
rect 13068 38106 13092 38108
rect 12930 38054 12932 38106
rect 12994 38054 13006 38106
rect 13068 38054 13070 38106
rect 12908 38052 12932 38054
rect 12988 38052 13012 38054
rect 13068 38052 13092 38054
rect 12852 38032 13148 38052
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12256 37936 12308 37942
rect 12256 37878 12308 37884
rect 12072 37868 12124 37874
rect 12072 37810 12124 37816
rect 12084 37466 12112 37810
rect 12072 37460 12124 37466
rect 12072 37402 12124 37408
rect 11888 35624 11940 35630
rect 11888 35566 11940 35572
rect 11900 35018 11928 35566
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 11888 35012 11940 35018
rect 11888 34954 11940 34960
rect 11992 34950 12020 35226
rect 11980 34944 12032 34950
rect 11980 34886 12032 34892
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11796 30864 11848 30870
rect 11796 30806 11848 30812
rect 11796 30320 11848 30326
rect 11796 30262 11848 30268
rect 11704 29708 11756 29714
rect 11704 29650 11756 29656
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 11532 26438 11652 26466
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11428 25832 11480 25838
rect 11428 25774 11480 25780
rect 11440 25362 11468 25774
rect 11532 25498 11560 26318
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11428 25356 11480 25362
rect 11480 25316 11560 25344
rect 11428 25298 11480 25304
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 10888 19446 10916 23666
rect 11256 23361 11284 24074
rect 11242 23352 11298 23361
rect 11242 23287 11298 23296
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 21486 11008 22510
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11164 22098 11192 22374
rect 11244 22160 11296 22166
rect 11348 22137 11376 24686
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 24449 11468 24550
rect 11426 24440 11482 24449
rect 11426 24375 11482 24384
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11440 23186 11468 24210
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11440 23089 11468 23122
rect 11426 23080 11482 23089
rect 11426 23015 11482 23024
rect 11244 22102 11296 22108
rect 11334 22128 11390 22137
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11152 21616 11204 21622
rect 11150 21584 11152 21593
rect 11204 21584 11206 21593
rect 11150 21519 11206 21528
rect 10968 21480 11020 21486
rect 11152 21480 11204 21486
rect 10968 21422 11020 21428
rect 11150 21448 11152 21457
rect 11204 21448 11206 21457
rect 11150 21383 11206 21392
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11164 20398 11192 21286
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 19446 11008 20266
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10612 19366 10824 19394
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10612 17218 10640 19366
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10704 17338 10732 19178
rect 10888 18970 10916 19178
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10796 18306 10824 18770
rect 10796 18278 10916 18306
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10796 17542 10824 18158
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10612 17190 10732 17218
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 5166 10364 6734
rect 10428 5574 10456 6870
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10428 4146 10456 5510
rect 10612 4842 10640 17070
rect 10704 7546 10732 17190
rect 10888 15042 10916 18278
rect 10980 16454 11008 19246
rect 11072 16726 11100 19858
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18358 11192 19178
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 11256 18290 11284 22102
rect 11334 22063 11390 22072
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11348 21690 11376 21830
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 20534 11376 20742
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10888 15014 11008 15042
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10796 11626 10824 12718
rect 10888 12186 10916 14894
rect 10980 12374 11008 15014
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10888 12158 11008 12186
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11898 10916 12038
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 10606 10824 11562
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 9722 10824 10542
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10782 9208 10838 9217
rect 10782 9143 10838 9152
rect 10796 8906 10824 9143
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10888 8294 10916 11834
rect 10980 11762 11008 12158
rect 11072 11898 11100 12242
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11164 11762 11192 16594
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11256 14074 11284 14418
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11348 13870 11376 20334
rect 11440 19922 11468 21966
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11440 17610 11468 19858
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14618 11468 14758
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 13870 11468 14418
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11348 12782 11376 13806
rect 11532 13716 11560 25316
rect 11624 23730 11652 26438
rect 11808 25514 11836 30262
rect 11716 25486 11836 25514
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11624 22574 11652 23666
rect 11716 22778 11744 25486
rect 11900 24886 11928 33934
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 12084 30734 12112 31826
rect 12176 30870 12204 33866
rect 12164 30864 12216 30870
rect 12164 30806 12216 30812
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12176 30546 12204 30806
rect 12084 30518 12204 30546
rect 12084 30122 12112 30518
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 12072 30116 12124 30122
rect 12072 30058 12124 30064
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11992 26450 12020 27066
rect 12084 27062 12112 30058
rect 12176 29714 12204 30126
rect 12164 29708 12216 29714
rect 12164 29650 12216 29656
rect 12176 29306 12204 29650
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 12268 26874 12296 37878
rect 13176 37664 13228 37670
rect 13176 37606 13228 37612
rect 13188 37330 13216 37606
rect 13176 37324 13228 37330
rect 13176 37266 13228 37272
rect 12852 37020 13148 37040
rect 12908 37018 12932 37020
rect 12988 37018 13012 37020
rect 13068 37018 13092 37020
rect 12930 36966 12932 37018
rect 12994 36966 13006 37018
rect 13068 36966 13070 37018
rect 12908 36964 12932 36966
rect 12988 36964 13012 36966
rect 13068 36964 13092 36966
rect 12852 36944 13148 36964
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 12452 34202 12480 36722
rect 12716 36032 12768 36038
rect 12716 35974 12768 35980
rect 12728 35698 12756 35974
rect 12852 35932 13148 35952
rect 12908 35930 12932 35932
rect 12988 35930 13012 35932
rect 13068 35930 13092 35932
rect 12930 35878 12932 35930
rect 12994 35878 13006 35930
rect 13068 35878 13070 35930
rect 12908 35876 12932 35878
rect 12988 35876 13012 35878
rect 13068 35876 13092 35878
rect 12852 35856 13148 35876
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 12532 35148 12584 35154
rect 12820 35136 12848 35634
rect 12584 35108 12848 35136
rect 12532 35090 12584 35096
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12452 32978 12480 34002
rect 12544 33454 12572 34954
rect 12852 34844 13148 34864
rect 12908 34842 12932 34844
rect 12988 34842 13012 34844
rect 13068 34842 13092 34844
rect 12930 34790 12932 34842
rect 12994 34790 13006 34842
rect 13068 34790 13070 34842
rect 12908 34788 12932 34790
rect 12988 34788 13012 34790
rect 13068 34788 13092 34790
rect 12852 34768 13148 34788
rect 13188 34746 13216 37266
rect 13176 34740 13228 34746
rect 13176 34682 13228 34688
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12624 34536 12676 34542
rect 12624 34478 12676 34484
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 12440 32972 12492 32978
rect 12440 32914 12492 32920
rect 12544 32434 12572 33390
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 12532 31884 12584 31890
rect 12532 31826 12584 31832
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 12360 31346 12388 31622
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12452 29050 12480 31214
rect 12544 31210 12572 31826
rect 12532 31204 12584 31210
rect 12532 31146 12584 31152
rect 12636 30258 12664 34478
rect 12820 34066 12848 34546
rect 12808 34060 12860 34066
rect 12808 34002 12860 34008
rect 12852 33756 13148 33776
rect 12908 33754 12932 33756
rect 12988 33754 13012 33756
rect 13068 33754 13092 33756
rect 12930 33702 12932 33754
rect 12994 33702 13006 33754
rect 13068 33702 13070 33754
rect 12908 33700 12932 33702
rect 12988 33700 13012 33702
rect 13068 33700 13092 33702
rect 12852 33680 13148 33700
rect 12716 33448 12768 33454
rect 12716 33390 12768 33396
rect 12728 33114 12756 33390
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12852 32668 13148 32688
rect 12908 32666 12932 32668
rect 12988 32666 13012 32668
rect 13068 32666 13092 32668
rect 12930 32614 12932 32666
rect 12994 32614 13006 32666
rect 13068 32614 13070 32666
rect 12908 32612 12932 32614
rect 12988 32612 13012 32614
rect 13068 32612 13092 32614
rect 12852 32592 13148 32612
rect 12852 31580 13148 31600
rect 12908 31578 12932 31580
rect 12988 31578 13012 31580
rect 13068 31578 13092 31580
rect 12930 31526 12932 31578
rect 12994 31526 13006 31578
rect 13068 31526 13070 31578
rect 12908 31524 12932 31526
rect 12988 31524 13012 31526
rect 13068 31524 13092 31526
rect 12852 31504 13148 31524
rect 12852 30492 13148 30512
rect 12908 30490 12932 30492
rect 12988 30490 13012 30492
rect 13068 30490 13092 30492
rect 12930 30438 12932 30490
rect 12994 30438 13006 30490
rect 13068 30438 13070 30490
rect 12908 30436 12932 30438
rect 12988 30436 13012 30438
rect 13068 30436 13092 30438
rect 12852 30416 13148 30436
rect 12624 30252 12676 30258
rect 12624 30194 12676 30200
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 12624 29708 12676 29714
rect 12624 29650 12676 29656
rect 12532 29096 12584 29102
rect 12360 29044 12532 29050
rect 12360 29038 12584 29044
rect 12360 29022 12572 29038
rect 12360 28558 12388 29022
rect 12636 28626 12664 29650
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12728 29238 12756 29446
rect 12852 29404 13148 29424
rect 12908 29402 12932 29404
rect 12988 29402 13012 29404
rect 13068 29402 13092 29404
rect 12930 29350 12932 29402
rect 12994 29350 13006 29402
rect 13068 29350 13070 29402
rect 12908 29348 12932 29350
rect 12988 29348 13012 29350
rect 13068 29348 13092 29350
rect 12852 29328 13148 29348
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 13188 29170 13216 30126
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12360 27130 12388 28494
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12176 26846 12296 26874
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 11980 26444 12032 26450
rect 11980 26386 12032 26392
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11808 23526 11836 23802
rect 11900 23526 11928 24278
rect 11992 24274 12020 26386
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 12084 24274 12112 25910
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11624 20874 11652 21626
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11716 20466 11744 22714
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11808 18952 11836 23258
rect 11888 23248 11940 23254
rect 11886 23216 11888 23225
rect 11940 23216 11942 23225
rect 11886 23151 11942 23160
rect 12070 23216 12126 23225
rect 12070 23151 12126 23160
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11900 21622 11928 22510
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11900 20806 11928 21558
rect 11992 21350 12020 21830
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11808 18924 11928 18952
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11624 17338 11652 17614
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11716 16726 11744 17478
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11440 13688 11560 13716
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10810 11100 11086
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11256 10742 11284 10950
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11348 10266 11376 12718
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9648 11020 9654
rect 10966 9616 10968 9625
rect 11020 9616 11022 9625
rect 10966 9551 11022 9560
rect 10966 9480 11022 9489
rect 10966 9415 11022 9424
rect 10980 9382 11008 9415
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11072 9042 11100 10066
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11152 8968 11204 8974
rect 10966 8936 11022 8945
rect 11152 8910 11204 8916
rect 10966 8871 11022 8880
rect 10980 8566 11008 8871
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10980 7993 11008 8026
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 11072 7290 11100 8230
rect 10980 7274 11100 7290
rect 10968 7268 11100 7274
rect 11020 7262 11100 7268
rect 10968 7210 11020 7216
rect 11060 7200 11112 7206
rect 11164 7188 11192 8910
rect 11256 8430 11284 9318
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11112 7160 11192 7188
rect 11060 7142 11112 7148
rect 11072 6866 11100 7142
rect 11256 6984 11284 8026
rect 11164 6956 11284 6984
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10704 5166 10732 6326
rect 11164 6322 11192 6956
rect 11348 6882 11376 8434
rect 11256 6854 11376 6882
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10796 5030 10824 6190
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5914 11100 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10612 4814 10824 4842
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10336 3194 10364 3334
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10244 1414 10456 1442
rect 10428 800 10456 1414
rect 10796 800 10824 4814
rect 10980 4622 11008 5850
rect 11164 5846 11192 6258
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11164 5216 11192 5782
rect 11072 5188 11192 5216
rect 11072 5098 11100 5188
rect 11256 5166 11284 6854
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11244 5160 11296 5166
rect 11164 5108 11244 5114
rect 11164 5102 11296 5108
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11164 5086 11284 5102
rect 10968 4616 11020 4622
rect 10888 4576 10968 4604
rect 10888 3534 10916 4576
rect 10968 4558 11020 4564
rect 11164 3738 11192 5086
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 4146 11284 4558
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 2990 11008 3470
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 11164 2650 11192 3674
rect 11348 3534 11376 6666
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11440 2496 11468 13688
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11532 11218 11560 12174
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10606 11560 11154
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11624 10554 11652 14418
rect 11716 14074 11744 14758
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11716 10674 11744 14010
rect 11808 13734 11836 18770
rect 11900 14618 11928 18924
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11900 13462 11928 14554
rect 11992 14074 12020 20402
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10554 11836 10610
rect 11624 10526 11836 10554
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9353 11560 9862
rect 11518 9344 11574 9353
rect 11518 9279 11574 9288
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8022 11560 8910
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7546 11744 7754
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 6934 11652 7346
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11624 4078 11652 6394
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11440 2468 11560 2496
rect 11152 1012 11204 1018
rect 11152 954 11204 960
rect 11164 800 11192 954
rect 11532 800 11560 2468
rect 11808 800 11836 10526
rect 11900 9586 11928 11698
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10062 12020 10950
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 6458 11928 9522
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 8498 12020 9454
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 4826 12020 7754
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12084 1018 12112 23151
rect 12176 22080 12204 26846
rect 12452 23769 12480 26862
rect 12438 23760 12494 23769
rect 12438 23695 12494 23704
rect 12348 23656 12400 23662
rect 12400 23616 12480 23644
rect 12348 23598 12400 23604
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12254 23352 12310 23361
rect 12254 23287 12256 23296
rect 12308 23287 12310 23296
rect 12256 23258 12308 23264
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 12268 23089 12296 23122
rect 12254 23080 12310 23089
rect 12254 23015 12310 23024
rect 12256 22092 12308 22098
rect 12176 22052 12256 22080
rect 12256 22034 12308 22040
rect 12360 19258 12388 23462
rect 12452 23254 12480 23616
rect 12440 23248 12492 23254
rect 12544 23225 12572 28494
rect 12636 28218 12664 28562
rect 12852 28316 13148 28336
rect 12908 28314 12932 28316
rect 12988 28314 13012 28316
rect 13068 28314 13092 28316
rect 12930 28262 12932 28314
rect 12994 28262 13006 28314
rect 13068 28262 13070 28314
rect 12908 28260 12932 28262
rect 12988 28260 13012 28262
rect 13068 28260 13092 28262
rect 12852 28240 13148 28260
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12636 25838 12664 28154
rect 13280 27606 13308 41006
rect 13832 40390 13860 44390
rect 13912 44328 13964 44334
rect 14016 44282 14044 47058
rect 14200 46714 14228 47058
rect 14280 46912 14332 46918
rect 14280 46854 14332 46860
rect 14188 46708 14240 46714
rect 14188 46650 14240 46656
rect 14096 46504 14148 46510
rect 14096 46446 14148 46452
rect 14108 45830 14136 46446
rect 14292 46102 14320 46854
rect 14832 46572 14884 46578
rect 14832 46514 14884 46520
rect 14280 46096 14332 46102
rect 14280 46038 14332 46044
rect 14844 46034 14872 46514
rect 14832 46028 14884 46034
rect 14832 45970 14884 45976
rect 14096 45824 14148 45830
rect 14096 45766 14148 45772
rect 14844 45422 14872 45970
rect 14832 45416 14884 45422
rect 14832 45358 14884 45364
rect 15200 45416 15252 45422
rect 15200 45358 15252 45364
rect 14844 44878 14872 45358
rect 15212 45014 15240 45358
rect 15200 45008 15252 45014
rect 15200 44950 15252 44956
rect 14832 44872 14884 44878
rect 14832 44814 14884 44820
rect 13964 44276 14044 44282
rect 13912 44270 14044 44276
rect 13924 44254 14044 44270
rect 13924 42362 13952 44254
rect 14844 43790 14872 44814
rect 15304 44554 15332 49200
rect 15660 47116 15712 47122
rect 15660 47058 15712 47064
rect 15752 47116 15804 47122
rect 15752 47058 15804 47064
rect 15476 46912 15528 46918
rect 15476 46854 15528 46860
rect 15488 46510 15516 46854
rect 15476 46504 15528 46510
rect 15476 46446 15528 46452
rect 15384 46436 15436 46442
rect 15384 46378 15436 46384
rect 15212 44538 15332 44554
rect 15200 44532 15332 44538
rect 15252 44526 15332 44532
rect 15200 44474 15252 44480
rect 14096 43784 14148 43790
rect 14096 43726 14148 43732
rect 14832 43784 14884 43790
rect 14832 43726 14884 43732
rect 14108 43314 14136 43726
rect 14096 43308 14148 43314
rect 14096 43250 14148 43256
rect 14844 43246 14872 43726
rect 15304 43450 15332 44526
rect 15396 44402 15424 46378
rect 15488 45898 15516 46446
rect 15476 45892 15528 45898
rect 15476 45834 15528 45840
rect 15672 45490 15700 47058
rect 15660 45484 15712 45490
rect 15660 45426 15712 45432
rect 15476 44532 15528 44538
rect 15476 44474 15528 44480
rect 15384 44396 15436 44402
rect 15384 44338 15436 44344
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 14832 43240 14884 43246
rect 14832 43182 14884 43188
rect 14280 43104 14332 43110
rect 14280 43046 14332 43052
rect 13912 42356 13964 42362
rect 13912 42298 13964 42304
rect 14292 42158 14320 43046
rect 14844 42634 14872 43182
rect 15384 42764 15436 42770
rect 15384 42706 15436 42712
rect 14832 42628 14884 42634
rect 14832 42570 14884 42576
rect 14280 42152 14332 42158
rect 14280 42094 14332 42100
rect 14648 42152 14700 42158
rect 14648 42094 14700 42100
rect 14556 42084 14608 42090
rect 14556 42026 14608 42032
rect 14568 41818 14596 42026
rect 14556 41812 14608 41818
rect 14556 41754 14608 41760
rect 14464 41676 14516 41682
rect 14464 41618 14516 41624
rect 14280 41540 14332 41546
rect 14280 41482 14332 41488
rect 13820 40384 13872 40390
rect 13820 40326 13872 40332
rect 13912 40384 13964 40390
rect 13912 40326 13964 40332
rect 13924 40202 13952 40326
rect 13832 40174 13952 40202
rect 13832 39982 13860 40174
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 13820 39976 13872 39982
rect 13820 39918 13872 39924
rect 13452 37868 13504 37874
rect 13556 37856 13584 39918
rect 13832 39642 13860 39918
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 14096 39296 14148 39302
rect 14096 39238 14148 39244
rect 14108 38865 14136 39238
rect 14094 38856 14150 38865
rect 14094 38791 14150 38800
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13832 38486 13860 38694
rect 13820 38480 13872 38486
rect 13820 38422 13872 38428
rect 13504 37828 13584 37856
rect 13452 37810 13504 37816
rect 13360 36712 13412 36718
rect 13360 36654 13412 36660
rect 13372 36242 13400 36654
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13372 34950 13400 36178
rect 13464 36174 13492 37810
rect 13832 37806 13860 38422
rect 14108 37806 14136 38791
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 14096 37800 14148 37806
rect 14096 37742 14148 37748
rect 13832 37330 13860 37742
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 13636 36644 13688 36650
rect 13636 36586 13688 36592
rect 13544 36576 13596 36582
rect 13544 36518 13596 36524
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13360 34944 13412 34950
rect 13360 34886 13412 34892
rect 13556 32978 13584 36518
rect 13648 36242 13676 36586
rect 13832 36310 13860 37266
rect 13820 36304 13872 36310
rect 13820 36246 13872 36252
rect 13636 36236 13688 36242
rect 13636 36178 13688 36184
rect 13648 35154 13676 36178
rect 13636 35148 13688 35154
rect 13636 35090 13688 35096
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13372 31890 13400 32710
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13452 31952 13504 31958
rect 13452 31894 13504 31900
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13464 31362 13492 31894
rect 13556 31482 13584 32370
rect 13648 31890 13676 35090
rect 13832 35086 13860 36246
rect 14096 36236 14148 36242
rect 14096 36178 14148 36184
rect 14108 35578 14136 36178
rect 14016 35550 14136 35578
rect 13820 35080 13872 35086
rect 13820 35022 13872 35028
rect 13820 34944 13872 34950
rect 13872 34904 13952 34932
rect 13820 34886 13872 34892
rect 13924 32842 13952 34904
rect 14016 34542 14044 35550
rect 14004 34536 14056 34542
rect 14004 34478 14056 34484
rect 14016 33658 14044 34478
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 13912 32836 13964 32842
rect 13912 32778 13964 32784
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13464 31334 13584 31362
rect 13452 30660 13504 30666
rect 13452 30602 13504 30608
rect 13268 27600 13320 27606
rect 13268 27542 13320 27548
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12728 26518 12756 27338
rect 12852 27228 13148 27248
rect 12908 27226 12932 27228
rect 12988 27226 13012 27228
rect 13068 27226 13092 27228
rect 12930 27174 12932 27226
rect 12994 27174 13006 27226
rect 13068 27174 13070 27226
rect 12908 27172 12932 27174
rect 12988 27172 13012 27174
rect 13068 27172 13092 27174
rect 12852 27152 13148 27172
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12624 24744 12676 24750
rect 12622 24712 12624 24721
rect 12676 24712 12678 24721
rect 12728 24698 12756 26318
rect 12852 26140 13148 26160
rect 12908 26138 12932 26140
rect 12988 26138 13012 26140
rect 13068 26138 13092 26140
rect 12930 26086 12932 26138
rect 12994 26086 13006 26138
rect 13068 26086 13070 26138
rect 12908 26084 12932 26086
rect 12988 26084 13012 26086
rect 13068 26084 13092 26086
rect 12852 26064 13148 26084
rect 13280 25430 13308 27406
rect 13268 25424 13320 25430
rect 13268 25366 13320 25372
rect 12852 25052 13148 25072
rect 12908 25050 12932 25052
rect 12988 25050 13012 25052
rect 13068 25050 13092 25052
rect 12930 24998 12932 25050
rect 12994 24998 13006 25050
rect 13068 24998 13070 25050
rect 12908 24996 12932 24998
rect 12988 24996 13012 24998
rect 13068 24996 13092 24998
rect 12852 24976 13148 24996
rect 12678 24670 12756 24698
rect 13464 24682 13492 30602
rect 12622 24647 12678 24656
rect 12622 24032 12678 24041
rect 12622 23967 12678 23976
rect 12636 23526 12664 23967
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12440 23190 12492 23196
rect 12530 23216 12586 23225
rect 12530 23151 12586 23160
rect 12728 23118 12756 24670
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 12852 23964 13148 23984
rect 12908 23962 12932 23964
rect 12988 23962 13012 23964
rect 13068 23962 13092 23964
rect 12930 23910 12932 23962
rect 12994 23910 13006 23962
rect 13068 23910 13070 23962
rect 12908 23908 12932 23910
rect 12988 23908 13012 23910
rect 13068 23908 13092 23910
rect 12852 23888 13148 23908
rect 13556 23610 13584 31334
rect 13648 30258 13676 31826
rect 13832 31754 13860 32710
rect 13924 31754 13952 32778
rect 14108 32570 14136 32846
rect 14096 32564 14148 32570
rect 14096 32506 14148 32512
rect 14200 32230 14228 32914
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14200 31822 14228 32166
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 13820 31748 13872 31754
rect 13820 31690 13872 31696
rect 13912 31748 13964 31754
rect 13912 31690 13964 31696
rect 14200 31482 14228 31758
rect 14188 31476 14240 31482
rect 14188 31418 14240 31424
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 13636 30252 13688 30258
rect 13636 30194 13688 30200
rect 13924 29714 13952 31078
rect 14004 30796 14056 30802
rect 14004 30738 14056 30744
rect 14016 30326 14044 30738
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14004 30320 14056 30326
rect 14004 30262 14056 30268
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13912 29708 13964 29714
rect 13964 29668 14044 29696
rect 13912 29650 13964 29656
rect 13740 28694 13768 29650
rect 13728 28688 13780 28694
rect 13728 28630 13780 28636
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13924 28082 13952 28358
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13728 26444 13780 26450
rect 13728 26386 13780 26392
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13084 23588 13136 23594
rect 13084 23530 13136 23536
rect 13280 23582 13584 23610
rect 13096 23322 13124 23530
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12852 22876 13148 22896
rect 12908 22874 12932 22876
rect 12988 22874 13012 22876
rect 13068 22874 13092 22876
rect 12930 22822 12932 22874
rect 12994 22822 13006 22874
rect 13068 22822 13070 22874
rect 12908 22820 12932 22822
rect 12988 22820 13012 22822
rect 13068 22820 13092 22822
rect 12852 22800 13148 22820
rect 13280 22778 13308 23582
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13372 23050 13400 23462
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13452 23044 13504 23050
rect 13452 22986 13504 22992
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 12852 21788 13148 21808
rect 12908 21786 12932 21788
rect 12988 21786 13012 21788
rect 13068 21786 13092 21788
rect 12930 21734 12932 21786
rect 12994 21734 13006 21786
rect 13068 21734 13070 21786
rect 12908 21732 12932 21734
rect 12988 21732 13012 21734
rect 13068 21732 13092 21734
rect 12852 21712 13148 21732
rect 13188 21554 13216 22578
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 21078 12756 21422
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12820 20890 12848 20946
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12728 20862 12848 20890
rect 12176 19230 12388 19258
rect 12176 18986 12204 19230
rect 12176 18958 12296 18986
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 16998 12204 17614
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16114 12204 16934
rect 12268 16250 12296 18958
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12452 17202 12480 17818
rect 12544 17202 12572 20810
rect 12636 19922 12664 20810
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12176 15570 12204 16050
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12176 14550 12204 14894
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12268 14482 12296 15982
rect 12452 15366 12480 17002
rect 12544 15586 12572 17138
rect 12636 17134 12664 18770
rect 12728 18290 12756 20862
rect 12852 20700 13148 20720
rect 12908 20698 12932 20700
rect 12988 20698 13012 20700
rect 13068 20698 13092 20700
rect 12930 20646 12932 20698
rect 12994 20646 13006 20698
rect 13068 20646 13070 20698
rect 12908 20644 12932 20646
rect 12988 20644 13012 20646
rect 13068 20644 13092 20646
rect 12852 20624 13148 20644
rect 13188 20058 13216 21354
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20466 13400 20946
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 12852 19612 13148 19632
rect 12908 19610 12932 19612
rect 12988 19610 13012 19612
rect 13068 19610 13092 19612
rect 12930 19558 12932 19610
rect 12994 19558 13006 19610
rect 13068 19558 13070 19610
rect 12908 19556 12932 19558
rect 12988 19556 13012 19558
rect 13068 19556 13092 19558
rect 12852 19536 13148 19556
rect 13372 19514 13400 20402
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 12852 18524 13148 18544
rect 12908 18522 12932 18524
rect 12988 18522 13012 18524
rect 13068 18522 13092 18524
rect 12930 18470 12932 18522
rect 12994 18470 13006 18522
rect 13068 18470 13070 18522
rect 12908 18468 12932 18470
rect 12988 18468 13012 18470
rect 13068 18468 13092 18470
rect 12852 18448 13148 18468
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 13188 17610 13216 19178
rect 13372 18358 13400 19246
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13464 18170 13492 22986
rect 13556 22234 13584 23122
rect 13648 23050 13676 25298
rect 13740 24342 13768 26386
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 19990 13676 22714
rect 13740 22574 13768 23598
rect 13832 23526 13860 27338
rect 14016 27010 14044 29668
rect 13924 26982 14044 27010
rect 13924 24290 13952 26982
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14016 26042 14044 26862
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 13924 24262 14044 24290
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13924 23730 13952 24142
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 14016 22710 14044 24262
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13556 19718 13584 19926
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13648 18834 13676 19926
rect 13740 19310 13768 22510
rect 14108 21457 14136 30534
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14200 24750 14228 26930
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21690 14228 21830
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14094 21448 14150 21457
rect 14094 21383 14150 21392
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13740 18970 13768 19246
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 14200 18834 14228 19178
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13280 18142 13492 18170
rect 13636 18148 13688 18154
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 12852 17436 13148 17456
rect 12908 17434 12932 17436
rect 12988 17434 13012 17436
rect 13068 17434 13092 17436
rect 12930 17382 12932 17434
rect 12994 17382 13006 17434
rect 13068 17382 13070 17434
rect 12908 17380 12932 17382
rect 12988 17380 13012 17382
rect 13068 17380 13092 17382
rect 12852 17360 13148 17380
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12852 16348 13148 16368
rect 12908 16346 12932 16348
rect 12988 16346 13012 16348
rect 13068 16346 13092 16348
rect 12930 16294 12932 16346
rect 12994 16294 13006 16346
rect 13068 16294 13070 16346
rect 12908 16292 12932 16294
rect 12988 16292 13012 16294
rect 13068 16292 13092 16294
rect 12852 16272 13148 16292
rect 13188 16232 13216 17546
rect 13280 16658 13308 18142
rect 13636 18090 13688 18096
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13096 16204 13216 16232
rect 13096 15722 13124 16204
rect 13280 15994 13308 16594
rect 13372 16454 13400 17614
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13188 15966 13308 15994
rect 13464 15978 13492 16526
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13452 15972 13504 15978
rect 13188 15910 13216 15966
rect 13452 15914 13504 15920
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13096 15694 13216 15722
rect 12544 15558 12664 15586
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12544 14414 12572 15438
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 11694 12204 13670
rect 12360 12306 12388 14010
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 7857 12204 11018
rect 12268 10130 12296 12038
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12360 10713 12388 11766
rect 12452 11676 12480 12718
rect 12544 12374 12572 13942
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12532 11688 12584 11694
rect 12452 11648 12532 11676
rect 12532 11630 12584 11636
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12452 11082 12480 11494
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12438 10976 12494 10985
rect 12438 10911 12494 10920
rect 12346 10704 12402 10713
rect 12346 10639 12402 10648
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12452 10062 12480 10911
rect 12544 10606 12572 11494
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12636 10452 12664 15558
rect 12852 15260 13148 15280
rect 12908 15258 12932 15260
rect 12988 15258 13012 15260
rect 13068 15258 13092 15260
rect 12930 15206 12932 15258
rect 12994 15206 13006 15258
rect 13068 15206 13070 15258
rect 12908 15204 12932 15206
rect 12988 15204 13012 15206
rect 13068 15204 13092 15206
rect 12852 15184 13148 15204
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 11257 12756 14894
rect 13188 14770 13216 15694
rect 13556 15094 13584 15982
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13648 15026 13676 18090
rect 13740 17626 13768 18294
rect 13924 18222 13952 18702
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17746 13860 18022
rect 13924 17814 13952 18158
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13740 17598 13860 17626
rect 13832 17542 13860 17598
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16658 13768 17070
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13268 14952 13320 14958
rect 13320 14912 13400 14940
rect 13268 14894 13320 14900
rect 13188 14742 13308 14770
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12912 14346 12940 14486
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12852 14172 13148 14192
rect 12908 14170 12932 14172
rect 12988 14170 13012 14172
rect 13068 14170 13092 14172
rect 12930 14118 12932 14170
rect 12994 14118 13006 14170
rect 13068 14118 13070 14170
rect 12908 14116 12932 14118
rect 12988 14116 13012 14118
rect 13068 14116 13092 14118
rect 12852 14096 13148 14116
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13188 13258 13216 13806
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13280 13138 13308 14742
rect 13372 14006 13400 14912
rect 13648 14362 13676 14962
rect 13740 14550 13768 16594
rect 14292 16454 14320 41482
rect 14476 41070 14504 41618
rect 14660 41614 14688 42094
rect 14648 41608 14700 41614
rect 14648 41550 14700 41556
rect 14844 41546 14872 42570
rect 15396 41682 15424 42706
rect 15488 42294 15516 44474
rect 15660 44328 15712 44334
rect 15660 44270 15712 44276
rect 15568 42560 15620 42566
rect 15568 42502 15620 42508
rect 15476 42288 15528 42294
rect 15476 42230 15528 42236
rect 15580 41682 15608 42502
rect 15384 41676 15436 41682
rect 15384 41618 15436 41624
rect 15568 41676 15620 41682
rect 15568 41618 15620 41624
rect 14832 41540 14884 41546
rect 14832 41482 14884 41488
rect 14372 41064 14424 41070
rect 14372 41006 14424 41012
rect 14464 41064 14516 41070
rect 14464 41006 14516 41012
rect 14384 30716 14412 41006
rect 14476 39506 14504 41006
rect 14844 39522 14872 41482
rect 15396 40662 15424 41618
rect 15384 40656 15436 40662
rect 15384 40598 15436 40604
rect 14924 40384 14976 40390
rect 14924 40326 14976 40332
rect 14936 39982 14964 40326
rect 15396 40186 15424 40598
rect 15384 40180 15436 40186
rect 15384 40122 15436 40128
rect 15200 40044 15252 40050
rect 15200 39986 15252 39992
rect 14924 39976 14976 39982
rect 14924 39918 14976 39924
rect 14464 39500 14516 39506
rect 14844 39494 14964 39522
rect 15212 39506 15240 39986
rect 15396 39914 15424 40122
rect 15384 39908 15436 39914
rect 15384 39850 15436 39856
rect 14464 39442 14516 39448
rect 14476 38418 14504 39442
rect 14832 39364 14884 39370
rect 14832 39306 14884 39312
rect 14464 38412 14516 38418
rect 14464 38354 14516 38360
rect 14476 37466 14504 38354
rect 14556 38344 14608 38350
rect 14556 38286 14608 38292
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 14464 36780 14516 36786
rect 14464 36722 14516 36728
rect 14476 35222 14504 36722
rect 14464 35216 14516 35222
rect 14464 35158 14516 35164
rect 14464 35080 14516 35086
rect 14464 35022 14516 35028
rect 14476 30938 14504 35022
rect 14464 30932 14516 30938
rect 14464 30874 14516 30880
rect 14384 30688 14504 30716
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23798 14412 24006
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14384 22098 14412 22374
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19514 14412 20334
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13556 14334 13676 14362
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13188 13110 13308 13138
rect 12852 13084 13148 13104
rect 12908 13082 12932 13084
rect 12988 13082 13012 13084
rect 13068 13082 13092 13084
rect 12930 13030 12932 13082
rect 12994 13030 13006 13082
rect 13068 13030 13070 13082
rect 12908 13028 12932 13030
rect 12988 13028 13012 13030
rect 13068 13028 13092 13030
rect 12852 13008 13148 13028
rect 12852 11996 13148 12016
rect 12908 11994 12932 11996
rect 12988 11994 13012 11996
rect 13068 11994 13092 11996
rect 12930 11942 12932 11994
rect 12994 11942 13006 11994
rect 13068 11942 13070 11994
rect 12908 11940 12932 11942
rect 12988 11940 13012 11942
rect 13068 11940 13092 11942
rect 12852 11920 13148 11940
rect 12714 11248 12770 11257
rect 12714 11183 12770 11192
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12544 10424 12664 10452
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9920 12400 9926
rect 12452 9897 12480 9998
rect 12348 9862 12400 9868
rect 12438 9888 12494 9897
rect 12360 9042 12388 9862
rect 12438 9823 12494 9832
rect 12544 9738 12572 10424
rect 12544 9710 12664 9738
rect 12440 9104 12492 9110
rect 12438 9072 12440 9081
rect 12492 9072 12494 9081
rect 12348 9036 12400 9042
rect 12438 9007 12494 9016
rect 12348 8978 12400 8984
rect 12532 8968 12584 8974
rect 12254 8936 12310 8945
rect 12532 8910 12584 8916
rect 12254 8871 12310 8880
rect 12268 8090 12296 8871
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8424 12400 8430
rect 12452 8401 12480 8774
rect 12348 8366 12400 8372
rect 12438 8392 12494 8401
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12162 7848 12218 7857
rect 12360 7818 12388 8366
rect 12438 8327 12494 8336
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12162 7783 12218 7792
rect 12348 7812 12400 7818
rect 12176 7002 12204 7783
rect 12348 7754 12400 7760
rect 12452 7274 12480 8026
rect 12544 7478 12572 8910
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12544 7002 12572 7414
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12176 4622 12204 4966
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12162 4448 12218 4457
rect 12162 4383 12218 4392
rect 12072 1012 12124 1018
rect 12072 954 12124 960
rect 12176 800 12204 4383
rect 12360 2990 12388 5102
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12452 2514 12480 3062
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12544 800 12572 6802
rect 12636 2938 12664 9710
rect 12728 8362 12756 11086
rect 12852 10908 13148 10928
rect 12908 10906 12932 10908
rect 12988 10906 13012 10908
rect 13068 10906 13092 10908
rect 12930 10854 12932 10906
rect 12994 10854 13006 10906
rect 13068 10854 13070 10906
rect 12908 10852 12932 10854
rect 12988 10852 13012 10854
rect 13068 10852 13092 10854
rect 12852 10832 13148 10852
rect 12852 9820 13148 9840
rect 12908 9818 12932 9820
rect 12988 9818 13012 9820
rect 13068 9818 13092 9820
rect 12930 9766 12932 9818
rect 12994 9766 13006 9818
rect 13068 9766 13070 9818
rect 12908 9764 12932 9766
rect 12988 9764 13012 9766
rect 13068 9764 13092 9766
rect 12852 9744 13148 9764
rect 12898 9344 12954 9353
rect 12898 9279 12954 9288
rect 12912 9042 12940 9279
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12852 8732 13148 8752
rect 12908 8730 12932 8732
rect 12988 8730 13012 8732
rect 13068 8730 13092 8732
rect 12930 8678 12932 8730
rect 12994 8678 13006 8730
rect 13068 8678 13070 8730
rect 12908 8676 12932 8678
rect 12988 8676 13012 8678
rect 13068 8676 13092 8678
rect 12852 8656 13148 8676
rect 13082 8392 13138 8401
rect 12716 8356 12768 8362
rect 13082 8327 13138 8336
rect 12716 8298 12768 8304
rect 12728 8090 12756 8298
rect 12898 8120 12954 8129
rect 12716 8084 12768 8090
rect 12898 8055 12954 8064
rect 12716 8026 12768 8032
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12728 6934 12756 7890
rect 12820 7818 12848 7890
rect 12912 7886 12940 8055
rect 13096 7954 13124 8327
rect 13188 8265 13216 13110
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13280 12442 13308 12718
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13372 12306 13400 13942
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11218 13400 11494
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 9994 13308 10542
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8634 13308 8774
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8514 13400 11154
rect 13280 8498 13400 8514
rect 13268 8492 13400 8498
rect 13320 8486 13400 8492
rect 13268 8434 13320 8440
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13268 8288 13320 8294
rect 13174 8256 13230 8265
rect 13268 8230 13320 8236
rect 13174 8191 13230 8200
rect 13280 8090 13308 8230
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13084 7948 13136 7954
rect 13136 7908 13216 7936
rect 13084 7890 13136 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12852 7644 13148 7664
rect 12908 7642 12932 7644
rect 12988 7642 13012 7644
rect 13068 7642 13092 7644
rect 12930 7590 12932 7642
rect 12994 7590 13006 7642
rect 13068 7590 13070 7642
rect 12908 7588 12932 7590
rect 12988 7588 13012 7590
rect 13068 7588 13092 7590
rect 12852 7568 13148 7588
rect 13188 7410 13216 7908
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12820 7206 12848 7346
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12716 6792 12768 6798
rect 12820 6780 12848 6938
rect 13372 6866 13400 8366
rect 13464 8129 13492 12922
rect 13450 8120 13506 8129
rect 13450 8055 13506 8064
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 12768 6752 12848 6780
rect 13176 6792 13228 6798
rect 12716 6734 12768 6740
rect 13176 6734 13228 6740
rect 12728 5166 12756 6734
rect 12852 6556 13148 6576
rect 12908 6554 12932 6556
rect 12988 6554 13012 6556
rect 13068 6554 13092 6556
rect 12930 6502 12932 6554
rect 12994 6502 13006 6554
rect 13068 6502 13070 6554
rect 12908 6500 12932 6502
rect 12988 6500 13012 6502
rect 13068 6500 13092 6502
rect 12852 6480 13148 6500
rect 13188 6458 13216 6734
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13280 5778 13308 6394
rect 13360 6316 13412 6322
rect 13464 6304 13492 8055
rect 13412 6276 13492 6304
rect 13360 6258 13412 6264
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13372 5710 13400 6258
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13360 5704 13412 5710
rect 13280 5652 13360 5658
rect 13280 5646 13412 5652
rect 13280 5630 13400 5646
rect 12852 5468 13148 5488
rect 12908 5466 12932 5468
rect 12988 5466 13012 5468
rect 13068 5466 13092 5468
rect 12930 5414 12932 5466
rect 12994 5414 13006 5466
rect 13068 5414 13070 5466
rect 12908 5412 12932 5414
rect 12988 5412 13012 5414
rect 13068 5412 13092 5414
rect 12852 5392 13148 5412
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 12852 4380 13148 4400
rect 12908 4378 12932 4380
rect 12988 4378 13012 4380
rect 13068 4378 13092 4380
rect 12930 4326 12932 4378
rect 12994 4326 13006 4378
rect 13068 4326 13070 4378
rect 12908 4324 12932 4326
rect 12988 4324 13012 4326
rect 13068 4324 13092 4326
rect 12852 4304 13148 4324
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3602 13032 4082
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3738 13124 4014
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13188 3516 13216 4762
rect 13280 4146 13308 5630
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5234 13400 5510
rect 13464 5370 13492 6122
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13372 4078 13400 4626
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13268 3528 13320 3534
rect 13188 3488 13268 3516
rect 13268 3470 13320 3476
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 3058 12756 3334
rect 12852 3292 13148 3312
rect 12908 3290 12932 3292
rect 12988 3290 13012 3292
rect 13068 3290 13092 3292
rect 12930 3238 12932 3290
rect 12994 3238 13006 3290
rect 13068 3238 13070 3290
rect 12908 3236 12932 3238
rect 12988 3236 13012 3238
rect 13068 3236 13092 3238
rect 12852 3216 13148 3236
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12636 2910 12756 2938
rect 12728 1358 12756 2910
rect 12852 2204 13148 2224
rect 12908 2202 12932 2204
rect 12988 2202 13012 2204
rect 13068 2202 13092 2204
rect 12930 2150 12932 2202
rect 12994 2150 13006 2202
rect 13068 2150 13070 2202
rect 12908 2148 12932 2150
rect 12988 2148 13012 2150
rect 13068 2148 13092 2150
rect 12852 2128 13148 2148
rect 13556 1442 13584 14334
rect 13924 14278 13952 15438
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13648 13530 13676 14214
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 13190 13676 13330
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13740 12986 13768 13670
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13924 12306 13952 14214
rect 14384 13734 14412 17818
rect 14476 15706 14504 30688
rect 14568 25906 14596 38286
rect 14648 36712 14700 36718
rect 14648 36654 14700 36660
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 14660 35290 14688 36654
rect 14752 36174 14780 36654
rect 14740 36168 14792 36174
rect 14740 36110 14792 36116
rect 14648 35284 14700 35290
rect 14648 35226 14700 35232
rect 14752 35086 14780 36110
rect 14740 35080 14792 35086
rect 14740 35022 14792 35028
rect 14740 33924 14792 33930
rect 14740 33866 14792 33872
rect 14648 30932 14700 30938
rect 14648 30874 14700 30880
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14660 24834 14688 30874
rect 14752 27044 14780 33866
rect 14844 31770 14872 39306
rect 14936 37398 14964 39494
rect 15200 39500 15252 39506
rect 15200 39442 15252 39448
rect 15384 39500 15436 39506
rect 15384 39442 15436 39448
rect 15108 37800 15160 37806
rect 15108 37742 15160 37748
rect 14924 37392 14976 37398
rect 14924 37334 14976 37340
rect 14936 35630 14964 37334
rect 15120 36786 15148 37742
rect 15212 36922 15240 39442
rect 15292 37732 15344 37738
rect 15292 37674 15344 37680
rect 15304 37330 15332 37674
rect 15292 37324 15344 37330
rect 15292 37266 15344 37272
rect 15396 37210 15424 39442
rect 15672 39438 15700 44270
rect 15660 39432 15712 39438
rect 15660 39374 15712 39380
rect 15764 38486 15792 47058
rect 16132 46374 16160 49200
rect 16960 47546 16988 49200
rect 16592 47518 16988 47546
rect 16212 47048 16264 47054
rect 16212 46990 16264 46996
rect 16120 46368 16172 46374
rect 16120 46310 16172 46316
rect 15936 45824 15988 45830
rect 15936 45766 15988 45772
rect 15948 44470 15976 45766
rect 16132 45626 16160 46310
rect 16120 45620 16172 45626
rect 16120 45562 16172 45568
rect 16224 44946 16252 46990
rect 16212 44940 16264 44946
rect 16212 44882 16264 44888
rect 15936 44464 15988 44470
rect 15936 44406 15988 44412
rect 16304 44260 16356 44266
rect 16304 44202 16356 44208
rect 16316 43858 16344 44202
rect 16304 43852 16356 43858
rect 16304 43794 16356 43800
rect 16592 43466 16620 47518
rect 16817 47356 17113 47376
rect 16873 47354 16897 47356
rect 16953 47354 16977 47356
rect 17033 47354 17057 47356
rect 16895 47302 16897 47354
rect 16959 47302 16971 47354
rect 17033 47302 17035 47354
rect 16873 47300 16897 47302
rect 16953 47300 16977 47302
rect 17033 47300 17057 47302
rect 16817 47280 17113 47300
rect 17696 46714 17724 49200
rect 18524 47546 18552 49200
rect 18248 47518 18552 47546
rect 17684 46708 17736 46714
rect 17684 46650 17736 46656
rect 17132 46504 17184 46510
rect 17132 46446 17184 46452
rect 16672 46436 16724 46442
rect 16672 46378 16724 46384
rect 16684 46034 16712 46378
rect 16817 46268 17113 46288
rect 16873 46266 16897 46268
rect 16953 46266 16977 46268
rect 17033 46266 17057 46268
rect 16895 46214 16897 46266
rect 16959 46214 16971 46266
rect 17033 46214 17035 46266
rect 16873 46212 16897 46214
rect 16953 46212 16977 46214
rect 17033 46212 17057 46214
rect 16817 46192 17113 46212
rect 16672 46028 16724 46034
rect 16672 45970 16724 45976
rect 16817 45180 17113 45200
rect 16873 45178 16897 45180
rect 16953 45178 16977 45180
rect 17033 45178 17057 45180
rect 16895 45126 16897 45178
rect 16959 45126 16971 45178
rect 17033 45126 17035 45178
rect 16873 45124 16897 45126
rect 16953 45124 16977 45126
rect 17033 45124 17057 45126
rect 16817 45104 17113 45124
rect 16817 44092 17113 44112
rect 16873 44090 16897 44092
rect 16953 44090 16977 44092
rect 17033 44090 17057 44092
rect 16895 44038 16897 44090
rect 16959 44038 16971 44090
rect 17033 44038 17035 44090
rect 16873 44036 16897 44038
rect 16953 44036 16977 44038
rect 17033 44036 17057 44038
rect 16817 44016 17113 44036
rect 16500 43438 16620 43466
rect 16500 43110 16528 43438
rect 16488 43104 16540 43110
rect 16488 43046 16540 43052
rect 16817 43004 17113 43024
rect 16873 43002 16897 43004
rect 16953 43002 16977 43004
rect 17033 43002 17057 43004
rect 16895 42950 16897 43002
rect 16959 42950 16971 43002
rect 17033 42950 17035 43002
rect 16873 42948 16897 42950
rect 16953 42948 16977 42950
rect 17033 42948 17057 42950
rect 16817 42928 17113 42948
rect 16120 42696 16172 42702
rect 16120 42638 16172 42644
rect 17040 42696 17092 42702
rect 17040 42638 17092 42644
rect 16028 42288 16080 42294
rect 16028 42230 16080 42236
rect 16040 41070 16068 42230
rect 16132 42090 16160 42638
rect 16580 42628 16632 42634
rect 16580 42570 16632 42576
rect 16212 42152 16264 42158
rect 16212 42094 16264 42100
rect 16120 42084 16172 42090
rect 16120 42026 16172 42032
rect 16224 41206 16252 42094
rect 16592 41614 16620 42570
rect 17052 42226 17080 42638
rect 17040 42220 17092 42226
rect 17040 42162 17092 42168
rect 16672 42084 16724 42090
rect 16672 42026 16724 42032
rect 16684 41682 16712 42026
rect 16817 41916 17113 41936
rect 16873 41914 16897 41916
rect 16953 41914 16977 41916
rect 17033 41914 17057 41916
rect 16895 41862 16897 41914
rect 16959 41862 16971 41914
rect 17033 41862 17035 41914
rect 16873 41860 16897 41862
rect 16953 41860 16977 41862
rect 17033 41860 17057 41862
rect 16817 41840 17113 41860
rect 16672 41676 16724 41682
rect 16672 41618 16724 41624
rect 16580 41608 16632 41614
rect 16580 41550 16632 41556
rect 16212 41200 16264 41206
rect 16212 41142 16264 41148
rect 16028 41064 16080 41070
rect 16028 41006 16080 41012
rect 16212 41064 16264 41070
rect 16212 41006 16264 41012
rect 16040 39964 16068 41006
rect 16120 40996 16172 41002
rect 16120 40938 16172 40944
rect 16132 40662 16160 40938
rect 16120 40656 16172 40662
rect 16120 40598 16172 40604
rect 16120 39976 16172 39982
rect 16040 39936 16120 39964
rect 16120 39918 16172 39924
rect 15844 38888 15896 38894
rect 15844 38830 15896 38836
rect 15752 38480 15804 38486
rect 15752 38422 15804 38428
rect 15856 38418 15884 38830
rect 16132 38758 16160 39918
rect 16224 38962 16252 41006
rect 16592 40526 16620 41550
rect 17144 41274 17172 46446
rect 17960 46436 18012 46442
rect 17960 46378 18012 46384
rect 17868 44328 17920 44334
rect 17868 44270 17920 44276
rect 17880 42158 17908 44270
rect 17972 43926 18000 46378
rect 18248 46102 18276 47518
rect 19260 47410 19288 49200
rect 18340 47382 19288 47410
rect 18236 46096 18288 46102
rect 18236 46038 18288 46044
rect 18340 45422 18368 47382
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 18420 46708 18472 46714
rect 18420 46650 18472 46656
rect 18144 45416 18196 45422
rect 18144 45358 18196 45364
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 18052 45348 18104 45354
rect 18052 45290 18104 45296
rect 17960 43920 18012 43926
rect 17960 43862 18012 43868
rect 17972 43246 18000 43862
rect 17960 43240 18012 43246
rect 17960 43182 18012 43188
rect 18064 43178 18092 45290
rect 18156 45014 18184 45358
rect 18144 45008 18196 45014
rect 18144 44950 18196 44956
rect 18328 44396 18380 44402
rect 18328 44338 18380 44344
rect 18340 43450 18368 44338
rect 18328 43444 18380 43450
rect 18328 43386 18380 43392
rect 18052 43172 18104 43178
rect 18052 43114 18104 43120
rect 18064 42362 18092 43114
rect 18328 42764 18380 42770
rect 18328 42706 18380 42712
rect 18052 42356 18104 42362
rect 18052 42298 18104 42304
rect 17868 42152 17920 42158
rect 17868 42094 17920 42100
rect 17132 41268 17184 41274
rect 17132 41210 17184 41216
rect 16672 40996 16724 41002
rect 16672 40938 16724 40944
rect 16684 40594 16712 40938
rect 16817 40828 17113 40848
rect 16873 40826 16897 40828
rect 16953 40826 16977 40828
rect 17033 40826 17057 40828
rect 16895 40774 16897 40826
rect 16959 40774 16971 40826
rect 17033 40774 17035 40826
rect 16873 40772 16897 40774
rect 16953 40772 16977 40774
rect 17033 40772 17057 40774
rect 16817 40752 17113 40772
rect 16672 40588 16724 40594
rect 16672 40530 16724 40536
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 16304 39976 16356 39982
rect 16304 39918 16356 39924
rect 16212 38956 16264 38962
rect 16212 38898 16264 38904
rect 16120 38752 16172 38758
rect 16120 38694 16172 38700
rect 15568 38412 15620 38418
rect 15568 38354 15620 38360
rect 15844 38412 15896 38418
rect 15844 38354 15896 38360
rect 15304 37182 15424 37210
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15108 36780 15160 36786
rect 15108 36722 15160 36728
rect 15016 36712 15068 36718
rect 15016 36654 15068 36660
rect 15028 36242 15056 36654
rect 15108 36644 15160 36650
rect 15108 36586 15160 36592
rect 15016 36236 15068 36242
rect 15016 36178 15068 36184
rect 15028 35850 15056 36178
rect 15120 35986 15148 36586
rect 15304 36106 15332 37182
rect 15476 36712 15528 36718
rect 15476 36654 15528 36660
rect 15384 36372 15436 36378
rect 15384 36314 15436 36320
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15120 35958 15240 35986
rect 15028 35834 15148 35850
rect 15028 35828 15160 35834
rect 15028 35822 15108 35828
rect 15108 35770 15160 35776
rect 15212 35698 15240 35958
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 14924 35624 14976 35630
rect 14924 35566 14976 35572
rect 14936 35494 14964 35566
rect 14924 35488 14976 35494
rect 14924 35430 14976 35436
rect 15304 35018 15332 36042
rect 15292 35012 15344 35018
rect 15292 34954 15344 34960
rect 15292 33924 15344 33930
rect 15292 33866 15344 33872
rect 14924 33448 14976 33454
rect 14924 33390 14976 33396
rect 14936 31890 14964 33390
rect 15016 33312 15068 33318
rect 15016 33254 15068 33260
rect 15028 32978 15056 33254
rect 15200 33040 15252 33046
rect 15200 32982 15252 32988
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 14844 31742 15056 31770
rect 14752 27016 14872 27044
rect 14568 24806 14688 24834
rect 14568 23594 14596 24806
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14660 23798 14688 24686
rect 14752 24274 14780 24686
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14646 23624 14702 23633
rect 14556 23588 14608 23594
rect 14646 23559 14702 23568
rect 14556 23530 14608 23536
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14568 22234 14596 22374
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14660 20058 14688 23559
rect 14844 22642 14872 27016
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14752 21554 14780 22442
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 16522 14688 19654
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14568 15638 14596 16390
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14660 14822 14688 15642
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 12918 14412 13670
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13648 10266 13676 11086
rect 13740 10554 13768 12106
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14016 11150 14044 11630
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13912 10600 13964 10606
rect 13740 10526 13860 10554
rect 13912 10542 13964 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13648 10084 13728 10112
rect 13648 9518 13676 10084
rect 13728 10066 13780 10072
rect 13832 10010 13860 10526
rect 13924 10470 13952 10542
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13740 9982 13860 10010
rect 13740 9586 13768 9982
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13740 8650 13768 9522
rect 13820 9036 13872 9042
rect 13924 9024 13952 10202
rect 14016 9926 14044 11086
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13872 8996 13952 9024
rect 13820 8978 13872 8984
rect 13648 8622 13768 8650
rect 13648 8022 13676 8622
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13740 7478 13768 8434
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 4758 13768 7142
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13634 4176 13690 4185
rect 13634 4111 13690 4120
rect 12912 1414 13584 1442
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 12912 800 12940 1414
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13280 800 13308 1294
rect 13648 800 13676 4111
rect 13740 4078 13768 4694
rect 13832 4690 13860 8502
rect 13924 6798 13952 8996
rect 14016 8974 14044 9862
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14016 8566 14044 8910
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6254 13952 6598
rect 14016 6322 14044 8366
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14016 5642 14044 6258
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13832 3602 13860 4626
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 3602 14044 4558
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13832 3126 13860 3538
rect 14108 3482 14136 11018
rect 14476 10742 14504 11630
rect 14752 11082 14780 21490
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14844 14958 14872 17070
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14936 14498 14964 24142
rect 15028 16114 15056 31742
rect 15212 30938 15240 32982
rect 15304 32026 15332 33866
rect 15396 32910 15424 36314
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15396 32434 15424 32710
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 15304 31822 15332 31962
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15304 30818 15332 31758
rect 15384 31204 15436 31210
rect 15384 31146 15436 31152
rect 15212 30790 15332 30818
rect 15212 29714 15240 30790
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15212 29322 15240 29650
rect 15120 29294 15240 29322
rect 15120 28762 15148 29294
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 15108 28756 15160 28762
rect 15108 28698 15160 28704
rect 15212 28626 15240 29174
rect 15304 29034 15332 30602
rect 15396 30598 15424 31146
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 15396 29034 15424 30534
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15384 29028 15436 29034
rect 15384 28970 15436 28976
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15200 28620 15252 28626
rect 15200 28562 15252 28568
rect 15212 27538 15240 28562
rect 15396 28014 15424 28698
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15212 26450 15240 26726
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 15304 25838 15332 27542
rect 15396 27538 15424 27950
rect 15384 27532 15436 27538
rect 15384 27474 15436 27480
rect 15396 26994 15424 27474
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15396 26382 15424 26930
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15120 23594 15148 23734
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15120 20602 15148 23530
rect 15212 23050 15240 25638
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15304 21894 15332 25774
rect 15396 25430 15424 25842
rect 15384 25424 15436 25430
rect 15384 25366 15436 25372
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15304 20330 15332 20946
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14844 14470 14964 14498
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14200 7410 14228 9862
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14292 7342 14320 8366
rect 14568 8022 14596 9046
rect 14660 8498 14688 9522
rect 14738 9208 14794 9217
rect 14738 9143 14794 9152
rect 14752 8498 14780 9143
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14556 8016 14608 8022
rect 14370 7984 14426 7993
rect 14556 7958 14608 7964
rect 14370 7919 14372 7928
rect 14424 7919 14426 7928
rect 14372 7890 14424 7896
rect 14464 7880 14516 7886
rect 14462 7848 14464 7857
rect 14516 7848 14518 7857
rect 14462 7783 14518 7792
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14292 7002 14320 7278
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 4758 14228 6734
rect 14292 6322 14320 6938
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14568 5710 14596 7958
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14476 5302 14504 5646
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14844 4826 14872 14470
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 7750 14964 8366
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15120 6254 15148 16458
rect 15212 14618 15240 18770
rect 15304 18086 15332 18770
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 15450 15332 18022
rect 15396 16130 15424 25230
rect 15488 19310 15516 36654
rect 15580 32994 15608 38354
rect 15856 37754 15884 38354
rect 16316 38350 16344 39918
rect 16488 39908 16540 39914
rect 16488 39850 16540 39856
rect 16396 38820 16448 38826
rect 16396 38762 16448 38768
rect 16304 38344 16356 38350
rect 16304 38286 16356 38292
rect 16212 38208 16264 38214
rect 16212 38150 16264 38156
rect 15764 37726 15884 37754
rect 16028 37800 16080 37806
rect 16028 37742 16080 37748
rect 15764 37670 15792 37726
rect 15752 37664 15804 37670
rect 15752 37606 15804 37612
rect 15764 36650 15792 37606
rect 16040 37126 16068 37742
rect 16224 37738 16252 38150
rect 16304 37800 16356 37806
rect 16304 37742 16356 37748
rect 16212 37732 16264 37738
rect 16212 37674 16264 37680
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 15936 36916 15988 36922
rect 15936 36858 15988 36864
rect 15752 36644 15804 36650
rect 15752 36586 15804 36592
rect 15764 34542 15792 36586
rect 15948 36242 15976 36858
rect 15936 36236 15988 36242
rect 15936 36178 15988 36184
rect 16040 34746 16068 37062
rect 16316 36922 16344 37742
rect 16304 36916 16356 36922
rect 16304 36858 16356 36864
rect 16408 35306 16436 38762
rect 16500 38486 16528 39850
rect 16592 39438 16620 40462
rect 17880 40390 17908 42094
rect 18340 41750 18368 42706
rect 18328 41744 18380 41750
rect 18328 41686 18380 41692
rect 17868 40384 17920 40390
rect 17868 40326 17920 40332
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 16672 39908 16724 39914
rect 16672 39850 16724 39856
rect 16684 39506 16712 39850
rect 16817 39740 17113 39760
rect 16873 39738 16897 39740
rect 16953 39738 16977 39740
rect 17033 39738 17057 39740
rect 16895 39686 16897 39738
rect 16959 39686 16971 39738
rect 17033 39686 17035 39738
rect 16873 39684 16897 39686
rect 16953 39684 16977 39686
rect 17033 39684 17057 39686
rect 16817 39664 17113 39684
rect 18340 39642 18368 39918
rect 18328 39636 18380 39642
rect 18328 39578 18380 39584
rect 16672 39500 16724 39506
rect 16672 39442 16724 39448
rect 16580 39432 16632 39438
rect 16580 39374 16632 39380
rect 16670 38992 16726 39001
rect 16670 38927 16726 38936
rect 16684 38894 16712 38927
rect 16672 38888 16724 38894
rect 16672 38830 16724 38836
rect 16817 38652 17113 38672
rect 16873 38650 16897 38652
rect 16953 38650 16977 38652
rect 17033 38650 17057 38652
rect 16895 38598 16897 38650
rect 16959 38598 16971 38650
rect 17033 38598 17035 38650
rect 16873 38596 16897 38598
rect 16953 38596 16977 38598
rect 17033 38596 17057 38598
rect 16817 38576 17113 38596
rect 16488 38480 16540 38486
rect 16488 38422 16540 38428
rect 16672 37732 16724 37738
rect 16672 37674 16724 37680
rect 16684 37346 16712 37674
rect 16817 37564 17113 37584
rect 16873 37562 16897 37564
rect 16953 37562 16977 37564
rect 17033 37562 17057 37564
rect 16895 37510 16897 37562
rect 16959 37510 16971 37562
rect 17033 37510 17035 37562
rect 16873 37508 16897 37510
rect 16953 37508 16977 37510
rect 17033 37508 17057 37510
rect 16817 37488 17113 37508
rect 16684 37330 16804 37346
rect 16684 37324 16816 37330
rect 16684 37318 16764 37324
rect 16764 37266 16816 37272
rect 16817 36476 17113 36496
rect 16873 36474 16897 36476
rect 16953 36474 16977 36476
rect 17033 36474 17057 36476
rect 16895 36422 16897 36474
rect 16959 36422 16971 36474
rect 17033 36422 17035 36474
rect 16873 36420 16897 36422
rect 16953 36420 16977 36422
rect 17033 36420 17057 36422
rect 16817 36400 17113 36420
rect 17132 36032 17184 36038
rect 17132 35974 17184 35980
rect 16580 35488 16632 35494
rect 16580 35430 16632 35436
rect 16408 35278 16528 35306
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15672 33130 15700 34478
rect 15764 34066 15792 34478
rect 15752 34060 15804 34066
rect 15752 34002 15804 34008
rect 16040 33658 16068 34682
rect 16304 34604 16356 34610
rect 16304 34546 16356 34552
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16028 33652 16080 33658
rect 16028 33594 16080 33600
rect 16316 33454 16344 34546
rect 16408 33998 16436 34546
rect 16396 33992 16448 33998
rect 16396 33934 16448 33940
rect 16500 33810 16528 35278
rect 16408 33782 16528 33810
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 15672 33102 15792 33130
rect 15580 32966 15700 32994
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15580 31482 15608 31758
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15580 29714 15608 30058
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15580 27538 15608 28358
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15580 26246 15608 27270
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15580 25838 15608 26182
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15568 22704 15620 22710
rect 15568 22646 15620 22652
rect 15580 22234 15608 22646
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15580 21010 15608 22170
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20262 15608 20810
rect 15672 20466 15700 32966
rect 15764 23730 15792 33102
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 15856 31278 15884 32846
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16212 32292 16264 32298
rect 16212 32234 16264 32240
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15856 30258 15884 31214
rect 16040 31210 16068 31962
rect 16224 31890 16252 32234
rect 16316 32026 16344 32302
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 16212 31884 16264 31890
rect 16212 31826 16264 31832
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16224 31346 16252 31826
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16028 31204 16080 31210
rect 16028 31146 16080 31152
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15856 28558 15884 30194
rect 15936 30184 15988 30190
rect 15936 30126 15988 30132
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15856 25294 15884 28494
rect 15948 28218 15976 30126
rect 16040 28490 16068 30670
rect 16316 30274 16344 31826
rect 16224 30258 16344 30274
rect 16212 30252 16344 30258
rect 16264 30246 16344 30252
rect 16212 30194 16264 30200
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16028 28484 16080 28490
rect 16028 28426 16080 28432
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 15948 26994 15976 28154
rect 16040 27470 16068 28426
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 16040 27130 16068 27406
rect 16132 27130 16160 28562
rect 16224 28014 16252 30194
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16316 27826 16344 29106
rect 16224 27798 16344 27826
rect 16224 27334 16252 27798
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 16224 26926 16252 27270
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15948 24886 15976 25434
rect 16040 25362 16068 26318
rect 16224 25906 16252 26862
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16120 25764 16172 25770
rect 16120 25706 16172 25712
rect 16028 25356 16080 25362
rect 16028 25298 16080 25304
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15580 19122 15608 20198
rect 15764 19258 15792 21830
rect 15856 21486 15884 24210
rect 16132 23610 16160 25706
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 23730 16252 25638
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16316 24410 16344 25230
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 16132 23582 16252 23610
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15488 19094 15608 19122
rect 15672 19230 15792 19258
rect 15488 18766 15516 19094
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18222 15516 18702
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15488 16658 15516 18158
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15580 16998 15608 17070
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15566 16688 15622 16697
rect 15476 16652 15528 16658
rect 15566 16623 15622 16632
rect 15476 16594 15528 16600
rect 15580 16590 15608 16623
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15396 16102 15516 16130
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15638 15424 15982
rect 15488 15706 15516 16102
rect 15672 16046 15700 19230
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18630 15792 19110
rect 15856 18714 15884 21422
rect 15948 20448 15976 22510
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16132 20942 16160 21966
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16028 20460 16080 20466
rect 15948 20420 16028 20448
rect 16028 20402 16080 20408
rect 16040 19310 16068 20402
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19378 16160 20198
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18902 16068 19246
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 15856 18686 16068 18714
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15764 17882 15792 18158
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 16040 17746 16068 18686
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15856 17134 15884 17682
rect 16040 17338 16068 17682
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 16040 16658 16068 17002
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15764 16538 15792 16594
rect 15764 16510 15884 16538
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15672 15570 15700 15982
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15304 15422 15424 15450
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 13870 15332 14350
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 13682 15332 13806
rect 15396 13802 15424 15422
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15304 13654 15424 13682
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15304 10606 15332 13398
rect 15396 13190 15424 13654
rect 15488 13190 15516 15506
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 15094 15792 15438
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 13938 15608 14758
rect 15764 14618 15792 14894
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 13938 15700 14486
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15764 13326 15792 14554
rect 15856 14414 15884 16510
rect 16132 16250 16160 16594
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16224 16114 16252 23582
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16316 21486 16344 22578
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16316 20806 16344 21422
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16408 20618 16436 33782
rect 16592 33386 16620 35430
rect 16817 35388 17113 35408
rect 16873 35386 16897 35388
rect 16953 35386 16977 35388
rect 17033 35386 17057 35388
rect 16895 35334 16897 35386
rect 16959 35334 16971 35386
rect 17033 35334 17035 35386
rect 16873 35332 16897 35334
rect 16953 35332 16977 35334
rect 17033 35332 17057 35334
rect 16817 35312 17113 35332
rect 17144 35154 17172 35974
rect 18432 35630 18460 46650
rect 18512 46164 18564 46170
rect 18512 46106 18564 46112
rect 18524 40730 18552 46106
rect 18512 40724 18564 40730
rect 18512 40666 18564 40672
rect 19996 38418 20024 46854
rect 20088 46442 20116 49200
rect 20824 47410 20852 49200
rect 20824 47382 21312 47410
rect 21180 47252 21232 47258
rect 21180 47194 21232 47200
rect 20782 46812 21078 46832
rect 20838 46810 20862 46812
rect 20918 46810 20942 46812
rect 20998 46810 21022 46812
rect 20860 46758 20862 46810
rect 20924 46758 20936 46810
rect 20998 46758 21000 46810
rect 20838 46756 20862 46758
rect 20918 46756 20942 46758
rect 20998 46756 21022 46758
rect 20782 46736 21078 46756
rect 20076 46436 20128 46442
rect 20076 46378 20128 46384
rect 20782 45724 21078 45744
rect 20838 45722 20862 45724
rect 20918 45722 20942 45724
rect 20998 45722 21022 45724
rect 20860 45670 20862 45722
rect 20924 45670 20936 45722
rect 20998 45670 21000 45722
rect 20838 45668 20862 45670
rect 20918 45668 20942 45670
rect 20998 45668 21022 45670
rect 20782 45648 21078 45668
rect 20782 44636 21078 44656
rect 20838 44634 20862 44636
rect 20918 44634 20942 44636
rect 20998 44634 21022 44636
rect 20860 44582 20862 44634
rect 20924 44582 20936 44634
rect 20998 44582 21000 44634
rect 20838 44580 20862 44582
rect 20918 44580 20942 44582
rect 20998 44580 21022 44582
rect 20782 44560 21078 44580
rect 20782 43548 21078 43568
rect 20838 43546 20862 43548
rect 20918 43546 20942 43548
rect 20998 43546 21022 43548
rect 20860 43494 20862 43546
rect 20924 43494 20936 43546
rect 20998 43494 21000 43546
rect 20838 43492 20862 43494
rect 20918 43492 20942 43494
rect 20998 43492 21022 43494
rect 20782 43472 21078 43492
rect 20782 42460 21078 42480
rect 20838 42458 20862 42460
rect 20918 42458 20942 42460
rect 20998 42458 21022 42460
rect 20860 42406 20862 42458
rect 20924 42406 20936 42458
rect 20998 42406 21000 42458
rect 20838 42404 20862 42406
rect 20918 42404 20942 42406
rect 20998 42404 21022 42406
rect 20782 42384 21078 42404
rect 21192 41750 21220 47194
rect 21284 42770 21312 47382
rect 21652 47258 21680 49200
rect 22100 49156 22152 49162
rect 22100 49098 22152 49104
rect 21640 47252 21692 47258
rect 21640 47194 21692 47200
rect 21364 46436 21416 46442
rect 21364 46378 21416 46384
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 21180 41744 21232 41750
rect 21180 41686 21232 41692
rect 20782 41372 21078 41392
rect 20838 41370 20862 41372
rect 20918 41370 20942 41372
rect 20998 41370 21022 41372
rect 20860 41318 20862 41370
rect 20924 41318 20936 41370
rect 20998 41318 21000 41370
rect 20838 41316 20862 41318
rect 20918 41316 20942 41318
rect 20998 41316 21022 41318
rect 20782 41296 21078 41316
rect 20782 40284 21078 40304
rect 20838 40282 20862 40284
rect 20918 40282 20942 40284
rect 20998 40282 21022 40284
rect 20860 40230 20862 40282
rect 20924 40230 20936 40282
rect 20998 40230 21000 40282
rect 20838 40228 20862 40230
rect 20918 40228 20942 40230
rect 20998 40228 21022 40230
rect 20782 40208 21078 40228
rect 20782 39196 21078 39216
rect 20838 39194 20862 39196
rect 20918 39194 20942 39196
rect 20998 39194 21022 39196
rect 20860 39142 20862 39194
rect 20924 39142 20936 39194
rect 20998 39142 21000 39194
rect 20838 39140 20862 39142
rect 20918 39140 20942 39142
rect 20998 39140 21022 39142
rect 20782 39120 21078 39140
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 19996 37398 20024 38354
rect 20782 38108 21078 38128
rect 20838 38106 20862 38108
rect 20918 38106 20942 38108
rect 20998 38106 21022 38108
rect 20860 38054 20862 38106
rect 20924 38054 20936 38106
rect 20998 38054 21000 38106
rect 20838 38052 20862 38054
rect 20918 38052 20942 38054
rect 20998 38052 21022 38054
rect 20782 38032 21078 38052
rect 19984 37392 20036 37398
rect 19984 37334 20036 37340
rect 20782 37020 21078 37040
rect 20838 37018 20862 37020
rect 20918 37018 20942 37020
rect 20998 37018 21022 37020
rect 20860 36966 20862 37018
rect 20924 36966 20936 37018
rect 20998 36966 21000 37018
rect 20838 36964 20862 36966
rect 20918 36964 20942 36966
rect 20998 36964 21022 36966
rect 20782 36944 21078 36964
rect 20782 35932 21078 35952
rect 20838 35930 20862 35932
rect 20918 35930 20942 35932
rect 20998 35930 21022 35932
rect 20860 35878 20862 35930
rect 20924 35878 20936 35930
rect 20998 35878 21000 35930
rect 20838 35876 20862 35878
rect 20918 35876 20942 35878
rect 20998 35876 21022 35878
rect 20782 35856 21078 35876
rect 18420 35624 18472 35630
rect 18420 35566 18472 35572
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 16580 33380 16632 33386
rect 16580 33322 16632 33328
rect 16684 32978 16712 35090
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 16817 34300 17113 34320
rect 16873 34298 16897 34300
rect 16953 34298 16977 34300
rect 17033 34298 17057 34300
rect 16895 34246 16897 34298
rect 16959 34246 16971 34298
rect 17033 34246 17035 34298
rect 16873 34244 16897 34246
rect 16953 34244 16977 34246
rect 17033 34244 17057 34246
rect 16817 34224 17113 34244
rect 17236 34066 17264 34886
rect 18432 34134 18460 35566
rect 19616 35556 19668 35562
rect 19616 35498 19668 35504
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18524 34746 18552 35022
rect 18512 34740 18564 34746
rect 18512 34682 18564 34688
rect 19628 34474 19656 35498
rect 21376 35222 21404 46378
rect 22112 39982 22140 49098
rect 22480 46170 22508 49200
rect 23216 49162 23244 49200
rect 23204 49156 23256 49162
rect 23204 49098 23256 49104
rect 24044 46918 24072 49200
rect 24032 46912 24084 46918
rect 24032 46854 24084 46860
rect 24780 46442 24808 49200
rect 25608 46714 25636 49200
rect 25596 46708 25648 46714
rect 25596 46650 25648 46656
rect 24768 46436 24820 46442
rect 24768 46378 24820 46384
rect 22468 46164 22520 46170
rect 22468 46106 22520 46112
rect 22100 39976 22152 39982
rect 22100 39918 22152 39924
rect 21364 35216 21416 35222
rect 21364 35158 21416 35164
rect 20782 34844 21078 34864
rect 20838 34842 20862 34844
rect 20918 34842 20942 34844
rect 20998 34842 21022 34844
rect 20860 34790 20862 34842
rect 20924 34790 20936 34842
rect 20998 34790 21000 34842
rect 20838 34788 20862 34790
rect 20918 34788 20942 34790
rect 20998 34788 21022 34790
rect 20782 34768 21078 34788
rect 21376 34542 21404 35158
rect 21364 34536 21416 34542
rect 21364 34478 21416 34484
rect 19616 34468 19668 34474
rect 19616 34410 19668 34416
rect 18420 34128 18472 34134
rect 18420 34070 18472 34076
rect 17224 34060 17276 34066
rect 17224 34002 17276 34008
rect 16764 33992 16816 33998
rect 16764 33934 16816 33940
rect 16776 33522 16804 33934
rect 20782 33756 21078 33776
rect 20838 33754 20862 33756
rect 20918 33754 20942 33756
rect 20998 33754 21022 33756
rect 20860 33702 20862 33754
rect 20924 33702 20936 33754
rect 20998 33702 21000 33754
rect 20838 33700 20862 33702
rect 20918 33700 20942 33702
rect 20998 33700 21022 33702
rect 20782 33680 21078 33700
rect 16764 33516 16816 33522
rect 16764 33458 16816 33464
rect 16817 33212 17113 33232
rect 16873 33210 16897 33212
rect 16953 33210 16977 33212
rect 17033 33210 17057 33212
rect 16895 33158 16897 33210
rect 16959 33158 16971 33210
rect 17033 33158 17035 33210
rect 16873 33156 16897 33158
rect 16953 33156 16977 33158
rect 17033 33156 17057 33158
rect 16817 33136 17113 33156
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16488 32292 16540 32298
rect 16488 32234 16540 32240
rect 16500 31890 16528 32234
rect 16592 32230 16620 32846
rect 20782 32668 21078 32688
rect 20838 32666 20862 32668
rect 20918 32666 20942 32668
rect 20998 32666 21022 32668
rect 20860 32614 20862 32666
rect 20924 32614 20936 32666
rect 20998 32614 21000 32666
rect 20838 32612 20862 32614
rect 20918 32612 20942 32614
rect 20998 32612 21022 32614
rect 20782 32592 21078 32612
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16488 31884 16540 31890
rect 16488 31826 16540 31832
rect 16592 30802 16620 32166
rect 16817 32124 17113 32144
rect 16873 32122 16897 32124
rect 16953 32122 16977 32124
rect 17033 32122 17057 32124
rect 16895 32070 16897 32122
rect 16959 32070 16971 32122
rect 17033 32070 17035 32122
rect 16873 32068 16897 32070
rect 16953 32068 16977 32070
rect 17033 32068 17057 32070
rect 16817 32048 17113 32068
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17880 31414 17908 31622
rect 20782 31580 21078 31600
rect 20838 31578 20862 31580
rect 20918 31578 20942 31580
rect 20998 31578 21022 31580
rect 20860 31526 20862 31578
rect 20924 31526 20936 31578
rect 20998 31526 21000 31578
rect 20838 31524 20862 31526
rect 20918 31524 20942 31526
rect 20998 31524 21022 31526
rect 20782 31504 21078 31524
rect 17868 31408 17920 31414
rect 17868 31350 17920 31356
rect 16817 31036 17113 31056
rect 16873 31034 16897 31036
rect 16953 31034 16977 31036
rect 17033 31034 17057 31036
rect 16895 30982 16897 31034
rect 16959 30982 16971 31034
rect 17033 30982 17035 31034
rect 16873 30980 16897 30982
rect 16953 30980 16977 30982
rect 17033 30980 17057 30982
rect 16817 30960 17113 30980
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16488 30592 16540 30598
rect 16488 30534 16540 30540
rect 16500 30190 16528 30534
rect 20782 30492 21078 30512
rect 20838 30490 20862 30492
rect 20918 30490 20942 30492
rect 20998 30490 21022 30492
rect 20860 30438 20862 30490
rect 20924 30438 20936 30490
rect 20998 30438 21000 30490
rect 20838 30436 20862 30438
rect 20918 30436 20942 30438
rect 20998 30436 21022 30438
rect 20782 30416 21078 30436
rect 16488 30184 16540 30190
rect 16488 30126 16540 30132
rect 16500 29510 16528 30126
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 16817 29948 17113 29968
rect 16873 29946 16897 29948
rect 16953 29946 16977 29948
rect 17033 29946 17057 29948
rect 16895 29894 16897 29946
rect 16959 29894 16971 29946
rect 17033 29894 17035 29946
rect 16873 29892 16897 29894
rect 16953 29892 16977 29894
rect 17033 29892 17057 29894
rect 16817 29872 17113 29892
rect 16488 29504 16540 29510
rect 16488 29446 16540 29452
rect 16500 29102 16528 29446
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 16500 28014 16528 29038
rect 16817 28860 17113 28880
rect 16873 28858 16897 28860
rect 16953 28858 16977 28860
rect 17033 28858 17057 28860
rect 16895 28806 16897 28858
rect 16959 28806 16971 28858
rect 17033 28806 17035 28858
rect 16873 28804 16897 28806
rect 16953 28804 16977 28806
rect 17033 28804 17057 28806
rect 16817 28784 17113 28804
rect 17604 28762 17632 29990
rect 20782 29404 21078 29424
rect 20838 29402 20862 29404
rect 20918 29402 20942 29404
rect 20998 29402 21022 29404
rect 20860 29350 20862 29402
rect 20924 29350 20936 29402
rect 20998 29350 21000 29402
rect 20838 29348 20862 29350
rect 20918 29348 20942 29350
rect 20998 29348 21022 29350
rect 20782 29328 21078 29348
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16592 28014 16620 28494
rect 20782 28316 21078 28336
rect 20838 28314 20862 28316
rect 20918 28314 20942 28316
rect 20998 28314 21022 28316
rect 20860 28262 20862 28314
rect 20924 28262 20936 28314
rect 20998 28262 21000 28314
rect 20838 28260 20862 28262
rect 20918 28260 20942 28262
rect 20998 28260 21022 28262
rect 20782 28240 21078 28260
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16580 28008 16632 28014
rect 16580 27950 16632 27956
rect 16817 27772 17113 27792
rect 16873 27770 16897 27772
rect 16953 27770 16977 27772
rect 17033 27770 17057 27772
rect 16895 27718 16897 27770
rect 16959 27718 16971 27770
rect 17033 27718 17035 27770
rect 16873 27716 16897 27718
rect 16953 27716 16977 27718
rect 17033 27716 17057 27718
rect 16817 27696 17113 27716
rect 20782 27228 21078 27248
rect 20838 27226 20862 27228
rect 20918 27226 20942 27228
rect 20998 27226 21022 27228
rect 20860 27174 20862 27226
rect 20924 27174 20936 27226
rect 20998 27174 21000 27226
rect 20838 27172 20862 27174
rect 20918 27172 20942 27174
rect 20998 27172 21022 27174
rect 20782 27152 21078 27172
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 16500 26518 16528 26862
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 16817 26684 17113 26704
rect 16873 26682 16897 26684
rect 16953 26682 16977 26684
rect 17033 26682 17057 26684
rect 16895 26630 16897 26682
rect 16959 26630 16971 26682
rect 17033 26630 17035 26682
rect 16873 26628 16897 26630
rect 16953 26628 16977 26630
rect 17033 26628 17057 26630
rect 16817 26608 17113 26628
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16488 24676 16540 24682
rect 16592 24664 16620 25774
rect 16540 24636 16620 24664
rect 16488 24618 16540 24624
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16500 23798 16528 24142
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16500 23322 16528 23598
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16500 22710 16528 23258
rect 16592 23254 16620 24636
rect 16684 24342 16712 26318
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 16817 25596 17113 25616
rect 16873 25594 16897 25596
rect 16953 25594 16977 25596
rect 17033 25594 17057 25596
rect 16895 25542 16897 25594
rect 16959 25542 16971 25594
rect 17033 25542 17035 25594
rect 16873 25540 16897 25542
rect 16953 25540 16977 25542
rect 17033 25540 17057 25542
rect 16817 25520 17113 25540
rect 17972 25430 18000 26182
rect 17960 25424 18012 25430
rect 17960 25366 18012 25372
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 16817 24508 17113 24528
rect 16873 24506 16897 24508
rect 16953 24506 16977 24508
rect 17033 24506 17057 24508
rect 16895 24454 16897 24506
rect 16959 24454 16971 24506
rect 17033 24454 17035 24506
rect 16873 24452 16897 24454
rect 16953 24452 16977 24454
rect 17033 24452 17057 24454
rect 16817 24432 17113 24452
rect 16672 24336 16724 24342
rect 16672 24278 16724 24284
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17144 23662 17172 24210
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16684 22574 16712 23598
rect 16817 23420 17113 23440
rect 16873 23418 16897 23420
rect 16953 23418 16977 23420
rect 17033 23418 17057 23420
rect 16895 23366 16897 23418
rect 16959 23366 16971 23418
rect 17033 23366 17035 23418
rect 16873 23364 16897 23366
rect 16953 23364 16977 23366
rect 17033 23364 17057 23366
rect 16817 23344 17113 23364
rect 17144 23186 17172 23598
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16592 22030 16620 22442
rect 16817 22332 17113 22352
rect 16873 22330 16897 22332
rect 16953 22330 16977 22332
rect 17033 22330 17057 22332
rect 16895 22278 16897 22330
rect 16959 22278 16971 22330
rect 17033 22278 17035 22330
rect 16873 22276 16897 22278
rect 16953 22276 16977 22278
rect 17033 22276 17057 22278
rect 16817 22256 17113 22276
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16500 21690 16528 21966
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16817 21244 17113 21264
rect 16873 21242 16897 21244
rect 16953 21242 16977 21244
rect 17033 21242 17057 21244
rect 16895 21190 16897 21242
rect 16959 21190 16971 21242
rect 17033 21190 17035 21242
rect 16873 21188 16897 21190
rect 16953 21188 16977 21190
rect 17033 21188 17057 21190
rect 16817 21168 17113 21188
rect 16316 20590 16436 20618
rect 16316 19174 16344 20590
rect 17144 20466 17172 22510
rect 17222 21448 17278 21457
rect 17222 21383 17278 21392
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17626 16436 18022
rect 16500 17746 16528 19246
rect 16592 19242 16620 20402
rect 16817 20156 17113 20176
rect 16873 20154 16897 20156
rect 16953 20154 16977 20156
rect 17033 20154 17057 20156
rect 16895 20102 16897 20154
rect 16959 20102 16971 20154
rect 17033 20102 17035 20154
rect 16873 20100 16897 20102
rect 16953 20100 16977 20102
rect 17033 20100 17057 20102
rect 16817 20080 17113 20100
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16684 18834 16712 19654
rect 17144 19378 17172 20402
rect 17236 20330 17264 21383
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16817 19068 17113 19088
rect 16873 19066 16897 19068
rect 16953 19066 16977 19068
rect 17033 19066 17057 19068
rect 16895 19014 16897 19066
rect 16959 19014 16971 19066
rect 17033 19014 17035 19066
rect 16873 19012 16897 19014
rect 16953 19012 16977 19014
rect 17033 19012 17057 19014
rect 16817 18992 17113 19012
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16817 17980 17113 18000
rect 16873 17978 16897 17980
rect 16953 17978 16977 17980
rect 17033 17978 17057 17980
rect 16895 17926 16897 17978
rect 16959 17926 16971 17978
rect 17033 17926 17035 17978
rect 16873 17924 16897 17926
rect 16953 17924 16977 17926
rect 17033 17924 17057 17926
rect 16817 17904 17113 17924
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16592 17626 16620 17682
rect 16408 17598 16620 17626
rect 17144 16998 17172 19178
rect 17512 17202 17540 24890
rect 17592 24676 17644 24682
rect 17592 24618 17644 24624
rect 17604 23526 17632 24618
rect 17972 24342 18000 25366
rect 17960 24336 18012 24342
rect 17960 24278 18012 24284
rect 18064 23662 18092 26386
rect 18156 25974 18184 26726
rect 20782 26140 21078 26160
rect 20838 26138 20862 26140
rect 20918 26138 20942 26140
rect 20998 26138 21022 26140
rect 20860 26086 20862 26138
rect 20924 26086 20936 26138
rect 20998 26086 21000 26138
rect 20838 26084 20862 26086
rect 20918 26084 20942 26086
rect 20998 26084 21022 26086
rect 20782 26064 21078 26084
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 20782 25052 21078 25072
rect 20838 25050 20862 25052
rect 20918 25050 20942 25052
rect 20998 25050 21022 25052
rect 20860 24998 20862 25050
rect 20924 24998 20936 25050
rect 20998 24998 21000 25050
rect 20838 24996 20862 24998
rect 20918 24996 20942 24998
rect 20998 24996 21022 24998
rect 20782 24976 21078 24996
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18052 23656 18104 23662
rect 17958 23624 18014 23633
rect 18052 23598 18104 23604
rect 17958 23559 18014 23568
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17880 23186 17908 23462
rect 17972 23186 18000 23559
rect 18156 23254 18184 24210
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17696 22234 17724 22646
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17604 19922 17632 21490
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17788 19922 17816 20402
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 16817 16892 17113 16912
rect 16873 16890 16897 16892
rect 16953 16890 16977 16892
rect 17033 16890 17057 16892
rect 16895 16838 16897 16890
rect 16959 16838 16971 16890
rect 17033 16838 17035 16890
rect 16873 16836 16897 16838
rect 16953 16836 16977 16838
rect 17033 16836 17057 16838
rect 16817 16816 17113 16836
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16212 16108 16264 16114
rect 16264 16068 16344 16096
rect 16212 16050 16264 16056
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16132 13462 16160 15982
rect 16316 15570 16344 16068
rect 16960 16046 16988 16390
rect 17144 16250 17172 16934
rect 17604 16810 17632 19858
rect 17788 18986 17816 19858
rect 17880 19310 17908 23122
rect 18248 22982 18276 24550
rect 18420 24336 18472 24342
rect 18420 24278 18472 24284
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18340 22778 18368 23666
rect 18432 23594 18460 24278
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18524 23662 18552 23802
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18248 22098 18276 22510
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 18052 21412 18104 21418
rect 18052 21354 18104 21360
rect 18064 21010 18092 21354
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 18248 20942 18276 22034
rect 18326 21584 18382 21593
rect 18326 21519 18382 21528
rect 18340 21418 18368 21519
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18236 20936 18288 20942
rect 18288 20884 18368 20890
rect 18236 20878 18368 20884
rect 18248 20862 18368 20878
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17788 18958 17908 18986
rect 17880 18834 17908 18958
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17880 18630 17908 18770
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18154 17908 18566
rect 17972 18222 18000 19858
rect 18248 19514 18276 20742
rect 18340 20602 18368 20862
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18432 20466 18460 23530
rect 18616 22642 18644 24142
rect 19168 24138 19196 24686
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 20782 23964 21078 23984
rect 20838 23962 20862 23964
rect 20918 23962 20942 23964
rect 20998 23962 21022 23964
rect 20860 23910 20862 23962
rect 20924 23910 20936 23962
rect 20998 23910 21000 23962
rect 20838 23908 20862 23910
rect 20918 23908 20942 23910
rect 20998 23908 21022 23910
rect 20782 23888 21078 23908
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18708 22098 18736 23122
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19260 22778 19288 23054
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 19168 21486 19196 22442
rect 19260 21554 19288 22714
rect 19444 22710 19472 22918
rect 20782 22876 21078 22896
rect 20838 22874 20862 22876
rect 20918 22874 20942 22876
rect 20998 22874 21022 22876
rect 20860 22822 20862 22874
rect 20924 22822 20936 22874
rect 20998 22822 21000 22874
rect 20838 22820 20862 22822
rect 20918 22820 20942 22822
rect 20998 22820 21022 22822
rect 20782 22800 21078 22820
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 22098 19564 22374
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 20782 21788 21078 21808
rect 20838 21786 20862 21788
rect 20918 21786 20942 21788
rect 20998 21786 21022 21788
rect 20860 21734 20862 21786
rect 20924 21734 20936 21786
rect 20998 21734 21000 21786
rect 20838 21732 20862 21734
rect 20918 21732 20942 21734
rect 20998 21732 21022 21734
rect 20782 21712 21078 21732
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19076 21010 19104 21422
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18248 18970 18276 19314
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17604 16782 17724 16810
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 16224 13394 16252 15438
rect 16592 14958 16620 15914
rect 16817 15804 17113 15824
rect 16873 15802 16897 15804
rect 16953 15802 16977 15804
rect 17033 15802 17057 15804
rect 16895 15750 16897 15802
rect 16959 15750 16971 15802
rect 17033 15750 17035 15802
rect 16873 15748 16897 15750
rect 16953 15748 16977 15750
rect 17033 15748 17057 15750
rect 16817 15728 17113 15748
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 6458 15240 10066
rect 15488 9450 15516 13126
rect 15672 12850 15700 13126
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 10810 15608 11290
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 16040 10690 16068 10950
rect 16040 10662 16160 10690
rect 16132 10606 16160 10662
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16040 10266 16068 10542
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15290 8936 15346 8945
rect 15290 8871 15346 8880
rect 15304 7954 15332 8871
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 16132 6798 16160 10542
rect 16224 10062 16252 13330
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12782 16344 13194
rect 16500 12918 16528 13398
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16684 12782 16712 15506
rect 17512 15434 17540 16050
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 16817 14716 17113 14736
rect 16873 14714 16897 14716
rect 16953 14714 16977 14716
rect 17033 14714 17057 14716
rect 16895 14662 16897 14714
rect 16959 14662 16971 14714
rect 17033 14662 17035 14714
rect 16873 14660 16897 14662
rect 16953 14660 16977 14662
rect 17033 14660 17057 14662
rect 16817 14640 17113 14660
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 13870 16896 14418
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16817 13628 17113 13648
rect 16873 13626 16897 13628
rect 16953 13626 16977 13628
rect 17033 13626 17057 13628
rect 16895 13574 16897 13626
rect 16959 13574 16971 13626
rect 17033 13574 17035 13626
rect 16873 13572 16897 13574
rect 16953 13572 16977 13574
rect 17033 13572 17057 13574
rect 16817 13552 17113 13572
rect 17144 13462 17172 14350
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 16684 12322 16712 12718
rect 16817 12540 17113 12560
rect 16873 12538 16897 12540
rect 16953 12538 16977 12540
rect 17033 12538 17057 12540
rect 16895 12486 16897 12538
rect 16959 12486 16971 12538
rect 17033 12486 17035 12538
rect 16873 12484 16897 12486
rect 16953 12484 16977 12486
rect 17033 12484 17057 12486
rect 16817 12464 17113 12484
rect 16684 12294 16804 12322
rect 17144 12306 17172 12718
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16592 11694 16620 11766
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10198 16344 10950
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16408 10606 16436 10746
rect 16500 10606 16528 11494
rect 16684 11370 16712 12174
rect 16776 11608 16804 12294
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11762 17172 12242
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16856 11620 16908 11626
rect 16776 11580 16856 11608
rect 16856 11562 16908 11568
rect 16817 11452 17113 11472
rect 16873 11450 16897 11452
rect 16953 11450 16977 11452
rect 17033 11450 17057 11452
rect 16895 11398 16897 11450
rect 16959 11398 16971 11450
rect 17033 11398 17035 11450
rect 16873 11396 16897 11398
rect 16953 11396 16977 11398
rect 17033 11396 17057 11398
rect 16817 11376 17113 11396
rect 16592 11342 16712 11370
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10198 16528 10542
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9382 16344 9522
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8022 16344 8910
rect 16408 8838 16436 9998
rect 16500 9353 16528 9998
rect 16592 9382 16620 11342
rect 17144 11286 17172 11698
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16684 10130 16712 10746
rect 16817 10364 17113 10384
rect 16873 10362 16897 10364
rect 16953 10362 16977 10364
rect 17033 10362 17057 10364
rect 16895 10310 16897 10362
rect 16959 10310 16971 10362
rect 17033 10310 17035 10362
rect 16873 10308 16897 10310
rect 16953 10308 16977 10310
rect 17033 10308 17057 10310
rect 16817 10288 17113 10308
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 17236 10062 17264 11766
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17236 9518 17264 9998
rect 17328 9994 17356 11834
rect 17512 11626 17540 15370
rect 17604 15366 17632 16186
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17604 12170 17632 15302
rect 17696 13394 17724 16782
rect 17972 15706 18000 18158
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 14958 18000 15642
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17880 14006 17908 14214
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 12238 17724 13330
rect 17880 12306 17908 13806
rect 17972 13394 18000 14214
rect 18064 13462 18092 14758
rect 18156 14278 18184 15438
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17604 11830 17632 12106
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17604 10810 17632 11766
rect 17880 11694 17908 12242
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11354 17908 11630
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17972 10198 18000 12106
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 11218 18092 12038
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18248 10606 18276 17070
rect 18340 12714 18368 19110
rect 18616 18290 18644 19858
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16114 18460 16390
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18432 15502 18460 16050
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18524 13530 18552 16934
rect 18708 16046 18736 20198
rect 19168 19922 19196 21422
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20180 21146 20208 21286
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20782 20700 21078 20720
rect 20838 20698 20862 20700
rect 20918 20698 20942 20700
rect 20998 20698 21022 20700
rect 20860 20646 20862 20698
rect 20924 20646 20936 20698
rect 20998 20646 21000 20698
rect 20838 20644 20862 20646
rect 20918 20644 20942 20646
rect 20998 20644 21022 20646
rect 20782 20624 21078 20644
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 20782 19612 21078 19632
rect 20838 19610 20862 19612
rect 20918 19610 20942 19612
rect 20998 19610 21022 19612
rect 20860 19558 20862 19610
rect 20924 19558 20936 19610
rect 20998 19558 21000 19610
rect 20838 19556 20862 19558
rect 20918 19556 20942 19558
rect 20998 19556 21022 19558
rect 20782 19536 21078 19556
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19536 18426 19564 18634
rect 20782 18524 21078 18544
rect 20838 18522 20862 18524
rect 20918 18522 20942 18524
rect 20998 18522 21022 18524
rect 20860 18470 20862 18522
rect 20924 18470 20936 18522
rect 20998 18470 21000 18522
rect 20838 18468 20862 18470
rect 20918 18468 20942 18470
rect 20998 18468 21022 18470
rect 20782 18448 21078 18468
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 20782 17436 21078 17456
rect 20838 17434 20862 17436
rect 20918 17434 20942 17436
rect 20998 17434 21022 17436
rect 20860 17382 20862 17434
rect 20924 17382 20936 17434
rect 20998 17382 21000 17434
rect 20838 17380 20862 17382
rect 20918 17380 20942 17382
rect 20998 17380 21022 17382
rect 20782 17360 21078 17380
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19076 16794 19104 17138
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16250 19288 16594
rect 20782 16348 21078 16368
rect 20838 16346 20862 16348
rect 20918 16346 20942 16348
rect 20998 16346 21022 16348
rect 20860 16294 20862 16346
rect 20924 16294 20936 16346
rect 20998 16294 21000 16346
rect 20838 16292 20862 16294
rect 20918 16292 20942 16294
rect 20998 16292 21022 16294
rect 20782 16272 21078 16292
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 20782 15260 21078 15280
rect 20838 15258 20862 15260
rect 20918 15258 20942 15260
rect 20998 15258 21022 15260
rect 20860 15206 20862 15258
rect 20924 15206 20936 15258
rect 20998 15206 21000 15258
rect 20838 15204 20862 15206
rect 20918 15204 20942 15206
rect 20998 15204 21022 15206
rect 20782 15184 21078 15204
rect 20782 14172 21078 14192
rect 20838 14170 20862 14172
rect 20918 14170 20942 14172
rect 20998 14170 21022 14172
rect 20860 14118 20862 14170
rect 20924 14118 20936 14170
rect 20998 14118 21000 14170
rect 20838 14116 20862 14118
rect 20918 14116 20942 14118
rect 20998 14116 21022 14118
rect 20782 14096 21078 14116
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 16580 9376 16632 9382
rect 16486 9344 16542 9353
rect 16580 9318 16632 9324
rect 16486 9279 16542 9288
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16592 7886 16620 9318
rect 16817 9276 17113 9296
rect 16873 9274 16897 9276
rect 16953 9274 16977 9276
rect 17033 9274 17057 9276
rect 16895 9222 16897 9274
rect 16959 9222 16971 9274
rect 17033 9222 17035 9274
rect 16873 9220 16897 9222
rect 16953 9220 16977 9222
rect 17033 9220 17057 9222
rect 16817 9200 17113 9220
rect 17236 8974 17264 9454
rect 17328 9110 17356 9930
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17498 9072 17554 9081
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 8566 17264 8910
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16817 8188 17113 8208
rect 16873 8186 16897 8188
rect 16953 8186 16977 8188
rect 17033 8186 17057 8188
rect 16895 8134 16897 8186
rect 16959 8134 16971 8186
rect 17033 8134 17035 8186
rect 16873 8132 16897 8134
rect 16953 8132 16977 8134
rect 17033 8132 17057 8134
rect 16817 8112 17113 8132
rect 17236 7954 17264 8502
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 7478 16896 7754
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 17328 7274 17356 9046
rect 17498 9007 17554 9016
rect 17512 8906 17540 9007
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17972 8430 18000 10134
rect 18248 9994 18276 10542
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9722 18184 9862
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18234 9480 18290 9489
rect 18156 9042 18184 9454
rect 18234 9415 18236 9424
rect 18288 9415 18290 9424
rect 18236 9386 18288 9392
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 8022 18184 8230
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18340 7954 18368 12378
rect 18984 12306 19012 13330
rect 20782 13084 21078 13104
rect 20838 13082 20862 13084
rect 20918 13082 20942 13084
rect 20998 13082 21022 13084
rect 20860 13030 20862 13082
rect 20924 13030 20936 13082
rect 20998 13030 21000 13082
rect 20838 13028 20862 13030
rect 20918 13028 20942 13030
rect 20998 13028 21022 13030
rect 20782 13008 21078 13028
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11898 19012 12242
rect 20782 11996 21078 12016
rect 20838 11994 20862 11996
rect 20918 11994 20942 11996
rect 20998 11994 21022 11996
rect 20860 11942 20862 11994
rect 20924 11942 20936 11994
rect 20998 11942 21000 11994
rect 20838 11940 20862 11942
rect 20918 11940 20942 11942
rect 20998 11940 21022 11942
rect 20782 11920 21078 11940
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10606 18460 10950
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18984 10130 19012 11562
rect 20782 10908 21078 10928
rect 20838 10906 20862 10908
rect 20918 10906 20942 10908
rect 20998 10906 21022 10908
rect 20860 10854 20862 10906
rect 20924 10854 20936 10906
rect 20998 10854 21000 10906
rect 20838 10852 20862 10854
rect 20918 10852 20942 10854
rect 20998 10852 21022 10854
rect 20782 10832 21078 10852
rect 19154 10704 19210 10713
rect 19154 10639 19210 10648
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 17512 7342 17540 7890
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7546 18460 7686
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 16592 6798 16620 7142
rect 16817 7100 17113 7120
rect 16873 7098 16897 7100
rect 16953 7098 16977 7100
rect 17033 7098 17057 7100
rect 16895 7046 16897 7098
rect 16959 7046 16971 7098
rect 17033 7046 17035 7098
rect 16873 7044 16897 7046
rect 16953 7044 16977 7046
rect 17033 7044 17057 7046
rect 16817 7024 17113 7044
rect 17144 6934 17172 7142
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17328 6882 17356 7210
rect 17512 7002 17540 7278
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17328 6866 17448 6882
rect 17328 6860 17460 6866
rect 17328 6854 17408 6860
rect 17408 6802 17460 6808
rect 18984 6798 19012 10066
rect 19168 8634 19196 10639
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 10033 20944 10066
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20782 9820 21078 9840
rect 20838 9818 20862 9820
rect 20918 9818 20942 9820
rect 20998 9818 21022 9820
rect 20860 9766 20862 9818
rect 20924 9766 20936 9818
rect 20998 9766 21000 9818
rect 20838 9764 20862 9766
rect 20918 9764 20942 9766
rect 20998 9764 21022 9766
rect 20782 9744 21078 9764
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 20180 8498 20208 9318
rect 20782 8732 21078 8752
rect 20838 8730 20862 8732
rect 20918 8730 20942 8732
rect 20998 8730 21022 8732
rect 20860 8678 20862 8730
rect 20924 8678 20936 8730
rect 20998 8678 21000 8730
rect 20838 8676 20862 8678
rect 20918 8676 20942 8678
rect 20998 8676 21022 8678
rect 20782 8656 21078 8676
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19076 7410 19104 8366
rect 21192 8362 21220 9862
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 20782 7644 21078 7664
rect 20838 7642 20862 7644
rect 20918 7642 20942 7644
rect 20998 7642 21022 7644
rect 20860 7590 20862 7642
rect 20924 7590 20936 7642
rect 20998 7590 21000 7642
rect 20838 7588 20862 7590
rect 20918 7588 20942 7590
rect 20998 7588 21022 7590
rect 20782 7568 21078 7588
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15396 6322 15424 6598
rect 16592 6458 16620 6734
rect 20782 6556 21078 6576
rect 20838 6554 20862 6556
rect 20918 6554 20942 6556
rect 20998 6554 21022 6556
rect 20860 6502 20862 6554
rect 20924 6502 20936 6554
rect 20998 6502 21000 6554
rect 20838 6500 20862 6502
rect 20918 6500 20942 6502
rect 20998 6500 21022 6502
rect 20782 6480 21078 6500
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14016 3454 14136 3482
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 2514 13952 2790
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14016 800 14044 3454
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14292 2106 14320 2246
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14384 800 14412 4762
rect 15120 4146 15148 6190
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 15396 5778 15424 6054
rect 16817 6012 17113 6032
rect 16873 6010 16897 6012
rect 16953 6010 16977 6012
rect 17033 6010 17057 6012
rect 16895 5958 16897 6010
rect 16959 5958 16971 6010
rect 17033 5958 17035 6010
rect 16873 5956 16897 5958
rect 16953 5956 16977 5958
rect 17033 5956 17057 5958
rect 16817 5936 17113 5956
rect 18156 5914 18184 6054
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15212 4826 15240 5714
rect 20782 5468 21078 5488
rect 20838 5466 20862 5468
rect 20918 5466 20942 5468
rect 20998 5466 21022 5468
rect 20860 5414 20862 5466
rect 20924 5414 20936 5466
rect 20998 5414 21000 5466
rect 20838 5412 20862 5414
rect 20918 5412 20942 5414
rect 20998 5412 21022 5414
rect 20782 5392 21078 5412
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 16817 4924 17113 4944
rect 16873 4922 16897 4924
rect 16953 4922 16977 4924
rect 17033 4922 17057 4924
rect 16895 4870 16897 4922
rect 16959 4870 16971 4922
rect 17033 4870 17035 4922
rect 16873 4868 16897 4870
rect 16953 4868 16977 4870
rect 17033 4868 17057 4870
rect 16817 4848 17113 4868
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14568 3602 14596 4082
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14660 2378 14688 3062
rect 14844 3058 14872 4082
rect 16040 4078 16068 4762
rect 18616 4282 18644 5034
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 20782 4380 21078 4400
rect 20838 4378 20862 4380
rect 20918 4378 20942 4380
rect 20998 4378 21022 4380
rect 20860 4326 20862 4378
rect 20924 4326 20936 4378
rect 20998 4326 21000 4378
rect 20838 4324 20862 4326
rect 20918 4324 20942 4326
rect 20998 4324 21022 4326
rect 20782 4304 21078 4324
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 14936 3126 14964 4014
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 15028 2650 15056 3946
rect 22204 3942 22232 4082
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 18512 3936 18564 3942
rect 22192 3936 22244 3942
rect 18564 3896 18644 3924
rect 18512 3878 18564 3884
rect 16132 3670 16160 3878
rect 16817 3836 17113 3856
rect 16873 3834 16897 3836
rect 16953 3834 16977 3836
rect 17033 3834 17057 3836
rect 16895 3782 16897 3834
rect 16959 3782 16971 3834
rect 17033 3782 17035 3834
rect 16873 3780 16897 3782
rect 16953 3780 16977 3782
rect 17033 3780 17057 3782
rect 16817 3760 17113 3780
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15120 2446 15148 2994
rect 15304 2854 15332 3538
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15396 3194 15424 3334
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15396 2514 15424 2858
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14660 800 14688 2314
rect 15120 1714 15148 2382
rect 15028 1686 15148 1714
rect 15028 800 15056 1686
rect 15396 800 15424 2450
rect 15764 800 15792 2790
rect 16132 800 16160 3334
rect 16500 800 16528 3470
rect 16684 1442 16712 3538
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 16817 2748 17113 2768
rect 16873 2746 16897 2748
rect 16953 2746 16977 2748
rect 17033 2746 17057 2748
rect 16895 2694 16897 2746
rect 16959 2694 16971 2746
rect 17033 2694 17035 2746
rect 16873 2692 16897 2694
rect 16953 2692 16977 2694
rect 17033 2692 17057 2694
rect 16817 2672 17113 2692
rect 16684 1414 16896 1442
rect 16868 800 16896 1414
rect 17236 800 17264 3402
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17328 2446 17356 3334
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17512 800 17540 3334
rect 17880 800 17908 3402
rect 18248 800 18276 3538
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18524 1442 18552 3470
rect 18616 2650 18644 3896
rect 22192 3878 22244 3884
rect 22100 3528 22152 3534
rect 22152 3488 22232 3516
rect 22100 3470 22152 3476
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18708 2582 18736 3334
rect 20782 3292 21078 3312
rect 20838 3290 20862 3292
rect 20918 3290 20942 3292
rect 20998 3290 21022 3292
rect 20860 3238 20862 3290
rect 20924 3238 20936 3290
rect 20998 3238 21000 3290
rect 20838 3236 20862 3238
rect 20918 3236 20942 3238
rect 20998 3236 21022 3238
rect 20782 3216 21078 3236
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 2038 18644 2246
rect 18604 2032 18656 2038
rect 18604 1974 18656 1980
rect 18524 1414 18644 1442
rect 18616 800 18644 1414
rect 18984 800 19012 3130
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 800 19380 2926
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19628 898 19656 2858
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 2514 19748 2790
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19628 870 19748 898
rect 19720 800 19748 870
rect 20088 800 20116 3062
rect 20364 800 20392 3062
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20732 2292 20760 2994
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21180 2916 21232 2922
rect 21180 2858 21232 2864
rect 20640 2264 20760 2292
rect 20640 1986 20668 2264
rect 20782 2204 21078 2224
rect 20838 2202 20862 2204
rect 20918 2202 20942 2204
rect 20998 2202 21022 2204
rect 20860 2150 20862 2202
rect 20924 2150 20936 2202
rect 20998 2150 21000 2202
rect 20838 2148 20862 2150
rect 20918 2148 20942 2150
rect 20998 2148 21022 2150
rect 20782 2128 21078 2148
rect 20640 1958 20760 1986
rect 20732 800 20760 1958
rect 21192 1170 21220 2858
rect 21100 1142 21220 1170
rect 21100 800 21128 1142
rect 21468 800 21496 2926
rect 21836 800 21864 3402
rect 22204 800 22232 3488
rect 22296 3194 22324 4150
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22388 3738 22416 4082
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22388 2582 22416 2858
rect 22376 2576 22428 2582
rect 22376 2518 22428 2524
rect 22572 800 22600 3606
rect 22928 3392 22980 3398
rect 22928 3334 22980 3340
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22756 2446 22784 2790
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22940 800 22968 3334
rect 23032 2650 23060 3878
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23308 2258 23336 4422
rect 23400 4010 23428 4422
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23400 2514 23428 2790
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23216 2230 23336 2258
rect 23216 800 23244 2230
rect 23584 800 23612 4558
rect 23952 800 23980 4626
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 24320 800 24348 4490
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24688 800 24716 2926
rect 25412 2916 25464 2922
rect 25412 2858 25464 2864
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 25056 800 25084 2246
rect 25424 800 25452 2858
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 800 25820 2790
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
<< via2 >>
rect 3054 47232 3110 47288
rect 3330 41656 3386 41712
rect 2410 38956 2466 38992
rect 2410 38936 2412 38956
rect 2412 38936 2464 38956
rect 2464 38936 2466 38956
rect 2962 38936 3018 38992
rect 4921 46810 4977 46812
rect 5001 46810 5057 46812
rect 5081 46810 5137 46812
rect 5161 46810 5217 46812
rect 4921 46758 4947 46810
rect 4947 46758 4977 46810
rect 5001 46758 5011 46810
rect 5011 46758 5057 46810
rect 5081 46758 5127 46810
rect 5127 46758 5137 46810
rect 5161 46758 5191 46810
rect 5191 46758 5217 46810
rect 4921 46756 4977 46758
rect 5001 46756 5057 46758
rect 5081 46756 5137 46758
rect 5161 46756 5217 46758
rect 3330 36080 3386 36136
rect 1674 22516 1676 22536
rect 1676 22516 1728 22536
rect 1728 22516 1730 22536
rect 1674 22480 1730 22516
rect 1582 19352 1638 19408
rect 3146 31320 3202 31376
rect 2594 26444 2650 26480
rect 2594 26424 2596 26444
rect 2596 26424 2648 26444
rect 2648 26424 2650 26444
rect 3514 30504 3570 30560
rect 3790 26460 3792 26480
rect 3792 26460 3844 26480
rect 3844 26460 3846 26480
rect 3790 26424 3846 26460
rect 4921 45722 4977 45724
rect 5001 45722 5057 45724
rect 5081 45722 5137 45724
rect 5161 45722 5217 45724
rect 4921 45670 4947 45722
rect 4947 45670 4977 45722
rect 5001 45670 5011 45722
rect 5011 45670 5057 45722
rect 5081 45670 5127 45722
rect 5127 45670 5137 45722
rect 5161 45670 5191 45722
rect 5191 45670 5217 45722
rect 4921 45668 4977 45670
rect 5001 45668 5057 45670
rect 5081 45668 5137 45670
rect 5161 45668 5217 45670
rect 4921 44634 4977 44636
rect 5001 44634 5057 44636
rect 5081 44634 5137 44636
rect 5161 44634 5217 44636
rect 4921 44582 4947 44634
rect 4947 44582 4977 44634
rect 5001 44582 5011 44634
rect 5011 44582 5057 44634
rect 5081 44582 5127 44634
rect 5127 44582 5137 44634
rect 5161 44582 5191 44634
rect 5191 44582 5217 44634
rect 4921 44580 4977 44582
rect 5001 44580 5057 44582
rect 5081 44580 5137 44582
rect 5161 44580 5217 44582
rect 4921 43546 4977 43548
rect 5001 43546 5057 43548
rect 5081 43546 5137 43548
rect 5161 43546 5217 43548
rect 4921 43494 4947 43546
rect 4947 43494 4977 43546
rect 5001 43494 5011 43546
rect 5011 43494 5057 43546
rect 5081 43494 5127 43546
rect 5127 43494 5137 43546
rect 5161 43494 5191 43546
rect 5191 43494 5217 43546
rect 4921 43492 4977 43494
rect 5001 43492 5057 43494
rect 5081 43492 5137 43494
rect 5161 43492 5217 43494
rect 4921 42458 4977 42460
rect 5001 42458 5057 42460
rect 5081 42458 5137 42460
rect 5161 42458 5217 42460
rect 4921 42406 4947 42458
rect 4947 42406 4977 42458
rect 5001 42406 5011 42458
rect 5011 42406 5057 42458
rect 5081 42406 5127 42458
rect 5127 42406 5137 42458
rect 5161 42406 5191 42458
rect 5191 42406 5217 42458
rect 4921 42404 4977 42406
rect 5001 42404 5057 42406
rect 5081 42404 5137 42406
rect 5161 42404 5217 42406
rect 4921 41370 4977 41372
rect 5001 41370 5057 41372
rect 5081 41370 5137 41372
rect 5161 41370 5217 41372
rect 4921 41318 4947 41370
rect 4947 41318 4977 41370
rect 5001 41318 5011 41370
rect 5011 41318 5057 41370
rect 5081 41318 5127 41370
rect 5127 41318 5137 41370
rect 5161 41318 5191 41370
rect 5191 41318 5217 41370
rect 4921 41316 4977 41318
rect 5001 41316 5057 41318
rect 5081 41316 5137 41318
rect 5161 41316 5217 41318
rect 4921 40282 4977 40284
rect 5001 40282 5057 40284
rect 5081 40282 5137 40284
rect 5161 40282 5217 40284
rect 4921 40230 4947 40282
rect 4947 40230 4977 40282
rect 5001 40230 5011 40282
rect 5011 40230 5057 40282
rect 5081 40230 5127 40282
rect 5127 40230 5137 40282
rect 5161 40230 5191 40282
rect 5191 40230 5217 40282
rect 4921 40228 4977 40230
rect 5001 40228 5057 40230
rect 5081 40228 5137 40230
rect 5161 40228 5217 40230
rect 4158 28600 4214 28656
rect 3422 19352 3478 19408
rect 2042 9988 2098 10024
rect 2042 9968 2044 9988
rect 2044 9968 2096 9988
rect 2096 9968 2098 9988
rect 2410 2760 2466 2816
rect 2962 4936 3018 4992
rect 4066 24928 4122 24984
rect 4921 39194 4977 39196
rect 5001 39194 5057 39196
rect 5081 39194 5137 39196
rect 5161 39194 5217 39196
rect 4921 39142 4947 39194
rect 4947 39142 4977 39194
rect 5001 39142 5011 39194
rect 5011 39142 5057 39194
rect 5081 39142 5127 39194
rect 5127 39142 5137 39194
rect 5161 39142 5191 39194
rect 5191 39142 5217 39194
rect 4921 39140 4977 39142
rect 5001 39140 5057 39142
rect 5081 39140 5137 39142
rect 5161 39140 5217 39142
rect 4921 38106 4977 38108
rect 5001 38106 5057 38108
rect 5081 38106 5137 38108
rect 5161 38106 5217 38108
rect 4921 38054 4947 38106
rect 4947 38054 4977 38106
rect 5001 38054 5011 38106
rect 5011 38054 5057 38106
rect 5081 38054 5127 38106
rect 5127 38054 5137 38106
rect 5161 38054 5191 38106
rect 5191 38054 5217 38106
rect 4921 38052 4977 38054
rect 5001 38052 5057 38054
rect 5081 38052 5137 38054
rect 5161 38052 5217 38054
rect 4921 37018 4977 37020
rect 5001 37018 5057 37020
rect 5081 37018 5137 37020
rect 5161 37018 5217 37020
rect 4921 36966 4947 37018
rect 4947 36966 4977 37018
rect 5001 36966 5011 37018
rect 5011 36966 5057 37018
rect 5081 36966 5127 37018
rect 5127 36966 5137 37018
rect 5161 36966 5191 37018
rect 5191 36966 5217 37018
rect 4921 36964 4977 36966
rect 5001 36964 5057 36966
rect 5081 36964 5137 36966
rect 5161 36964 5217 36966
rect 4921 35930 4977 35932
rect 5001 35930 5057 35932
rect 5081 35930 5137 35932
rect 5161 35930 5217 35932
rect 4921 35878 4947 35930
rect 4947 35878 4977 35930
rect 5001 35878 5011 35930
rect 5011 35878 5057 35930
rect 5081 35878 5127 35930
rect 5127 35878 5137 35930
rect 5161 35878 5191 35930
rect 5191 35878 5217 35930
rect 4921 35876 4977 35878
rect 5001 35876 5057 35878
rect 5081 35876 5137 35878
rect 5161 35876 5217 35878
rect 4921 34842 4977 34844
rect 5001 34842 5057 34844
rect 5081 34842 5137 34844
rect 5161 34842 5217 34844
rect 4921 34790 4947 34842
rect 4947 34790 4977 34842
rect 5001 34790 5011 34842
rect 5011 34790 5057 34842
rect 5081 34790 5127 34842
rect 5127 34790 5137 34842
rect 5161 34790 5191 34842
rect 5191 34790 5217 34842
rect 4921 34788 4977 34790
rect 5001 34788 5057 34790
rect 5081 34788 5137 34790
rect 5161 34788 5217 34790
rect 4921 33754 4977 33756
rect 5001 33754 5057 33756
rect 5081 33754 5137 33756
rect 5161 33754 5217 33756
rect 4921 33702 4947 33754
rect 4947 33702 4977 33754
rect 5001 33702 5011 33754
rect 5011 33702 5057 33754
rect 5081 33702 5127 33754
rect 5127 33702 5137 33754
rect 5161 33702 5191 33754
rect 5191 33702 5217 33754
rect 4921 33700 4977 33702
rect 5001 33700 5057 33702
rect 5081 33700 5137 33702
rect 5161 33700 5217 33702
rect 4526 28328 4582 28384
rect 4921 32666 4977 32668
rect 5001 32666 5057 32668
rect 5081 32666 5137 32668
rect 5161 32666 5217 32668
rect 4921 32614 4947 32666
rect 4947 32614 4977 32666
rect 5001 32614 5011 32666
rect 5011 32614 5057 32666
rect 5081 32614 5127 32666
rect 5127 32614 5137 32666
rect 5161 32614 5191 32666
rect 5191 32614 5217 32666
rect 4921 32612 4977 32614
rect 5001 32612 5057 32614
rect 5081 32612 5137 32614
rect 5161 32612 5217 32614
rect 5354 34176 5410 34232
rect 4921 31578 4977 31580
rect 5001 31578 5057 31580
rect 5081 31578 5137 31580
rect 5161 31578 5217 31580
rect 4921 31526 4947 31578
rect 4947 31526 4977 31578
rect 5001 31526 5011 31578
rect 5011 31526 5057 31578
rect 5081 31526 5127 31578
rect 5127 31526 5137 31578
rect 5161 31526 5191 31578
rect 5191 31526 5217 31578
rect 4921 31524 4977 31526
rect 5001 31524 5057 31526
rect 5081 31524 5137 31526
rect 5161 31524 5217 31526
rect 4894 31320 4950 31376
rect 8886 47354 8942 47356
rect 8966 47354 9022 47356
rect 9046 47354 9102 47356
rect 9126 47354 9182 47356
rect 8886 47302 8912 47354
rect 8912 47302 8942 47354
rect 8966 47302 8976 47354
rect 8976 47302 9022 47354
rect 9046 47302 9092 47354
rect 9092 47302 9102 47354
rect 9126 47302 9156 47354
rect 9156 47302 9182 47354
rect 8886 47300 8942 47302
rect 8966 47300 9022 47302
rect 9046 47300 9102 47302
rect 9126 47300 9182 47302
rect 5446 31592 5502 31648
rect 4921 30490 4977 30492
rect 5001 30490 5057 30492
rect 5081 30490 5137 30492
rect 5161 30490 5217 30492
rect 4921 30438 4947 30490
rect 4947 30438 4977 30490
rect 5001 30438 5011 30490
rect 5011 30438 5057 30490
rect 5081 30438 5127 30490
rect 5127 30438 5137 30490
rect 5161 30438 5191 30490
rect 5191 30438 5217 30490
rect 4921 30436 4977 30438
rect 5001 30436 5057 30438
rect 5081 30436 5137 30438
rect 5161 30436 5217 30438
rect 4921 29402 4977 29404
rect 5001 29402 5057 29404
rect 5081 29402 5137 29404
rect 5161 29402 5217 29404
rect 4921 29350 4947 29402
rect 4947 29350 4977 29402
rect 5001 29350 5011 29402
rect 5011 29350 5057 29402
rect 5081 29350 5127 29402
rect 5127 29350 5137 29402
rect 5161 29350 5191 29402
rect 5191 29350 5217 29402
rect 4921 29348 4977 29350
rect 5001 29348 5057 29350
rect 5081 29348 5137 29350
rect 5161 29348 5217 29350
rect 4802 28600 4858 28656
rect 4802 28500 4804 28520
rect 4804 28500 4856 28520
rect 4856 28500 4858 28520
rect 4802 28464 4858 28500
rect 5078 28464 5134 28520
rect 4250 21528 4306 21584
rect 4342 20848 4398 20904
rect 4066 8200 4122 8256
rect 4921 28314 4977 28316
rect 5001 28314 5057 28316
rect 5081 28314 5137 28316
rect 5161 28314 5217 28316
rect 4921 28262 4947 28314
rect 4947 28262 4977 28314
rect 5001 28262 5011 28314
rect 5011 28262 5057 28314
rect 5081 28262 5127 28314
rect 5127 28262 5137 28314
rect 5161 28262 5191 28314
rect 5191 28262 5217 28314
rect 4921 28260 4977 28262
rect 5001 28260 5057 28262
rect 5081 28260 5137 28262
rect 5161 28260 5217 28262
rect 4894 28056 4950 28112
rect 4921 27226 4977 27228
rect 5001 27226 5057 27228
rect 5081 27226 5137 27228
rect 5161 27226 5217 27228
rect 4921 27174 4947 27226
rect 4947 27174 4977 27226
rect 5001 27174 5011 27226
rect 5011 27174 5057 27226
rect 5081 27174 5127 27226
rect 5127 27174 5137 27226
rect 5161 27174 5191 27226
rect 5191 27174 5217 27226
rect 4921 27172 4977 27174
rect 5001 27172 5057 27174
rect 5081 27172 5137 27174
rect 5161 27172 5217 27174
rect 4921 26138 4977 26140
rect 5001 26138 5057 26140
rect 5081 26138 5137 26140
rect 5161 26138 5217 26140
rect 4921 26086 4947 26138
rect 4947 26086 4977 26138
rect 5001 26086 5011 26138
rect 5011 26086 5057 26138
rect 5081 26086 5127 26138
rect 5127 26086 5137 26138
rect 5161 26086 5191 26138
rect 5191 26086 5217 26138
rect 4921 26084 4977 26086
rect 5001 26084 5057 26086
rect 5081 26084 5137 26086
rect 5161 26084 5217 26086
rect 4921 25050 4977 25052
rect 5001 25050 5057 25052
rect 5081 25050 5137 25052
rect 5161 25050 5217 25052
rect 4921 24998 4947 25050
rect 4947 24998 4977 25050
rect 5001 24998 5011 25050
rect 5011 24998 5057 25050
rect 5081 24998 5127 25050
rect 5127 24998 5137 25050
rect 5161 24998 5191 25050
rect 5191 24998 5217 25050
rect 4921 24996 4977 24998
rect 5001 24996 5057 24998
rect 5081 24996 5137 24998
rect 5161 24996 5217 24998
rect 4921 23962 4977 23964
rect 5001 23962 5057 23964
rect 5081 23962 5137 23964
rect 5161 23962 5217 23964
rect 4921 23910 4947 23962
rect 4947 23910 4977 23962
rect 5001 23910 5011 23962
rect 5011 23910 5057 23962
rect 5081 23910 5127 23962
rect 5127 23910 5137 23962
rect 5161 23910 5191 23962
rect 5191 23910 5217 23962
rect 4921 23908 4977 23910
rect 5001 23908 5057 23910
rect 5081 23908 5137 23910
rect 5161 23908 5217 23910
rect 4921 22874 4977 22876
rect 5001 22874 5057 22876
rect 5081 22874 5137 22876
rect 5161 22874 5217 22876
rect 4921 22822 4947 22874
rect 4947 22822 4977 22874
rect 5001 22822 5011 22874
rect 5011 22822 5057 22874
rect 5081 22822 5127 22874
rect 5127 22822 5137 22874
rect 5161 22822 5191 22874
rect 5191 22822 5217 22874
rect 4921 22820 4977 22822
rect 5001 22820 5057 22822
rect 5081 22820 5137 22822
rect 5161 22820 5217 22822
rect 5354 23024 5410 23080
rect 4921 21786 4977 21788
rect 5001 21786 5057 21788
rect 5081 21786 5137 21788
rect 5161 21786 5217 21788
rect 4921 21734 4947 21786
rect 4947 21734 4977 21786
rect 5001 21734 5011 21786
rect 5011 21734 5057 21786
rect 5081 21734 5127 21786
rect 5127 21734 5137 21786
rect 5161 21734 5191 21786
rect 5191 21734 5217 21786
rect 4921 21732 4977 21734
rect 5001 21732 5057 21734
rect 5081 21732 5137 21734
rect 5161 21732 5217 21734
rect 4921 20698 4977 20700
rect 5001 20698 5057 20700
rect 5081 20698 5137 20700
rect 5161 20698 5217 20700
rect 4921 20646 4947 20698
rect 4947 20646 4977 20698
rect 5001 20646 5011 20698
rect 5011 20646 5057 20698
rect 5081 20646 5127 20698
rect 5127 20646 5137 20698
rect 5161 20646 5191 20698
rect 5191 20646 5217 20698
rect 4921 20644 4977 20646
rect 5001 20644 5057 20646
rect 5081 20644 5137 20646
rect 5161 20644 5217 20646
rect 4921 19610 4977 19612
rect 5001 19610 5057 19612
rect 5081 19610 5137 19612
rect 5161 19610 5217 19612
rect 4921 19558 4947 19610
rect 4947 19558 4977 19610
rect 5001 19558 5011 19610
rect 5011 19558 5057 19610
rect 5081 19558 5127 19610
rect 5127 19558 5137 19610
rect 5161 19558 5191 19610
rect 5191 19558 5217 19610
rect 4921 19556 4977 19558
rect 5001 19556 5057 19558
rect 5081 19556 5137 19558
rect 5161 19556 5217 19558
rect 4986 19352 5042 19408
rect 4986 18672 5042 18728
rect 4921 18522 4977 18524
rect 5001 18522 5057 18524
rect 5081 18522 5137 18524
rect 5161 18522 5217 18524
rect 4921 18470 4947 18522
rect 4947 18470 4977 18522
rect 5001 18470 5011 18522
rect 5011 18470 5057 18522
rect 5081 18470 5127 18522
rect 5127 18470 5137 18522
rect 5161 18470 5191 18522
rect 5191 18470 5217 18522
rect 4921 18468 4977 18470
rect 5001 18468 5057 18470
rect 5081 18468 5137 18470
rect 5161 18468 5217 18470
rect 4921 17434 4977 17436
rect 5001 17434 5057 17436
rect 5081 17434 5137 17436
rect 5161 17434 5217 17436
rect 4921 17382 4947 17434
rect 4947 17382 4977 17434
rect 5001 17382 5011 17434
rect 5011 17382 5057 17434
rect 5081 17382 5127 17434
rect 5127 17382 5137 17434
rect 5161 17382 5191 17434
rect 5191 17382 5217 17434
rect 4921 17380 4977 17382
rect 5001 17380 5057 17382
rect 5081 17380 5137 17382
rect 5161 17380 5217 17382
rect 4921 16346 4977 16348
rect 5001 16346 5057 16348
rect 5081 16346 5137 16348
rect 5161 16346 5217 16348
rect 4921 16294 4947 16346
rect 4947 16294 4977 16346
rect 5001 16294 5011 16346
rect 5011 16294 5057 16346
rect 5081 16294 5127 16346
rect 5127 16294 5137 16346
rect 5161 16294 5191 16346
rect 5191 16294 5217 16346
rect 4921 16292 4977 16294
rect 5001 16292 5057 16294
rect 5081 16292 5137 16294
rect 5161 16292 5217 16294
rect 4921 15258 4977 15260
rect 5001 15258 5057 15260
rect 5081 15258 5137 15260
rect 5161 15258 5217 15260
rect 4921 15206 4947 15258
rect 4947 15206 4977 15258
rect 5001 15206 5011 15258
rect 5011 15206 5057 15258
rect 5081 15206 5127 15258
rect 5127 15206 5137 15258
rect 5161 15206 5191 15258
rect 5191 15206 5217 15258
rect 4921 15204 4977 15206
rect 5001 15204 5057 15206
rect 5081 15204 5137 15206
rect 5161 15204 5217 15206
rect 4921 14170 4977 14172
rect 5001 14170 5057 14172
rect 5081 14170 5137 14172
rect 5161 14170 5217 14172
rect 4921 14118 4947 14170
rect 4947 14118 4977 14170
rect 5001 14118 5011 14170
rect 5011 14118 5057 14170
rect 5081 14118 5127 14170
rect 5127 14118 5137 14170
rect 5161 14118 5191 14170
rect 5191 14118 5217 14170
rect 4921 14116 4977 14118
rect 5001 14116 5057 14118
rect 5081 14116 5137 14118
rect 5161 14116 5217 14118
rect 4921 13082 4977 13084
rect 5001 13082 5057 13084
rect 5081 13082 5137 13084
rect 5161 13082 5217 13084
rect 4921 13030 4947 13082
rect 4947 13030 4977 13082
rect 5001 13030 5011 13082
rect 5011 13030 5057 13082
rect 5081 13030 5127 13082
rect 5127 13030 5137 13082
rect 5161 13030 5191 13082
rect 5191 13030 5217 13082
rect 4921 13028 4977 13030
rect 5001 13028 5057 13030
rect 5081 13028 5137 13030
rect 5161 13028 5217 13030
rect 5170 12844 5226 12880
rect 5170 12824 5172 12844
rect 5172 12824 5224 12844
rect 5224 12824 5226 12844
rect 4434 9016 4490 9072
rect 4434 8492 4490 8528
rect 4434 8472 4436 8492
rect 4436 8472 4488 8492
rect 4488 8472 4490 8492
rect 4921 11994 4977 11996
rect 5001 11994 5057 11996
rect 5081 11994 5137 11996
rect 5161 11994 5217 11996
rect 4921 11942 4947 11994
rect 4947 11942 4977 11994
rect 5001 11942 5011 11994
rect 5011 11942 5057 11994
rect 5081 11942 5127 11994
rect 5127 11942 5137 11994
rect 5161 11942 5191 11994
rect 5191 11942 5217 11994
rect 4921 11940 4977 11942
rect 5001 11940 5057 11942
rect 5081 11940 5137 11942
rect 5161 11940 5217 11942
rect 4921 10906 4977 10908
rect 5001 10906 5057 10908
rect 5081 10906 5137 10908
rect 5161 10906 5217 10908
rect 4921 10854 4947 10906
rect 4947 10854 4977 10906
rect 5001 10854 5011 10906
rect 5011 10854 5057 10906
rect 5081 10854 5127 10906
rect 5127 10854 5137 10906
rect 5161 10854 5191 10906
rect 5191 10854 5217 10906
rect 4921 10852 4977 10854
rect 5001 10852 5057 10854
rect 5081 10852 5137 10854
rect 5161 10852 5217 10854
rect 4921 9818 4977 9820
rect 5001 9818 5057 9820
rect 5081 9818 5137 9820
rect 5161 9818 5217 9820
rect 4921 9766 4947 9818
rect 4947 9766 4977 9818
rect 5001 9766 5011 9818
rect 5011 9766 5057 9818
rect 5081 9766 5127 9818
rect 5127 9766 5137 9818
rect 5161 9766 5191 9818
rect 5191 9766 5217 9818
rect 4921 9764 4977 9766
rect 5001 9764 5057 9766
rect 5081 9764 5137 9766
rect 5161 9764 5217 9766
rect 4894 9560 4950 9616
rect 5170 9424 5226 9480
rect 4921 8730 4977 8732
rect 5001 8730 5057 8732
rect 5081 8730 5137 8732
rect 5161 8730 5217 8732
rect 4921 8678 4947 8730
rect 4947 8678 4977 8730
rect 5001 8678 5011 8730
rect 5011 8678 5057 8730
rect 5081 8678 5127 8730
rect 5127 8678 5137 8730
rect 5161 8678 5191 8730
rect 5191 8678 5217 8730
rect 4921 8676 4977 8678
rect 5001 8676 5057 8678
rect 5081 8676 5137 8678
rect 5161 8676 5217 8678
rect 5446 13776 5502 13832
rect 4921 7642 4977 7644
rect 5001 7642 5057 7644
rect 5081 7642 5137 7644
rect 5161 7642 5217 7644
rect 4921 7590 4947 7642
rect 4947 7590 4977 7642
rect 5001 7590 5011 7642
rect 5011 7590 5057 7642
rect 5081 7590 5127 7642
rect 5127 7590 5137 7642
rect 5161 7590 5191 7642
rect 5191 7590 5217 7642
rect 4921 7588 4977 7590
rect 5001 7588 5057 7590
rect 5081 7588 5137 7590
rect 5161 7588 5217 7590
rect 4921 6554 4977 6556
rect 5001 6554 5057 6556
rect 5081 6554 5137 6556
rect 5161 6554 5217 6556
rect 4921 6502 4947 6554
rect 4947 6502 4977 6554
rect 5001 6502 5011 6554
rect 5011 6502 5057 6554
rect 5081 6502 5127 6554
rect 5127 6502 5137 6554
rect 5161 6502 5191 6554
rect 5191 6502 5217 6554
rect 4921 6500 4977 6502
rect 5001 6500 5057 6502
rect 5081 6500 5137 6502
rect 5161 6500 5217 6502
rect 5630 9424 5686 9480
rect 4921 5466 4977 5468
rect 5001 5466 5057 5468
rect 5081 5466 5137 5468
rect 5161 5466 5217 5468
rect 4921 5414 4947 5466
rect 4947 5414 4977 5466
rect 5001 5414 5011 5466
rect 5011 5414 5057 5466
rect 5081 5414 5127 5466
rect 5127 5414 5137 5466
rect 5161 5414 5191 5466
rect 5191 5414 5217 5466
rect 4921 5412 4977 5414
rect 5001 5412 5057 5414
rect 5081 5412 5137 5414
rect 5161 5412 5217 5414
rect 4921 4378 4977 4380
rect 5001 4378 5057 4380
rect 5081 4378 5137 4380
rect 5161 4378 5217 4380
rect 4921 4326 4947 4378
rect 4947 4326 4977 4378
rect 5001 4326 5011 4378
rect 5011 4326 5057 4378
rect 5081 4326 5127 4378
rect 5127 4326 5137 4378
rect 5161 4326 5191 4378
rect 5191 4326 5217 4378
rect 4921 4324 4977 4326
rect 5001 4324 5057 4326
rect 5081 4324 5137 4326
rect 5161 4324 5217 4326
rect 4921 3290 4977 3292
rect 5001 3290 5057 3292
rect 5081 3290 5137 3292
rect 5161 3290 5217 3292
rect 4921 3238 4947 3290
rect 4947 3238 4977 3290
rect 5001 3238 5011 3290
rect 5011 3238 5057 3290
rect 5081 3238 5127 3290
rect 5127 3238 5137 3290
rect 5161 3238 5191 3290
rect 5191 3238 5217 3290
rect 4921 3236 4977 3238
rect 5001 3236 5057 3238
rect 5081 3236 5137 3238
rect 5161 3236 5217 3238
rect 5906 9560 5962 9616
rect 4921 2202 4977 2204
rect 5001 2202 5057 2204
rect 5081 2202 5137 2204
rect 5161 2202 5217 2204
rect 4921 2150 4947 2202
rect 4947 2150 4977 2202
rect 5001 2150 5011 2202
rect 5011 2150 5057 2202
rect 5081 2150 5127 2202
rect 5127 2150 5137 2202
rect 5161 2150 5191 2202
rect 5191 2150 5217 2202
rect 4921 2148 4977 2150
rect 5001 2148 5057 2150
rect 5081 2148 5137 2150
rect 5161 2148 5217 2150
rect 5446 1808 5502 1864
rect 6090 9560 6146 9616
rect 6550 21528 6606 21584
rect 8886 46266 8942 46268
rect 8966 46266 9022 46268
rect 9046 46266 9102 46268
rect 9126 46266 9182 46268
rect 8886 46214 8912 46266
rect 8912 46214 8942 46266
rect 8966 46214 8976 46266
rect 8976 46214 9022 46266
rect 9046 46214 9092 46266
rect 9092 46214 9102 46266
rect 9126 46214 9156 46266
rect 9156 46214 9182 46266
rect 8886 46212 8942 46214
rect 8966 46212 9022 46214
rect 9046 46212 9102 46214
rect 9126 46212 9182 46214
rect 7930 38936 7986 38992
rect 6826 22344 6882 22400
rect 6826 20748 6828 20768
rect 6828 20748 6880 20768
rect 6880 20748 6882 20768
rect 6826 20712 6882 20748
rect 7194 22344 7250 22400
rect 6918 19896 6974 19952
rect 7562 22752 7618 22808
rect 7470 21936 7526 21992
rect 7470 21800 7526 21856
rect 7378 18944 7434 19000
rect 7562 21664 7618 21720
rect 7746 21548 7802 21584
rect 7746 21528 7748 21548
rect 7748 21528 7800 21548
rect 7800 21528 7802 21548
rect 7102 10240 7158 10296
rect 7930 22752 7986 22808
rect 8886 45178 8942 45180
rect 8966 45178 9022 45180
rect 9046 45178 9102 45180
rect 9126 45178 9182 45180
rect 8886 45126 8912 45178
rect 8912 45126 8942 45178
rect 8966 45126 8976 45178
rect 8976 45126 9022 45178
rect 9046 45126 9092 45178
rect 9092 45126 9102 45178
rect 9126 45126 9156 45178
rect 9156 45126 9182 45178
rect 8886 45124 8942 45126
rect 8966 45124 9022 45126
rect 9046 45124 9102 45126
rect 9126 45124 9182 45126
rect 8886 44090 8942 44092
rect 8966 44090 9022 44092
rect 9046 44090 9102 44092
rect 9126 44090 9182 44092
rect 8886 44038 8912 44090
rect 8912 44038 8942 44090
rect 8966 44038 8976 44090
rect 8976 44038 9022 44090
rect 9046 44038 9092 44090
rect 9092 44038 9102 44090
rect 9126 44038 9156 44090
rect 9156 44038 9182 44090
rect 8886 44036 8942 44038
rect 8966 44036 9022 44038
rect 9046 44036 9102 44038
rect 9126 44036 9182 44038
rect 8886 43002 8942 43004
rect 8966 43002 9022 43004
rect 9046 43002 9102 43004
rect 9126 43002 9182 43004
rect 8886 42950 8912 43002
rect 8912 42950 8942 43002
rect 8966 42950 8976 43002
rect 8976 42950 9022 43002
rect 9046 42950 9092 43002
rect 9092 42950 9102 43002
rect 9126 42950 9156 43002
rect 9156 42950 9182 43002
rect 8886 42948 8942 42950
rect 8966 42948 9022 42950
rect 9046 42948 9102 42950
rect 9126 42948 9182 42950
rect 8886 41914 8942 41916
rect 8966 41914 9022 41916
rect 9046 41914 9102 41916
rect 9126 41914 9182 41916
rect 8886 41862 8912 41914
rect 8912 41862 8942 41914
rect 8966 41862 8976 41914
rect 8976 41862 9022 41914
rect 9046 41862 9092 41914
rect 9092 41862 9102 41914
rect 9126 41862 9156 41914
rect 9156 41862 9182 41914
rect 8886 41860 8942 41862
rect 8966 41860 9022 41862
rect 9046 41860 9102 41862
rect 9126 41860 9182 41862
rect 8886 40826 8942 40828
rect 8966 40826 9022 40828
rect 9046 40826 9102 40828
rect 9126 40826 9182 40828
rect 8886 40774 8912 40826
rect 8912 40774 8942 40826
rect 8966 40774 8976 40826
rect 8976 40774 9022 40826
rect 9046 40774 9092 40826
rect 9092 40774 9102 40826
rect 9126 40774 9156 40826
rect 9156 40774 9182 40826
rect 8886 40772 8942 40774
rect 8966 40772 9022 40774
rect 9046 40772 9102 40774
rect 9126 40772 9182 40774
rect 8886 39738 8942 39740
rect 8966 39738 9022 39740
rect 9046 39738 9102 39740
rect 9126 39738 9182 39740
rect 8886 39686 8912 39738
rect 8912 39686 8942 39738
rect 8966 39686 8976 39738
rect 8976 39686 9022 39738
rect 9046 39686 9092 39738
rect 9092 39686 9102 39738
rect 9126 39686 9156 39738
rect 9156 39686 9182 39738
rect 8886 39684 8942 39686
rect 8966 39684 9022 39686
rect 9046 39684 9102 39686
rect 9126 39684 9182 39686
rect 8298 28464 8354 28520
rect 8886 38650 8942 38652
rect 8966 38650 9022 38652
rect 9046 38650 9102 38652
rect 9126 38650 9182 38652
rect 8886 38598 8912 38650
rect 8912 38598 8942 38650
rect 8966 38598 8976 38650
rect 8976 38598 9022 38650
rect 9046 38598 9092 38650
rect 9092 38598 9102 38650
rect 9126 38598 9156 38650
rect 9156 38598 9182 38650
rect 8886 38596 8942 38598
rect 8966 38596 9022 38598
rect 9046 38596 9102 38598
rect 9126 38596 9182 38598
rect 8886 37562 8942 37564
rect 8966 37562 9022 37564
rect 9046 37562 9102 37564
rect 9126 37562 9182 37564
rect 8886 37510 8912 37562
rect 8912 37510 8942 37562
rect 8966 37510 8976 37562
rect 8976 37510 9022 37562
rect 9046 37510 9092 37562
rect 9092 37510 9102 37562
rect 9126 37510 9156 37562
rect 9156 37510 9182 37562
rect 8886 37508 8942 37510
rect 8966 37508 9022 37510
rect 9046 37508 9102 37510
rect 9126 37508 9182 37510
rect 8886 36474 8942 36476
rect 8966 36474 9022 36476
rect 9046 36474 9102 36476
rect 9126 36474 9182 36476
rect 8886 36422 8912 36474
rect 8912 36422 8942 36474
rect 8966 36422 8976 36474
rect 8976 36422 9022 36474
rect 9046 36422 9092 36474
rect 9092 36422 9102 36474
rect 9126 36422 9156 36474
rect 9156 36422 9182 36474
rect 8886 36420 8942 36422
rect 8966 36420 9022 36422
rect 9046 36420 9102 36422
rect 9126 36420 9182 36422
rect 8886 35386 8942 35388
rect 8966 35386 9022 35388
rect 9046 35386 9102 35388
rect 9126 35386 9182 35388
rect 8886 35334 8912 35386
rect 8912 35334 8942 35386
rect 8966 35334 8976 35386
rect 8976 35334 9022 35386
rect 9046 35334 9092 35386
rect 9092 35334 9102 35386
rect 9126 35334 9156 35386
rect 9156 35334 9182 35386
rect 8886 35332 8942 35334
rect 8966 35332 9022 35334
rect 9046 35332 9102 35334
rect 9126 35332 9182 35334
rect 8886 34298 8942 34300
rect 8966 34298 9022 34300
rect 9046 34298 9102 34300
rect 9126 34298 9182 34300
rect 8886 34246 8912 34298
rect 8912 34246 8942 34298
rect 8966 34246 8976 34298
rect 8976 34246 9022 34298
rect 9046 34246 9092 34298
rect 9092 34246 9102 34298
rect 9126 34246 9156 34298
rect 9156 34246 9182 34298
rect 8886 34244 8942 34246
rect 8966 34244 9022 34246
rect 9046 34244 9102 34246
rect 9126 34244 9182 34246
rect 8886 33210 8942 33212
rect 8966 33210 9022 33212
rect 9046 33210 9102 33212
rect 9126 33210 9182 33212
rect 8886 33158 8912 33210
rect 8912 33158 8942 33210
rect 8966 33158 8976 33210
rect 8976 33158 9022 33210
rect 9046 33158 9092 33210
rect 9092 33158 9102 33210
rect 9126 33158 9156 33210
rect 9156 33158 9182 33210
rect 8886 33156 8942 33158
rect 8966 33156 9022 33158
rect 9046 33156 9102 33158
rect 9126 33156 9182 33158
rect 9586 38972 9588 38992
rect 9588 38972 9640 38992
rect 9640 38972 9642 38992
rect 9586 38936 9642 38972
rect 8886 32122 8942 32124
rect 8966 32122 9022 32124
rect 9046 32122 9102 32124
rect 9126 32122 9182 32124
rect 8886 32070 8912 32122
rect 8912 32070 8942 32122
rect 8966 32070 8976 32122
rect 8976 32070 9022 32122
rect 9046 32070 9092 32122
rect 9092 32070 9102 32122
rect 9126 32070 9156 32122
rect 9156 32070 9182 32122
rect 8886 32068 8942 32070
rect 8966 32068 9022 32070
rect 9046 32068 9102 32070
rect 9126 32068 9182 32070
rect 8886 31034 8942 31036
rect 8966 31034 9022 31036
rect 9046 31034 9102 31036
rect 9126 31034 9182 31036
rect 8886 30982 8912 31034
rect 8912 30982 8942 31034
rect 8966 30982 8976 31034
rect 8976 30982 9022 31034
rect 9046 30982 9092 31034
rect 9092 30982 9102 31034
rect 9126 30982 9156 31034
rect 9156 30982 9182 31034
rect 8886 30980 8942 30982
rect 8966 30980 9022 30982
rect 9046 30980 9102 30982
rect 9126 30980 9182 30982
rect 8482 27240 8538 27296
rect 8298 27004 8300 27024
rect 8300 27004 8352 27024
rect 8352 27004 8354 27024
rect 8298 26968 8354 27004
rect 8298 26732 8300 26752
rect 8300 26732 8352 26752
rect 8352 26732 8354 26752
rect 8298 26696 8354 26732
rect 8206 22072 8262 22128
rect 8886 29946 8942 29948
rect 8966 29946 9022 29948
rect 9046 29946 9102 29948
rect 9126 29946 9182 29948
rect 8886 29894 8912 29946
rect 8912 29894 8942 29946
rect 8966 29894 8976 29946
rect 8976 29894 9022 29946
rect 9046 29894 9092 29946
rect 9092 29894 9102 29946
rect 9126 29894 9156 29946
rect 9156 29894 9182 29946
rect 8886 29892 8942 29894
rect 8966 29892 9022 29894
rect 9046 29892 9102 29894
rect 9126 29892 9182 29894
rect 8666 26968 8722 27024
rect 8666 26696 8722 26752
rect 8482 22616 8538 22672
rect 8390 20712 8446 20768
rect 8390 19760 8446 19816
rect 6826 4936 6882 4992
rect 7286 7792 7342 7848
rect 8206 12416 8262 12472
rect 8206 12280 8262 12336
rect 8298 9052 8300 9072
rect 8300 9052 8352 9072
rect 8352 9052 8354 9072
rect 8298 9016 8354 9052
rect 8886 28858 8942 28860
rect 8966 28858 9022 28860
rect 9046 28858 9102 28860
rect 9126 28858 9182 28860
rect 8886 28806 8912 28858
rect 8912 28806 8942 28858
rect 8966 28806 8976 28858
rect 8976 28806 9022 28858
rect 9046 28806 9092 28858
rect 9092 28806 9102 28858
rect 9126 28806 9156 28858
rect 9156 28806 9182 28858
rect 8886 28804 8942 28806
rect 8966 28804 9022 28806
rect 9046 28804 9102 28806
rect 9126 28804 9182 28806
rect 8886 27770 8942 27772
rect 8966 27770 9022 27772
rect 9046 27770 9102 27772
rect 9126 27770 9182 27772
rect 8886 27718 8912 27770
rect 8912 27718 8942 27770
rect 8966 27718 8976 27770
rect 8976 27718 9022 27770
rect 9046 27718 9092 27770
rect 9092 27718 9102 27770
rect 9126 27718 9156 27770
rect 9156 27718 9182 27770
rect 8886 27716 8942 27718
rect 8966 27716 9022 27718
rect 9046 27716 9102 27718
rect 9126 27716 9182 27718
rect 8886 26682 8942 26684
rect 8966 26682 9022 26684
rect 9046 26682 9102 26684
rect 9126 26682 9182 26684
rect 8886 26630 8912 26682
rect 8912 26630 8942 26682
rect 8966 26630 8976 26682
rect 8976 26630 9022 26682
rect 9046 26630 9092 26682
rect 9092 26630 9102 26682
rect 9126 26630 9156 26682
rect 9156 26630 9182 26682
rect 8886 26628 8942 26630
rect 8966 26628 9022 26630
rect 9046 26628 9102 26630
rect 9126 26628 9182 26630
rect 8886 25594 8942 25596
rect 8966 25594 9022 25596
rect 9046 25594 9102 25596
rect 9126 25594 9182 25596
rect 8886 25542 8912 25594
rect 8912 25542 8942 25594
rect 8966 25542 8976 25594
rect 8976 25542 9022 25594
rect 9046 25542 9092 25594
rect 9092 25542 9102 25594
rect 9126 25542 9156 25594
rect 9156 25542 9182 25594
rect 8886 25540 8942 25542
rect 8966 25540 9022 25542
rect 9046 25540 9102 25542
rect 9126 25540 9182 25542
rect 9218 24792 9274 24848
rect 8886 24506 8942 24508
rect 8966 24506 9022 24508
rect 9046 24506 9102 24508
rect 9126 24506 9182 24508
rect 8886 24454 8912 24506
rect 8912 24454 8942 24506
rect 8966 24454 8976 24506
rect 8976 24454 9022 24506
rect 9046 24454 9092 24506
rect 9092 24454 9102 24506
rect 9126 24454 9156 24506
rect 9156 24454 9182 24506
rect 8886 24452 8942 24454
rect 8966 24452 9022 24454
rect 9046 24452 9102 24454
rect 9126 24452 9182 24454
rect 8886 23418 8942 23420
rect 8966 23418 9022 23420
rect 9046 23418 9102 23420
rect 9126 23418 9182 23420
rect 8886 23366 8912 23418
rect 8912 23366 8942 23418
rect 8966 23366 8976 23418
rect 8976 23366 9022 23418
rect 9046 23366 9092 23418
rect 9092 23366 9102 23418
rect 9126 23366 9156 23418
rect 9156 23366 9182 23418
rect 8886 23364 8942 23366
rect 8966 23364 9022 23366
rect 9046 23364 9102 23366
rect 9126 23364 9182 23366
rect 8886 22330 8942 22332
rect 8966 22330 9022 22332
rect 9046 22330 9102 22332
rect 9126 22330 9182 22332
rect 8886 22278 8912 22330
rect 8912 22278 8942 22330
rect 8966 22278 8976 22330
rect 8976 22278 9022 22330
rect 9046 22278 9092 22330
rect 9092 22278 9102 22330
rect 9126 22278 9156 22330
rect 9156 22278 9182 22330
rect 8886 22276 8942 22278
rect 8966 22276 9022 22278
rect 9046 22276 9102 22278
rect 9126 22276 9182 22278
rect 9218 21392 9274 21448
rect 8886 21242 8942 21244
rect 8966 21242 9022 21244
rect 9046 21242 9102 21244
rect 9126 21242 9182 21244
rect 8886 21190 8912 21242
rect 8912 21190 8942 21242
rect 8966 21190 8976 21242
rect 8976 21190 9022 21242
rect 9046 21190 9092 21242
rect 9092 21190 9102 21242
rect 9126 21190 9156 21242
rect 9156 21190 9182 21242
rect 8886 21188 8942 21190
rect 8966 21188 9022 21190
rect 9046 21188 9102 21190
rect 9126 21188 9182 21190
rect 9126 21004 9182 21040
rect 9126 20984 9128 21004
rect 9128 20984 9180 21004
rect 9180 20984 9182 21004
rect 8850 20440 8906 20496
rect 8886 20154 8942 20156
rect 8966 20154 9022 20156
rect 9046 20154 9102 20156
rect 9126 20154 9182 20156
rect 8886 20102 8912 20154
rect 8912 20102 8942 20154
rect 8966 20102 8976 20154
rect 8976 20102 9022 20154
rect 9046 20102 9092 20154
rect 9092 20102 9102 20154
rect 9126 20102 9156 20154
rect 9156 20102 9182 20154
rect 8886 20100 8942 20102
rect 8966 20100 9022 20102
rect 9046 20100 9102 20102
rect 9126 20100 9182 20102
rect 8886 19066 8942 19068
rect 8966 19066 9022 19068
rect 9046 19066 9102 19068
rect 9126 19066 9182 19068
rect 8886 19014 8912 19066
rect 8912 19014 8942 19066
rect 8966 19014 8976 19066
rect 8976 19014 9022 19066
rect 9046 19014 9092 19066
rect 9092 19014 9102 19066
rect 9126 19014 9156 19066
rect 9156 19014 9182 19066
rect 8886 19012 8942 19014
rect 8966 19012 9022 19014
rect 9046 19012 9102 19014
rect 9126 19012 9182 19014
rect 8886 17978 8942 17980
rect 8966 17978 9022 17980
rect 9046 17978 9102 17980
rect 9126 17978 9182 17980
rect 8886 17926 8912 17978
rect 8912 17926 8942 17978
rect 8966 17926 8976 17978
rect 8976 17926 9022 17978
rect 9046 17926 9092 17978
rect 9092 17926 9102 17978
rect 9126 17926 9156 17978
rect 9156 17926 9182 17978
rect 8886 17924 8942 17926
rect 8966 17924 9022 17926
rect 9046 17924 9102 17926
rect 9126 17924 9182 17926
rect 8886 16890 8942 16892
rect 8966 16890 9022 16892
rect 9046 16890 9102 16892
rect 9126 16890 9182 16892
rect 8886 16838 8912 16890
rect 8912 16838 8942 16890
rect 8966 16838 8976 16890
rect 8976 16838 9022 16890
rect 9046 16838 9092 16890
rect 9092 16838 9102 16890
rect 9126 16838 9156 16890
rect 9156 16838 9182 16890
rect 8886 16836 8942 16838
rect 8966 16836 9022 16838
rect 9046 16836 9102 16838
rect 9126 16836 9182 16838
rect 8886 15802 8942 15804
rect 8966 15802 9022 15804
rect 9046 15802 9102 15804
rect 9126 15802 9182 15804
rect 8886 15750 8912 15802
rect 8912 15750 8942 15802
rect 8966 15750 8976 15802
rect 8976 15750 9022 15802
rect 9046 15750 9092 15802
rect 9092 15750 9102 15802
rect 9126 15750 9156 15802
rect 9156 15750 9182 15802
rect 8886 15748 8942 15750
rect 8966 15748 9022 15750
rect 9046 15748 9102 15750
rect 9126 15748 9182 15750
rect 8886 14714 8942 14716
rect 8966 14714 9022 14716
rect 9046 14714 9102 14716
rect 9126 14714 9182 14716
rect 8886 14662 8912 14714
rect 8912 14662 8942 14714
rect 8966 14662 8976 14714
rect 8976 14662 9022 14714
rect 9046 14662 9092 14714
rect 9092 14662 9102 14714
rect 9126 14662 9156 14714
rect 9156 14662 9182 14714
rect 8886 14660 8942 14662
rect 8966 14660 9022 14662
rect 9046 14660 9102 14662
rect 9126 14660 9182 14662
rect 8886 13626 8942 13628
rect 8966 13626 9022 13628
rect 9046 13626 9102 13628
rect 9126 13626 9182 13628
rect 8886 13574 8912 13626
rect 8912 13574 8942 13626
rect 8966 13574 8976 13626
rect 8976 13574 9022 13626
rect 9046 13574 9092 13626
rect 9092 13574 9102 13626
rect 9126 13574 9156 13626
rect 9156 13574 9182 13626
rect 8886 13572 8942 13574
rect 8966 13572 9022 13574
rect 9046 13572 9102 13574
rect 9126 13572 9182 13574
rect 8886 12538 8942 12540
rect 8966 12538 9022 12540
rect 9046 12538 9102 12540
rect 9126 12538 9182 12540
rect 8886 12486 8912 12538
rect 8912 12486 8942 12538
rect 8966 12486 8976 12538
rect 8976 12486 9022 12538
rect 9046 12486 9092 12538
rect 9092 12486 9102 12538
rect 9126 12486 9156 12538
rect 9156 12486 9182 12538
rect 8886 12484 8942 12486
rect 8966 12484 9022 12486
rect 9046 12484 9102 12486
rect 9126 12484 9182 12486
rect 8886 11450 8942 11452
rect 8966 11450 9022 11452
rect 9046 11450 9102 11452
rect 9126 11450 9182 11452
rect 8886 11398 8912 11450
rect 8912 11398 8942 11450
rect 8966 11398 8976 11450
rect 8976 11398 9022 11450
rect 9046 11398 9092 11450
rect 9092 11398 9102 11450
rect 9126 11398 9156 11450
rect 9156 11398 9182 11450
rect 8886 11396 8942 11398
rect 8966 11396 9022 11398
rect 9046 11396 9102 11398
rect 9126 11396 9182 11398
rect 8886 10362 8942 10364
rect 8966 10362 9022 10364
rect 9046 10362 9102 10364
rect 9126 10362 9182 10364
rect 8886 10310 8912 10362
rect 8912 10310 8942 10362
rect 8966 10310 8976 10362
rect 8976 10310 9022 10362
rect 9046 10310 9092 10362
rect 9092 10310 9102 10362
rect 9126 10310 9156 10362
rect 9156 10310 9182 10362
rect 8886 10308 8942 10310
rect 8966 10308 9022 10310
rect 9046 10308 9102 10310
rect 9126 10308 9182 10310
rect 8886 9274 8942 9276
rect 8966 9274 9022 9276
rect 9046 9274 9102 9276
rect 9126 9274 9182 9276
rect 8886 9222 8912 9274
rect 8912 9222 8942 9274
rect 8966 9222 8976 9274
rect 8976 9222 9022 9274
rect 9046 9222 9092 9274
rect 9092 9222 9102 9274
rect 9126 9222 9156 9274
rect 9156 9222 9182 9274
rect 8886 9220 8942 9222
rect 8966 9220 9022 9222
rect 9046 9220 9102 9222
rect 9126 9220 9182 9222
rect 8886 8186 8942 8188
rect 8966 8186 9022 8188
rect 9046 8186 9102 8188
rect 9126 8186 9182 8188
rect 8886 8134 8912 8186
rect 8912 8134 8942 8186
rect 8966 8134 8976 8186
rect 8976 8134 9022 8186
rect 9046 8134 9092 8186
rect 9092 8134 9102 8186
rect 9126 8134 9156 8186
rect 9156 8134 9182 8186
rect 8886 8132 8942 8134
rect 8966 8132 9022 8134
rect 9046 8132 9102 8134
rect 9126 8132 9182 8134
rect 8886 7098 8942 7100
rect 8966 7098 9022 7100
rect 9046 7098 9102 7100
rect 9126 7098 9182 7100
rect 8886 7046 8912 7098
rect 8912 7046 8942 7098
rect 8966 7046 8976 7098
rect 8976 7046 9022 7098
rect 9046 7046 9092 7098
rect 9092 7046 9102 7098
rect 9126 7046 9156 7098
rect 9156 7046 9182 7098
rect 8886 7044 8942 7046
rect 8966 7044 9022 7046
rect 9046 7044 9102 7046
rect 9126 7044 9182 7046
rect 8886 6010 8942 6012
rect 8966 6010 9022 6012
rect 9046 6010 9102 6012
rect 9126 6010 9182 6012
rect 8886 5958 8912 6010
rect 8912 5958 8942 6010
rect 8966 5958 8976 6010
rect 8976 5958 9022 6010
rect 9046 5958 9092 6010
rect 9092 5958 9102 6010
rect 9126 5958 9156 6010
rect 9156 5958 9182 6010
rect 8886 5956 8942 5958
rect 8966 5956 9022 5958
rect 9046 5956 9102 5958
rect 9126 5956 9182 5958
rect 8886 4922 8942 4924
rect 8966 4922 9022 4924
rect 9046 4922 9102 4924
rect 9126 4922 9182 4924
rect 8886 4870 8912 4922
rect 8912 4870 8942 4922
rect 8966 4870 8976 4922
rect 8976 4870 9022 4922
rect 9046 4870 9092 4922
rect 9092 4870 9102 4922
rect 9126 4870 9156 4922
rect 9156 4870 9182 4922
rect 8886 4868 8942 4870
rect 8966 4868 9022 4870
rect 9046 4868 9102 4870
rect 9126 4868 9182 4870
rect 8886 3834 8942 3836
rect 8966 3834 9022 3836
rect 9046 3834 9102 3836
rect 9126 3834 9182 3836
rect 8886 3782 8912 3834
rect 8912 3782 8942 3834
rect 8966 3782 8976 3834
rect 8976 3782 9022 3834
rect 9046 3782 9092 3834
rect 9092 3782 9102 3834
rect 9126 3782 9156 3834
rect 9156 3782 9182 3834
rect 8886 3780 8942 3782
rect 8966 3780 9022 3782
rect 9046 3780 9102 3782
rect 9126 3780 9182 3782
rect 9494 26036 9550 26072
rect 9494 26016 9496 26036
rect 9496 26016 9548 26036
rect 9548 26016 9550 26036
rect 9494 24656 9550 24712
rect 9678 26832 9734 26888
rect 9770 24112 9826 24168
rect 9678 24012 9680 24032
rect 9680 24012 9732 24032
rect 9732 24012 9734 24032
rect 9678 23976 9734 24012
rect 9678 23704 9734 23760
rect 9494 21936 9550 21992
rect 9402 13096 9458 13152
rect 9586 21528 9642 21584
rect 10138 24384 10194 24440
rect 10138 24112 10194 24168
rect 9954 19080 10010 19136
rect 10138 16652 10194 16688
rect 10138 16632 10140 16652
rect 10140 16632 10192 16652
rect 10192 16632 10194 16652
rect 8886 2746 8942 2748
rect 8966 2746 9022 2748
rect 9046 2746 9102 2748
rect 9126 2746 9182 2748
rect 8886 2694 8912 2746
rect 8912 2694 8942 2746
rect 8966 2694 8976 2746
rect 8976 2694 9022 2746
rect 9046 2694 9092 2746
rect 9092 2694 9102 2746
rect 9126 2694 9156 2746
rect 9156 2694 9182 2746
rect 8886 2692 8942 2694
rect 8966 2692 9022 2694
rect 9046 2692 9102 2694
rect 9126 2692 9182 2694
rect 9310 3168 9366 3224
rect 10414 8336 10470 8392
rect 10782 26968 10838 27024
rect 12852 46810 12908 46812
rect 12932 46810 12988 46812
rect 13012 46810 13068 46812
rect 13092 46810 13148 46812
rect 12852 46758 12878 46810
rect 12878 46758 12908 46810
rect 12932 46758 12942 46810
rect 12942 46758 12988 46810
rect 13012 46758 13058 46810
rect 13058 46758 13068 46810
rect 13092 46758 13122 46810
rect 13122 46758 13148 46810
rect 12852 46756 12908 46758
rect 12932 46756 12988 46758
rect 13012 46756 13068 46758
rect 13092 46756 13148 46758
rect 12852 45722 12908 45724
rect 12932 45722 12988 45724
rect 13012 45722 13068 45724
rect 13092 45722 13148 45724
rect 12852 45670 12878 45722
rect 12878 45670 12908 45722
rect 12932 45670 12942 45722
rect 12942 45670 12988 45722
rect 13012 45670 13058 45722
rect 13058 45670 13068 45722
rect 13092 45670 13122 45722
rect 13122 45670 13148 45722
rect 12852 45668 12908 45670
rect 12932 45668 12988 45670
rect 13012 45668 13068 45670
rect 13092 45668 13148 45670
rect 11334 38836 11336 38856
rect 11336 38836 11388 38856
rect 11388 38836 11390 38856
rect 11334 38800 11390 38836
rect 10690 24268 10746 24304
rect 10690 24248 10692 24268
rect 10692 24248 10744 24268
rect 10744 24248 10746 24268
rect 12852 44634 12908 44636
rect 12932 44634 12988 44636
rect 13012 44634 13068 44636
rect 13092 44634 13148 44636
rect 12852 44582 12878 44634
rect 12878 44582 12908 44634
rect 12932 44582 12942 44634
rect 12942 44582 12988 44634
rect 13012 44582 13058 44634
rect 13058 44582 13068 44634
rect 13092 44582 13122 44634
rect 13122 44582 13148 44634
rect 12852 44580 12908 44582
rect 12932 44580 12988 44582
rect 13012 44580 13068 44582
rect 13092 44580 13148 44582
rect 12852 43546 12908 43548
rect 12932 43546 12988 43548
rect 13012 43546 13068 43548
rect 13092 43546 13148 43548
rect 12852 43494 12878 43546
rect 12878 43494 12908 43546
rect 12932 43494 12942 43546
rect 12942 43494 12988 43546
rect 13012 43494 13058 43546
rect 13058 43494 13068 43546
rect 13092 43494 13122 43546
rect 13122 43494 13148 43546
rect 12852 43492 12908 43494
rect 12932 43492 12988 43494
rect 13012 43492 13068 43494
rect 13092 43492 13148 43494
rect 12852 42458 12908 42460
rect 12932 42458 12988 42460
rect 13012 42458 13068 42460
rect 13092 42458 13148 42460
rect 12852 42406 12878 42458
rect 12878 42406 12908 42458
rect 12932 42406 12942 42458
rect 12942 42406 12988 42458
rect 13012 42406 13058 42458
rect 13058 42406 13068 42458
rect 13092 42406 13122 42458
rect 13122 42406 13148 42458
rect 12852 42404 12908 42406
rect 12932 42404 12988 42406
rect 13012 42404 13068 42406
rect 13092 42404 13148 42406
rect 12852 41370 12908 41372
rect 12932 41370 12988 41372
rect 13012 41370 13068 41372
rect 13092 41370 13148 41372
rect 12852 41318 12878 41370
rect 12878 41318 12908 41370
rect 12932 41318 12942 41370
rect 12942 41318 12988 41370
rect 13012 41318 13058 41370
rect 13058 41318 13068 41370
rect 13092 41318 13122 41370
rect 13122 41318 13148 41370
rect 12852 41316 12908 41318
rect 12932 41316 12988 41318
rect 13012 41316 13068 41318
rect 13092 41316 13148 41318
rect 12852 40282 12908 40284
rect 12932 40282 12988 40284
rect 13012 40282 13068 40284
rect 13092 40282 13148 40284
rect 12852 40230 12878 40282
rect 12878 40230 12908 40282
rect 12932 40230 12942 40282
rect 12942 40230 12988 40282
rect 13012 40230 13058 40282
rect 13058 40230 13068 40282
rect 13092 40230 13122 40282
rect 13122 40230 13148 40282
rect 12852 40228 12908 40230
rect 12932 40228 12988 40230
rect 13012 40228 13068 40230
rect 13092 40228 13148 40230
rect 12070 38972 12072 38992
rect 12072 38972 12124 38992
rect 12124 38972 12126 38992
rect 12070 38936 12126 38972
rect 12852 39194 12908 39196
rect 12932 39194 12988 39196
rect 13012 39194 13068 39196
rect 13092 39194 13148 39196
rect 12852 39142 12878 39194
rect 12878 39142 12908 39194
rect 12932 39142 12942 39194
rect 12942 39142 12988 39194
rect 13012 39142 13058 39194
rect 13058 39142 13068 39194
rect 13092 39142 13122 39194
rect 13122 39142 13148 39194
rect 12852 39140 12908 39142
rect 12932 39140 12988 39142
rect 13012 39140 13068 39142
rect 13092 39140 13148 39142
rect 12852 38106 12908 38108
rect 12932 38106 12988 38108
rect 13012 38106 13068 38108
rect 13092 38106 13148 38108
rect 12852 38054 12878 38106
rect 12878 38054 12908 38106
rect 12932 38054 12942 38106
rect 12942 38054 12988 38106
rect 13012 38054 13058 38106
rect 13058 38054 13068 38106
rect 13092 38054 13122 38106
rect 13122 38054 13148 38106
rect 12852 38052 12908 38054
rect 12932 38052 12988 38054
rect 13012 38052 13068 38054
rect 13092 38052 13148 38054
rect 11242 23296 11298 23352
rect 11426 24384 11482 24440
rect 11426 23024 11482 23080
rect 11150 21564 11152 21584
rect 11152 21564 11204 21584
rect 11204 21564 11206 21584
rect 11150 21528 11206 21564
rect 11150 21428 11152 21448
rect 11152 21428 11204 21448
rect 11204 21428 11206 21448
rect 11150 21392 11206 21428
rect 11334 22072 11390 22128
rect 10782 9152 10838 9208
rect 12852 37018 12908 37020
rect 12932 37018 12988 37020
rect 13012 37018 13068 37020
rect 13092 37018 13148 37020
rect 12852 36966 12878 37018
rect 12878 36966 12908 37018
rect 12932 36966 12942 37018
rect 12942 36966 12988 37018
rect 13012 36966 13058 37018
rect 13058 36966 13068 37018
rect 13092 36966 13122 37018
rect 13122 36966 13148 37018
rect 12852 36964 12908 36966
rect 12932 36964 12988 36966
rect 13012 36964 13068 36966
rect 13092 36964 13148 36966
rect 12852 35930 12908 35932
rect 12932 35930 12988 35932
rect 13012 35930 13068 35932
rect 13092 35930 13148 35932
rect 12852 35878 12878 35930
rect 12878 35878 12908 35930
rect 12932 35878 12942 35930
rect 12942 35878 12988 35930
rect 13012 35878 13058 35930
rect 13058 35878 13068 35930
rect 13092 35878 13122 35930
rect 13122 35878 13148 35930
rect 12852 35876 12908 35878
rect 12932 35876 12988 35878
rect 13012 35876 13068 35878
rect 13092 35876 13148 35878
rect 12852 34842 12908 34844
rect 12932 34842 12988 34844
rect 13012 34842 13068 34844
rect 13092 34842 13148 34844
rect 12852 34790 12878 34842
rect 12878 34790 12908 34842
rect 12932 34790 12942 34842
rect 12942 34790 12988 34842
rect 13012 34790 13058 34842
rect 13058 34790 13068 34842
rect 13092 34790 13122 34842
rect 13122 34790 13148 34842
rect 12852 34788 12908 34790
rect 12932 34788 12988 34790
rect 13012 34788 13068 34790
rect 13092 34788 13148 34790
rect 12852 33754 12908 33756
rect 12932 33754 12988 33756
rect 13012 33754 13068 33756
rect 13092 33754 13148 33756
rect 12852 33702 12878 33754
rect 12878 33702 12908 33754
rect 12932 33702 12942 33754
rect 12942 33702 12988 33754
rect 13012 33702 13058 33754
rect 13058 33702 13068 33754
rect 13092 33702 13122 33754
rect 13122 33702 13148 33754
rect 12852 33700 12908 33702
rect 12932 33700 12988 33702
rect 13012 33700 13068 33702
rect 13092 33700 13148 33702
rect 12852 32666 12908 32668
rect 12932 32666 12988 32668
rect 13012 32666 13068 32668
rect 13092 32666 13148 32668
rect 12852 32614 12878 32666
rect 12878 32614 12908 32666
rect 12932 32614 12942 32666
rect 12942 32614 12988 32666
rect 13012 32614 13058 32666
rect 13058 32614 13068 32666
rect 13092 32614 13122 32666
rect 13122 32614 13148 32666
rect 12852 32612 12908 32614
rect 12932 32612 12988 32614
rect 13012 32612 13068 32614
rect 13092 32612 13148 32614
rect 12852 31578 12908 31580
rect 12932 31578 12988 31580
rect 13012 31578 13068 31580
rect 13092 31578 13148 31580
rect 12852 31526 12878 31578
rect 12878 31526 12908 31578
rect 12932 31526 12942 31578
rect 12942 31526 12988 31578
rect 13012 31526 13058 31578
rect 13058 31526 13068 31578
rect 13092 31526 13122 31578
rect 13122 31526 13148 31578
rect 12852 31524 12908 31526
rect 12932 31524 12988 31526
rect 13012 31524 13068 31526
rect 13092 31524 13148 31526
rect 12852 30490 12908 30492
rect 12932 30490 12988 30492
rect 13012 30490 13068 30492
rect 13092 30490 13148 30492
rect 12852 30438 12878 30490
rect 12878 30438 12908 30490
rect 12932 30438 12942 30490
rect 12942 30438 12988 30490
rect 13012 30438 13058 30490
rect 13058 30438 13068 30490
rect 13092 30438 13122 30490
rect 13122 30438 13148 30490
rect 12852 30436 12908 30438
rect 12932 30436 12988 30438
rect 13012 30436 13068 30438
rect 13092 30436 13148 30438
rect 12852 29402 12908 29404
rect 12932 29402 12988 29404
rect 13012 29402 13068 29404
rect 13092 29402 13148 29404
rect 12852 29350 12878 29402
rect 12878 29350 12908 29402
rect 12932 29350 12942 29402
rect 12942 29350 12988 29402
rect 13012 29350 13058 29402
rect 13058 29350 13068 29402
rect 13092 29350 13122 29402
rect 13122 29350 13148 29402
rect 12852 29348 12908 29350
rect 12932 29348 12988 29350
rect 13012 29348 13068 29350
rect 13092 29348 13148 29350
rect 11886 23196 11888 23216
rect 11888 23196 11940 23216
rect 11940 23196 11942 23216
rect 11886 23160 11942 23196
rect 12070 23160 12126 23216
rect 10966 9596 10968 9616
rect 10968 9596 11020 9616
rect 11020 9596 11022 9616
rect 10966 9560 11022 9596
rect 10966 9424 11022 9480
rect 10966 8880 11022 8936
rect 10966 7928 11022 7984
rect 11518 9288 11574 9344
rect 12438 23704 12494 23760
rect 12254 23316 12310 23352
rect 12254 23296 12256 23316
rect 12256 23296 12308 23316
rect 12308 23296 12310 23316
rect 12254 23024 12310 23080
rect 12852 28314 12908 28316
rect 12932 28314 12988 28316
rect 13012 28314 13068 28316
rect 13092 28314 13148 28316
rect 12852 28262 12878 28314
rect 12878 28262 12908 28314
rect 12932 28262 12942 28314
rect 12942 28262 12988 28314
rect 13012 28262 13058 28314
rect 13058 28262 13068 28314
rect 13092 28262 13122 28314
rect 13122 28262 13148 28314
rect 12852 28260 12908 28262
rect 12932 28260 12988 28262
rect 13012 28260 13068 28262
rect 13092 28260 13148 28262
rect 14094 38800 14150 38856
rect 12852 27226 12908 27228
rect 12932 27226 12988 27228
rect 13012 27226 13068 27228
rect 13092 27226 13148 27228
rect 12852 27174 12878 27226
rect 12878 27174 12908 27226
rect 12932 27174 12942 27226
rect 12942 27174 12988 27226
rect 13012 27174 13058 27226
rect 13058 27174 13068 27226
rect 13092 27174 13122 27226
rect 13122 27174 13148 27226
rect 12852 27172 12908 27174
rect 12932 27172 12988 27174
rect 13012 27172 13068 27174
rect 13092 27172 13148 27174
rect 12622 24692 12624 24712
rect 12624 24692 12676 24712
rect 12676 24692 12678 24712
rect 12852 26138 12908 26140
rect 12932 26138 12988 26140
rect 13012 26138 13068 26140
rect 13092 26138 13148 26140
rect 12852 26086 12878 26138
rect 12878 26086 12908 26138
rect 12932 26086 12942 26138
rect 12942 26086 12988 26138
rect 13012 26086 13058 26138
rect 13058 26086 13068 26138
rect 13092 26086 13122 26138
rect 13122 26086 13148 26138
rect 12852 26084 12908 26086
rect 12932 26084 12988 26086
rect 13012 26084 13068 26086
rect 13092 26084 13148 26086
rect 12852 25050 12908 25052
rect 12932 25050 12988 25052
rect 13012 25050 13068 25052
rect 13092 25050 13148 25052
rect 12852 24998 12878 25050
rect 12878 24998 12908 25050
rect 12932 24998 12942 25050
rect 12942 24998 12988 25050
rect 13012 24998 13058 25050
rect 13058 24998 13068 25050
rect 13092 24998 13122 25050
rect 13122 24998 13148 25050
rect 12852 24996 12908 24998
rect 12932 24996 12988 24998
rect 13012 24996 13068 24998
rect 13092 24996 13148 24998
rect 12622 24656 12678 24692
rect 12622 23976 12678 24032
rect 12530 23160 12586 23216
rect 12852 23962 12908 23964
rect 12932 23962 12988 23964
rect 13012 23962 13068 23964
rect 13092 23962 13148 23964
rect 12852 23910 12878 23962
rect 12878 23910 12908 23962
rect 12932 23910 12942 23962
rect 12942 23910 12988 23962
rect 13012 23910 13058 23962
rect 13058 23910 13068 23962
rect 13092 23910 13122 23962
rect 13122 23910 13148 23962
rect 12852 23908 12908 23910
rect 12932 23908 12988 23910
rect 13012 23908 13068 23910
rect 13092 23908 13148 23910
rect 12852 22874 12908 22876
rect 12932 22874 12988 22876
rect 13012 22874 13068 22876
rect 13092 22874 13148 22876
rect 12852 22822 12878 22874
rect 12878 22822 12908 22874
rect 12932 22822 12942 22874
rect 12942 22822 12988 22874
rect 13012 22822 13058 22874
rect 13058 22822 13068 22874
rect 13092 22822 13122 22874
rect 13122 22822 13148 22874
rect 12852 22820 12908 22822
rect 12932 22820 12988 22822
rect 13012 22820 13068 22822
rect 13092 22820 13148 22822
rect 12852 21786 12908 21788
rect 12932 21786 12988 21788
rect 13012 21786 13068 21788
rect 13092 21786 13148 21788
rect 12852 21734 12878 21786
rect 12878 21734 12908 21786
rect 12932 21734 12942 21786
rect 12942 21734 12988 21786
rect 13012 21734 13058 21786
rect 13058 21734 13068 21786
rect 13092 21734 13122 21786
rect 13122 21734 13148 21786
rect 12852 21732 12908 21734
rect 12932 21732 12988 21734
rect 13012 21732 13068 21734
rect 13092 21732 13148 21734
rect 12852 20698 12908 20700
rect 12932 20698 12988 20700
rect 13012 20698 13068 20700
rect 13092 20698 13148 20700
rect 12852 20646 12878 20698
rect 12878 20646 12908 20698
rect 12932 20646 12942 20698
rect 12942 20646 12988 20698
rect 13012 20646 13058 20698
rect 13058 20646 13068 20698
rect 13092 20646 13122 20698
rect 13122 20646 13148 20698
rect 12852 20644 12908 20646
rect 12932 20644 12988 20646
rect 13012 20644 13068 20646
rect 13092 20644 13148 20646
rect 12852 19610 12908 19612
rect 12932 19610 12988 19612
rect 13012 19610 13068 19612
rect 13092 19610 13148 19612
rect 12852 19558 12878 19610
rect 12878 19558 12908 19610
rect 12932 19558 12942 19610
rect 12942 19558 12988 19610
rect 13012 19558 13058 19610
rect 13058 19558 13068 19610
rect 13092 19558 13122 19610
rect 13122 19558 13148 19610
rect 12852 19556 12908 19558
rect 12932 19556 12988 19558
rect 13012 19556 13068 19558
rect 13092 19556 13148 19558
rect 12852 18522 12908 18524
rect 12932 18522 12988 18524
rect 13012 18522 13068 18524
rect 13092 18522 13148 18524
rect 12852 18470 12878 18522
rect 12878 18470 12908 18522
rect 12932 18470 12942 18522
rect 12942 18470 12988 18522
rect 13012 18470 13058 18522
rect 13058 18470 13068 18522
rect 13092 18470 13122 18522
rect 13122 18470 13148 18522
rect 12852 18468 12908 18470
rect 12932 18468 12988 18470
rect 13012 18468 13068 18470
rect 13092 18468 13148 18470
rect 14094 21392 14150 21448
rect 12852 17434 12908 17436
rect 12932 17434 12988 17436
rect 13012 17434 13068 17436
rect 13092 17434 13148 17436
rect 12852 17382 12878 17434
rect 12878 17382 12908 17434
rect 12932 17382 12942 17434
rect 12942 17382 12988 17434
rect 13012 17382 13058 17434
rect 13058 17382 13068 17434
rect 13092 17382 13122 17434
rect 13122 17382 13148 17434
rect 12852 17380 12908 17382
rect 12932 17380 12988 17382
rect 13012 17380 13068 17382
rect 13092 17380 13148 17382
rect 12852 16346 12908 16348
rect 12932 16346 12988 16348
rect 13012 16346 13068 16348
rect 13092 16346 13148 16348
rect 12852 16294 12878 16346
rect 12878 16294 12908 16346
rect 12932 16294 12942 16346
rect 12942 16294 12988 16346
rect 13012 16294 13058 16346
rect 13058 16294 13068 16346
rect 13092 16294 13122 16346
rect 13122 16294 13148 16346
rect 12852 16292 12908 16294
rect 12932 16292 12988 16294
rect 13012 16292 13068 16294
rect 13092 16292 13148 16294
rect 12438 10920 12494 10976
rect 12346 10648 12402 10704
rect 12852 15258 12908 15260
rect 12932 15258 12988 15260
rect 13012 15258 13068 15260
rect 13092 15258 13148 15260
rect 12852 15206 12878 15258
rect 12878 15206 12908 15258
rect 12932 15206 12942 15258
rect 12942 15206 12988 15258
rect 13012 15206 13058 15258
rect 13058 15206 13068 15258
rect 13092 15206 13122 15258
rect 13122 15206 13148 15258
rect 12852 15204 12908 15206
rect 12932 15204 12988 15206
rect 13012 15204 13068 15206
rect 13092 15204 13148 15206
rect 12852 14170 12908 14172
rect 12932 14170 12988 14172
rect 13012 14170 13068 14172
rect 13092 14170 13148 14172
rect 12852 14118 12878 14170
rect 12878 14118 12908 14170
rect 12932 14118 12942 14170
rect 12942 14118 12988 14170
rect 13012 14118 13058 14170
rect 13058 14118 13068 14170
rect 13092 14118 13122 14170
rect 13122 14118 13148 14170
rect 12852 14116 12908 14118
rect 12932 14116 12988 14118
rect 13012 14116 13068 14118
rect 13092 14116 13148 14118
rect 12852 13082 12908 13084
rect 12932 13082 12988 13084
rect 13012 13082 13068 13084
rect 13092 13082 13148 13084
rect 12852 13030 12878 13082
rect 12878 13030 12908 13082
rect 12932 13030 12942 13082
rect 12942 13030 12988 13082
rect 13012 13030 13058 13082
rect 13058 13030 13068 13082
rect 13092 13030 13122 13082
rect 13122 13030 13148 13082
rect 12852 13028 12908 13030
rect 12932 13028 12988 13030
rect 13012 13028 13068 13030
rect 13092 13028 13148 13030
rect 12852 11994 12908 11996
rect 12932 11994 12988 11996
rect 13012 11994 13068 11996
rect 13092 11994 13148 11996
rect 12852 11942 12878 11994
rect 12878 11942 12908 11994
rect 12932 11942 12942 11994
rect 12942 11942 12988 11994
rect 13012 11942 13058 11994
rect 13058 11942 13068 11994
rect 13092 11942 13122 11994
rect 13122 11942 13148 11994
rect 12852 11940 12908 11942
rect 12932 11940 12988 11942
rect 13012 11940 13068 11942
rect 13092 11940 13148 11942
rect 12714 11192 12770 11248
rect 12438 9832 12494 9888
rect 12438 9052 12440 9072
rect 12440 9052 12492 9072
rect 12492 9052 12494 9072
rect 12438 9016 12494 9052
rect 12254 8880 12310 8936
rect 12162 7792 12218 7848
rect 12438 8336 12494 8392
rect 12162 4392 12218 4448
rect 12852 10906 12908 10908
rect 12932 10906 12988 10908
rect 13012 10906 13068 10908
rect 13092 10906 13148 10908
rect 12852 10854 12878 10906
rect 12878 10854 12908 10906
rect 12932 10854 12942 10906
rect 12942 10854 12988 10906
rect 13012 10854 13058 10906
rect 13058 10854 13068 10906
rect 13092 10854 13122 10906
rect 13122 10854 13148 10906
rect 12852 10852 12908 10854
rect 12932 10852 12988 10854
rect 13012 10852 13068 10854
rect 13092 10852 13148 10854
rect 12852 9818 12908 9820
rect 12932 9818 12988 9820
rect 13012 9818 13068 9820
rect 13092 9818 13148 9820
rect 12852 9766 12878 9818
rect 12878 9766 12908 9818
rect 12932 9766 12942 9818
rect 12942 9766 12988 9818
rect 13012 9766 13058 9818
rect 13058 9766 13068 9818
rect 13092 9766 13122 9818
rect 13122 9766 13148 9818
rect 12852 9764 12908 9766
rect 12932 9764 12988 9766
rect 13012 9764 13068 9766
rect 13092 9764 13148 9766
rect 12898 9288 12954 9344
rect 12852 8730 12908 8732
rect 12932 8730 12988 8732
rect 13012 8730 13068 8732
rect 13092 8730 13148 8732
rect 12852 8678 12878 8730
rect 12878 8678 12908 8730
rect 12932 8678 12942 8730
rect 12942 8678 12988 8730
rect 13012 8678 13058 8730
rect 13058 8678 13068 8730
rect 13092 8678 13122 8730
rect 13122 8678 13148 8730
rect 12852 8676 12908 8678
rect 12932 8676 12988 8678
rect 13012 8676 13068 8678
rect 13092 8676 13148 8678
rect 13082 8336 13138 8392
rect 12898 8064 12954 8120
rect 13174 8200 13230 8256
rect 12852 7642 12908 7644
rect 12932 7642 12988 7644
rect 13012 7642 13068 7644
rect 13092 7642 13148 7644
rect 12852 7590 12878 7642
rect 12878 7590 12908 7642
rect 12932 7590 12942 7642
rect 12942 7590 12988 7642
rect 13012 7590 13058 7642
rect 13058 7590 13068 7642
rect 13092 7590 13122 7642
rect 13122 7590 13148 7642
rect 12852 7588 12908 7590
rect 12932 7588 12988 7590
rect 13012 7588 13068 7590
rect 13092 7588 13148 7590
rect 13450 8064 13506 8120
rect 12852 6554 12908 6556
rect 12932 6554 12988 6556
rect 13012 6554 13068 6556
rect 13092 6554 13148 6556
rect 12852 6502 12878 6554
rect 12878 6502 12908 6554
rect 12932 6502 12942 6554
rect 12942 6502 12988 6554
rect 13012 6502 13058 6554
rect 13058 6502 13068 6554
rect 13092 6502 13122 6554
rect 13122 6502 13148 6554
rect 12852 6500 12908 6502
rect 12932 6500 12988 6502
rect 13012 6500 13068 6502
rect 13092 6500 13148 6502
rect 12852 5466 12908 5468
rect 12932 5466 12988 5468
rect 13012 5466 13068 5468
rect 13092 5466 13148 5468
rect 12852 5414 12878 5466
rect 12878 5414 12908 5466
rect 12932 5414 12942 5466
rect 12942 5414 12988 5466
rect 13012 5414 13058 5466
rect 13058 5414 13068 5466
rect 13092 5414 13122 5466
rect 13122 5414 13148 5466
rect 12852 5412 12908 5414
rect 12932 5412 12988 5414
rect 13012 5412 13068 5414
rect 13092 5412 13148 5414
rect 12852 4378 12908 4380
rect 12932 4378 12988 4380
rect 13012 4378 13068 4380
rect 13092 4378 13148 4380
rect 12852 4326 12878 4378
rect 12878 4326 12908 4378
rect 12932 4326 12942 4378
rect 12942 4326 12988 4378
rect 13012 4326 13058 4378
rect 13058 4326 13068 4378
rect 13092 4326 13122 4378
rect 13122 4326 13148 4378
rect 12852 4324 12908 4326
rect 12932 4324 12988 4326
rect 13012 4324 13068 4326
rect 13092 4324 13148 4326
rect 12852 3290 12908 3292
rect 12932 3290 12988 3292
rect 13012 3290 13068 3292
rect 13092 3290 13148 3292
rect 12852 3238 12878 3290
rect 12878 3238 12908 3290
rect 12932 3238 12942 3290
rect 12942 3238 12988 3290
rect 13012 3238 13058 3290
rect 13058 3238 13068 3290
rect 13092 3238 13122 3290
rect 13122 3238 13148 3290
rect 12852 3236 12908 3238
rect 12932 3236 12988 3238
rect 13012 3236 13068 3238
rect 13092 3236 13148 3238
rect 12852 2202 12908 2204
rect 12932 2202 12988 2204
rect 13012 2202 13068 2204
rect 13092 2202 13148 2204
rect 12852 2150 12878 2202
rect 12878 2150 12908 2202
rect 12932 2150 12942 2202
rect 12942 2150 12988 2202
rect 13012 2150 13058 2202
rect 13058 2150 13068 2202
rect 13092 2150 13122 2202
rect 13122 2150 13148 2202
rect 12852 2148 12908 2150
rect 12932 2148 12988 2150
rect 13012 2148 13068 2150
rect 13092 2148 13148 2150
rect 16817 47354 16873 47356
rect 16897 47354 16953 47356
rect 16977 47354 17033 47356
rect 17057 47354 17113 47356
rect 16817 47302 16843 47354
rect 16843 47302 16873 47354
rect 16897 47302 16907 47354
rect 16907 47302 16953 47354
rect 16977 47302 17023 47354
rect 17023 47302 17033 47354
rect 17057 47302 17087 47354
rect 17087 47302 17113 47354
rect 16817 47300 16873 47302
rect 16897 47300 16953 47302
rect 16977 47300 17033 47302
rect 17057 47300 17113 47302
rect 16817 46266 16873 46268
rect 16897 46266 16953 46268
rect 16977 46266 17033 46268
rect 17057 46266 17113 46268
rect 16817 46214 16843 46266
rect 16843 46214 16873 46266
rect 16897 46214 16907 46266
rect 16907 46214 16953 46266
rect 16977 46214 17023 46266
rect 17023 46214 17033 46266
rect 17057 46214 17087 46266
rect 17087 46214 17113 46266
rect 16817 46212 16873 46214
rect 16897 46212 16953 46214
rect 16977 46212 17033 46214
rect 17057 46212 17113 46214
rect 16817 45178 16873 45180
rect 16897 45178 16953 45180
rect 16977 45178 17033 45180
rect 17057 45178 17113 45180
rect 16817 45126 16843 45178
rect 16843 45126 16873 45178
rect 16897 45126 16907 45178
rect 16907 45126 16953 45178
rect 16977 45126 17023 45178
rect 17023 45126 17033 45178
rect 17057 45126 17087 45178
rect 17087 45126 17113 45178
rect 16817 45124 16873 45126
rect 16897 45124 16953 45126
rect 16977 45124 17033 45126
rect 17057 45124 17113 45126
rect 16817 44090 16873 44092
rect 16897 44090 16953 44092
rect 16977 44090 17033 44092
rect 17057 44090 17113 44092
rect 16817 44038 16843 44090
rect 16843 44038 16873 44090
rect 16897 44038 16907 44090
rect 16907 44038 16953 44090
rect 16977 44038 17023 44090
rect 17023 44038 17033 44090
rect 17057 44038 17087 44090
rect 17087 44038 17113 44090
rect 16817 44036 16873 44038
rect 16897 44036 16953 44038
rect 16977 44036 17033 44038
rect 17057 44036 17113 44038
rect 16817 43002 16873 43004
rect 16897 43002 16953 43004
rect 16977 43002 17033 43004
rect 17057 43002 17113 43004
rect 16817 42950 16843 43002
rect 16843 42950 16873 43002
rect 16897 42950 16907 43002
rect 16907 42950 16953 43002
rect 16977 42950 17023 43002
rect 17023 42950 17033 43002
rect 17057 42950 17087 43002
rect 17087 42950 17113 43002
rect 16817 42948 16873 42950
rect 16897 42948 16953 42950
rect 16977 42948 17033 42950
rect 17057 42948 17113 42950
rect 16817 41914 16873 41916
rect 16897 41914 16953 41916
rect 16977 41914 17033 41916
rect 17057 41914 17113 41916
rect 16817 41862 16843 41914
rect 16843 41862 16873 41914
rect 16897 41862 16907 41914
rect 16907 41862 16953 41914
rect 16977 41862 17023 41914
rect 17023 41862 17033 41914
rect 17057 41862 17087 41914
rect 17087 41862 17113 41914
rect 16817 41860 16873 41862
rect 16897 41860 16953 41862
rect 16977 41860 17033 41862
rect 17057 41860 17113 41862
rect 16817 40826 16873 40828
rect 16897 40826 16953 40828
rect 16977 40826 17033 40828
rect 17057 40826 17113 40828
rect 16817 40774 16843 40826
rect 16843 40774 16873 40826
rect 16897 40774 16907 40826
rect 16907 40774 16953 40826
rect 16977 40774 17023 40826
rect 17023 40774 17033 40826
rect 17057 40774 17087 40826
rect 17087 40774 17113 40826
rect 16817 40772 16873 40774
rect 16897 40772 16953 40774
rect 16977 40772 17033 40774
rect 17057 40772 17113 40774
rect 14646 23568 14702 23624
rect 13634 4120 13690 4176
rect 14738 9152 14794 9208
rect 14370 7948 14426 7984
rect 14370 7928 14372 7948
rect 14372 7928 14424 7948
rect 14424 7928 14426 7948
rect 14462 7828 14464 7848
rect 14464 7828 14516 7848
rect 14516 7828 14518 7848
rect 14462 7792 14518 7828
rect 16817 39738 16873 39740
rect 16897 39738 16953 39740
rect 16977 39738 17033 39740
rect 17057 39738 17113 39740
rect 16817 39686 16843 39738
rect 16843 39686 16873 39738
rect 16897 39686 16907 39738
rect 16907 39686 16953 39738
rect 16977 39686 17023 39738
rect 17023 39686 17033 39738
rect 17057 39686 17087 39738
rect 17087 39686 17113 39738
rect 16817 39684 16873 39686
rect 16897 39684 16953 39686
rect 16977 39684 17033 39686
rect 17057 39684 17113 39686
rect 16670 38936 16726 38992
rect 16817 38650 16873 38652
rect 16897 38650 16953 38652
rect 16977 38650 17033 38652
rect 17057 38650 17113 38652
rect 16817 38598 16843 38650
rect 16843 38598 16873 38650
rect 16897 38598 16907 38650
rect 16907 38598 16953 38650
rect 16977 38598 17023 38650
rect 17023 38598 17033 38650
rect 17057 38598 17087 38650
rect 17087 38598 17113 38650
rect 16817 38596 16873 38598
rect 16897 38596 16953 38598
rect 16977 38596 17033 38598
rect 17057 38596 17113 38598
rect 16817 37562 16873 37564
rect 16897 37562 16953 37564
rect 16977 37562 17033 37564
rect 17057 37562 17113 37564
rect 16817 37510 16843 37562
rect 16843 37510 16873 37562
rect 16897 37510 16907 37562
rect 16907 37510 16953 37562
rect 16977 37510 17023 37562
rect 17023 37510 17033 37562
rect 17057 37510 17087 37562
rect 17087 37510 17113 37562
rect 16817 37508 16873 37510
rect 16897 37508 16953 37510
rect 16977 37508 17033 37510
rect 17057 37508 17113 37510
rect 16817 36474 16873 36476
rect 16897 36474 16953 36476
rect 16977 36474 17033 36476
rect 17057 36474 17113 36476
rect 16817 36422 16843 36474
rect 16843 36422 16873 36474
rect 16897 36422 16907 36474
rect 16907 36422 16953 36474
rect 16977 36422 17023 36474
rect 17023 36422 17033 36474
rect 17057 36422 17087 36474
rect 17087 36422 17113 36474
rect 16817 36420 16873 36422
rect 16897 36420 16953 36422
rect 16977 36420 17033 36422
rect 17057 36420 17113 36422
rect 15566 16632 15622 16688
rect 16817 35386 16873 35388
rect 16897 35386 16953 35388
rect 16977 35386 17033 35388
rect 17057 35386 17113 35388
rect 16817 35334 16843 35386
rect 16843 35334 16873 35386
rect 16897 35334 16907 35386
rect 16907 35334 16953 35386
rect 16977 35334 17023 35386
rect 17023 35334 17033 35386
rect 17057 35334 17087 35386
rect 17087 35334 17113 35386
rect 16817 35332 16873 35334
rect 16897 35332 16953 35334
rect 16977 35332 17033 35334
rect 17057 35332 17113 35334
rect 20782 46810 20838 46812
rect 20862 46810 20918 46812
rect 20942 46810 20998 46812
rect 21022 46810 21078 46812
rect 20782 46758 20808 46810
rect 20808 46758 20838 46810
rect 20862 46758 20872 46810
rect 20872 46758 20918 46810
rect 20942 46758 20988 46810
rect 20988 46758 20998 46810
rect 21022 46758 21052 46810
rect 21052 46758 21078 46810
rect 20782 46756 20838 46758
rect 20862 46756 20918 46758
rect 20942 46756 20998 46758
rect 21022 46756 21078 46758
rect 20782 45722 20838 45724
rect 20862 45722 20918 45724
rect 20942 45722 20998 45724
rect 21022 45722 21078 45724
rect 20782 45670 20808 45722
rect 20808 45670 20838 45722
rect 20862 45670 20872 45722
rect 20872 45670 20918 45722
rect 20942 45670 20988 45722
rect 20988 45670 20998 45722
rect 21022 45670 21052 45722
rect 21052 45670 21078 45722
rect 20782 45668 20838 45670
rect 20862 45668 20918 45670
rect 20942 45668 20998 45670
rect 21022 45668 21078 45670
rect 20782 44634 20838 44636
rect 20862 44634 20918 44636
rect 20942 44634 20998 44636
rect 21022 44634 21078 44636
rect 20782 44582 20808 44634
rect 20808 44582 20838 44634
rect 20862 44582 20872 44634
rect 20872 44582 20918 44634
rect 20942 44582 20988 44634
rect 20988 44582 20998 44634
rect 21022 44582 21052 44634
rect 21052 44582 21078 44634
rect 20782 44580 20838 44582
rect 20862 44580 20918 44582
rect 20942 44580 20998 44582
rect 21022 44580 21078 44582
rect 20782 43546 20838 43548
rect 20862 43546 20918 43548
rect 20942 43546 20998 43548
rect 21022 43546 21078 43548
rect 20782 43494 20808 43546
rect 20808 43494 20838 43546
rect 20862 43494 20872 43546
rect 20872 43494 20918 43546
rect 20942 43494 20988 43546
rect 20988 43494 20998 43546
rect 21022 43494 21052 43546
rect 21052 43494 21078 43546
rect 20782 43492 20838 43494
rect 20862 43492 20918 43494
rect 20942 43492 20998 43494
rect 21022 43492 21078 43494
rect 20782 42458 20838 42460
rect 20862 42458 20918 42460
rect 20942 42458 20998 42460
rect 21022 42458 21078 42460
rect 20782 42406 20808 42458
rect 20808 42406 20838 42458
rect 20862 42406 20872 42458
rect 20872 42406 20918 42458
rect 20942 42406 20988 42458
rect 20988 42406 20998 42458
rect 21022 42406 21052 42458
rect 21052 42406 21078 42458
rect 20782 42404 20838 42406
rect 20862 42404 20918 42406
rect 20942 42404 20998 42406
rect 21022 42404 21078 42406
rect 20782 41370 20838 41372
rect 20862 41370 20918 41372
rect 20942 41370 20998 41372
rect 21022 41370 21078 41372
rect 20782 41318 20808 41370
rect 20808 41318 20838 41370
rect 20862 41318 20872 41370
rect 20872 41318 20918 41370
rect 20942 41318 20988 41370
rect 20988 41318 20998 41370
rect 21022 41318 21052 41370
rect 21052 41318 21078 41370
rect 20782 41316 20838 41318
rect 20862 41316 20918 41318
rect 20942 41316 20998 41318
rect 21022 41316 21078 41318
rect 20782 40282 20838 40284
rect 20862 40282 20918 40284
rect 20942 40282 20998 40284
rect 21022 40282 21078 40284
rect 20782 40230 20808 40282
rect 20808 40230 20838 40282
rect 20862 40230 20872 40282
rect 20872 40230 20918 40282
rect 20942 40230 20988 40282
rect 20988 40230 20998 40282
rect 21022 40230 21052 40282
rect 21052 40230 21078 40282
rect 20782 40228 20838 40230
rect 20862 40228 20918 40230
rect 20942 40228 20998 40230
rect 21022 40228 21078 40230
rect 20782 39194 20838 39196
rect 20862 39194 20918 39196
rect 20942 39194 20998 39196
rect 21022 39194 21078 39196
rect 20782 39142 20808 39194
rect 20808 39142 20838 39194
rect 20862 39142 20872 39194
rect 20872 39142 20918 39194
rect 20942 39142 20988 39194
rect 20988 39142 20998 39194
rect 21022 39142 21052 39194
rect 21052 39142 21078 39194
rect 20782 39140 20838 39142
rect 20862 39140 20918 39142
rect 20942 39140 20998 39142
rect 21022 39140 21078 39142
rect 20782 38106 20838 38108
rect 20862 38106 20918 38108
rect 20942 38106 20998 38108
rect 21022 38106 21078 38108
rect 20782 38054 20808 38106
rect 20808 38054 20838 38106
rect 20862 38054 20872 38106
rect 20872 38054 20918 38106
rect 20942 38054 20988 38106
rect 20988 38054 20998 38106
rect 21022 38054 21052 38106
rect 21052 38054 21078 38106
rect 20782 38052 20838 38054
rect 20862 38052 20918 38054
rect 20942 38052 20998 38054
rect 21022 38052 21078 38054
rect 20782 37018 20838 37020
rect 20862 37018 20918 37020
rect 20942 37018 20998 37020
rect 21022 37018 21078 37020
rect 20782 36966 20808 37018
rect 20808 36966 20838 37018
rect 20862 36966 20872 37018
rect 20872 36966 20918 37018
rect 20942 36966 20988 37018
rect 20988 36966 20998 37018
rect 21022 36966 21052 37018
rect 21052 36966 21078 37018
rect 20782 36964 20838 36966
rect 20862 36964 20918 36966
rect 20942 36964 20998 36966
rect 21022 36964 21078 36966
rect 20782 35930 20838 35932
rect 20862 35930 20918 35932
rect 20942 35930 20998 35932
rect 21022 35930 21078 35932
rect 20782 35878 20808 35930
rect 20808 35878 20838 35930
rect 20862 35878 20872 35930
rect 20872 35878 20918 35930
rect 20942 35878 20988 35930
rect 20988 35878 20998 35930
rect 21022 35878 21052 35930
rect 21052 35878 21078 35930
rect 20782 35876 20838 35878
rect 20862 35876 20918 35878
rect 20942 35876 20998 35878
rect 21022 35876 21078 35878
rect 16817 34298 16873 34300
rect 16897 34298 16953 34300
rect 16977 34298 17033 34300
rect 17057 34298 17113 34300
rect 16817 34246 16843 34298
rect 16843 34246 16873 34298
rect 16897 34246 16907 34298
rect 16907 34246 16953 34298
rect 16977 34246 17023 34298
rect 17023 34246 17033 34298
rect 17057 34246 17087 34298
rect 17087 34246 17113 34298
rect 16817 34244 16873 34246
rect 16897 34244 16953 34246
rect 16977 34244 17033 34246
rect 17057 34244 17113 34246
rect 20782 34842 20838 34844
rect 20862 34842 20918 34844
rect 20942 34842 20998 34844
rect 21022 34842 21078 34844
rect 20782 34790 20808 34842
rect 20808 34790 20838 34842
rect 20862 34790 20872 34842
rect 20872 34790 20918 34842
rect 20942 34790 20988 34842
rect 20988 34790 20998 34842
rect 21022 34790 21052 34842
rect 21052 34790 21078 34842
rect 20782 34788 20838 34790
rect 20862 34788 20918 34790
rect 20942 34788 20998 34790
rect 21022 34788 21078 34790
rect 20782 33754 20838 33756
rect 20862 33754 20918 33756
rect 20942 33754 20998 33756
rect 21022 33754 21078 33756
rect 20782 33702 20808 33754
rect 20808 33702 20838 33754
rect 20862 33702 20872 33754
rect 20872 33702 20918 33754
rect 20942 33702 20988 33754
rect 20988 33702 20998 33754
rect 21022 33702 21052 33754
rect 21052 33702 21078 33754
rect 20782 33700 20838 33702
rect 20862 33700 20918 33702
rect 20942 33700 20998 33702
rect 21022 33700 21078 33702
rect 16817 33210 16873 33212
rect 16897 33210 16953 33212
rect 16977 33210 17033 33212
rect 17057 33210 17113 33212
rect 16817 33158 16843 33210
rect 16843 33158 16873 33210
rect 16897 33158 16907 33210
rect 16907 33158 16953 33210
rect 16977 33158 17023 33210
rect 17023 33158 17033 33210
rect 17057 33158 17087 33210
rect 17087 33158 17113 33210
rect 16817 33156 16873 33158
rect 16897 33156 16953 33158
rect 16977 33156 17033 33158
rect 17057 33156 17113 33158
rect 20782 32666 20838 32668
rect 20862 32666 20918 32668
rect 20942 32666 20998 32668
rect 21022 32666 21078 32668
rect 20782 32614 20808 32666
rect 20808 32614 20838 32666
rect 20862 32614 20872 32666
rect 20872 32614 20918 32666
rect 20942 32614 20988 32666
rect 20988 32614 20998 32666
rect 21022 32614 21052 32666
rect 21052 32614 21078 32666
rect 20782 32612 20838 32614
rect 20862 32612 20918 32614
rect 20942 32612 20998 32614
rect 21022 32612 21078 32614
rect 16817 32122 16873 32124
rect 16897 32122 16953 32124
rect 16977 32122 17033 32124
rect 17057 32122 17113 32124
rect 16817 32070 16843 32122
rect 16843 32070 16873 32122
rect 16897 32070 16907 32122
rect 16907 32070 16953 32122
rect 16977 32070 17023 32122
rect 17023 32070 17033 32122
rect 17057 32070 17087 32122
rect 17087 32070 17113 32122
rect 16817 32068 16873 32070
rect 16897 32068 16953 32070
rect 16977 32068 17033 32070
rect 17057 32068 17113 32070
rect 20782 31578 20838 31580
rect 20862 31578 20918 31580
rect 20942 31578 20998 31580
rect 21022 31578 21078 31580
rect 20782 31526 20808 31578
rect 20808 31526 20838 31578
rect 20862 31526 20872 31578
rect 20872 31526 20918 31578
rect 20942 31526 20988 31578
rect 20988 31526 20998 31578
rect 21022 31526 21052 31578
rect 21052 31526 21078 31578
rect 20782 31524 20838 31526
rect 20862 31524 20918 31526
rect 20942 31524 20998 31526
rect 21022 31524 21078 31526
rect 16817 31034 16873 31036
rect 16897 31034 16953 31036
rect 16977 31034 17033 31036
rect 17057 31034 17113 31036
rect 16817 30982 16843 31034
rect 16843 30982 16873 31034
rect 16897 30982 16907 31034
rect 16907 30982 16953 31034
rect 16977 30982 17023 31034
rect 17023 30982 17033 31034
rect 17057 30982 17087 31034
rect 17087 30982 17113 31034
rect 16817 30980 16873 30982
rect 16897 30980 16953 30982
rect 16977 30980 17033 30982
rect 17057 30980 17113 30982
rect 20782 30490 20838 30492
rect 20862 30490 20918 30492
rect 20942 30490 20998 30492
rect 21022 30490 21078 30492
rect 20782 30438 20808 30490
rect 20808 30438 20838 30490
rect 20862 30438 20872 30490
rect 20872 30438 20918 30490
rect 20942 30438 20988 30490
rect 20988 30438 20998 30490
rect 21022 30438 21052 30490
rect 21052 30438 21078 30490
rect 20782 30436 20838 30438
rect 20862 30436 20918 30438
rect 20942 30436 20998 30438
rect 21022 30436 21078 30438
rect 16817 29946 16873 29948
rect 16897 29946 16953 29948
rect 16977 29946 17033 29948
rect 17057 29946 17113 29948
rect 16817 29894 16843 29946
rect 16843 29894 16873 29946
rect 16897 29894 16907 29946
rect 16907 29894 16953 29946
rect 16977 29894 17023 29946
rect 17023 29894 17033 29946
rect 17057 29894 17087 29946
rect 17087 29894 17113 29946
rect 16817 29892 16873 29894
rect 16897 29892 16953 29894
rect 16977 29892 17033 29894
rect 17057 29892 17113 29894
rect 16817 28858 16873 28860
rect 16897 28858 16953 28860
rect 16977 28858 17033 28860
rect 17057 28858 17113 28860
rect 16817 28806 16843 28858
rect 16843 28806 16873 28858
rect 16897 28806 16907 28858
rect 16907 28806 16953 28858
rect 16977 28806 17023 28858
rect 17023 28806 17033 28858
rect 17057 28806 17087 28858
rect 17087 28806 17113 28858
rect 16817 28804 16873 28806
rect 16897 28804 16953 28806
rect 16977 28804 17033 28806
rect 17057 28804 17113 28806
rect 20782 29402 20838 29404
rect 20862 29402 20918 29404
rect 20942 29402 20998 29404
rect 21022 29402 21078 29404
rect 20782 29350 20808 29402
rect 20808 29350 20838 29402
rect 20862 29350 20872 29402
rect 20872 29350 20918 29402
rect 20942 29350 20988 29402
rect 20988 29350 20998 29402
rect 21022 29350 21052 29402
rect 21052 29350 21078 29402
rect 20782 29348 20838 29350
rect 20862 29348 20918 29350
rect 20942 29348 20998 29350
rect 21022 29348 21078 29350
rect 20782 28314 20838 28316
rect 20862 28314 20918 28316
rect 20942 28314 20998 28316
rect 21022 28314 21078 28316
rect 20782 28262 20808 28314
rect 20808 28262 20838 28314
rect 20862 28262 20872 28314
rect 20872 28262 20918 28314
rect 20942 28262 20988 28314
rect 20988 28262 20998 28314
rect 21022 28262 21052 28314
rect 21052 28262 21078 28314
rect 20782 28260 20838 28262
rect 20862 28260 20918 28262
rect 20942 28260 20998 28262
rect 21022 28260 21078 28262
rect 16817 27770 16873 27772
rect 16897 27770 16953 27772
rect 16977 27770 17033 27772
rect 17057 27770 17113 27772
rect 16817 27718 16843 27770
rect 16843 27718 16873 27770
rect 16897 27718 16907 27770
rect 16907 27718 16953 27770
rect 16977 27718 17023 27770
rect 17023 27718 17033 27770
rect 17057 27718 17087 27770
rect 17087 27718 17113 27770
rect 16817 27716 16873 27718
rect 16897 27716 16953 27718
rect 16977 27716 17033 27718
rect 17057 27716 17113 27718
rect 20782 27226 20838 27228
rect 20862 27226 20918 27228
rect 20942 27226 20998 27228
rect 21022 27226 21078 27228
rect 20782 27174 20808 27226
rect 20808 27174 20838 27226
rect 20862 27174 20872 27226
rect 20872 27174 20918 27226
rect 20942 27174 20988 27226
rect 20988 27174 20998 27226
rect 21022 27174 21052 27226
rect 21052 27174 21078 27226
rect 20782 27172 20838 27174
rect 20862 27172 20918 27174
rect 20942 27172 20998 27174
rect 21022 27172 21078 27174
rect 16817 26682 16873 26684
rect 16897 26682 16953 26684
rect 16977 26682 17033 26684
rect 17057 26682 17113 26684
rect 16817 26630 16843 26682
rect 16843 26630 16873 26682
rect 16897 26630 16907 26682
rect 16907 26630 16953 26682
rect 16977 26630 17023 26682
rect 17023 26630 17033 26682
rect 17057 26630 17087 26682
rect 17087 26630 17113 26682
rect 16817 26628 16873 26630
rect 16897 26628 16953 26630
rect 16977 26628 17033 26630
rect 17057 26628 17113 26630
rect 16817 25594 16873 25596
rect 16897 25594 16953 25596
rect 16977 25594 17033 25596
rect 17057 25594 17113 25596
rect 16817 25542 16843 25594
rect 16843 25542 16873 25594
rect 16897 25542 16907 25594
rect 16907 25542 16953 25594
rect 16977 25542 17023 25594
rect 17023 25542 17033 25594
rect 17057 25542 17087 25594
rect 17087 25542 17113 25594
rect 16817 25540 16873 25542
rect 16897 25540 16953 25542
rect 16977 25540 17033 25542
rect 17057 25540 17113 25542
rect 16817 24506 16873 24508
rect 16897 24506 16953 24508
rect 16977 24506 17033 24508
rect 17057 24506 17113 24508
rect 16817 24454 16843 24506
rect 16843 24454 16873 24506
rect 16897 24454 16907 24506
rect 16907 24454 16953 24506
rect 16977 24454 17023 24506
rect 17023 24454 17033 24506
rect 17057 24454 17087 24506
rect 17087 24454 17113 24506
rect 16817 24452 16873 24454
rect 16897 24452 16953 24454
rect 16977 24452 17033 24454
rect 17057 24452 17113 24454
rect 16817 23418 16873 23420
rect 16897 23418 16953 23420
rect 16977 23418 17033 23420
rect 17057 23418 17113 23420
rect 16817 23366 16843 23418
rect 16843 23366 16873 23418
rect 16897 23366 16907 23418
rect 16907 23366 16953 23418
rect 16977 23366 17023 23418
rect 17023 23366 17033 23418
rect 17057 23366 17087 23418
rect 17087 23366 17113 23418
rect 16817 23364 16873 23366
rect 16897 23364 16953 23366
rect 16977 23364 17033 23366
rect 17057 23364 17113 23366
rect 16817 22330 16873 22332
rect 16897 22330 16953 22332
rect 16977 22330 17033 22332
rect 17057 22330 17113 22332
rect 16817 22278 16843 22330
rect 16843 22278 16873 22330
rect 16897 22278 16907 22330
rect 16907 22278 16953 22330
rect 16977 22278 17023 22330
rect 17023 22278 17033 22330
rect 17057 22278 17087 22330
rect 17087 22278 17113 22330
rect 16817 22276 16873 22278
rect 16897 22276 16953 22278
rect 16977 22276 17033 22278
rect 17057 22276 17113 22278
rect 16817 21242 16873 21244
rect 16897 21242 16953 21244
rect 16977 21242 17033 21244
rect 17057 21242 17113 21244
rect 16817 21190 16843 21242
rect 16843 21190 16873 21242
rect 16897 21190 16907 21242
rect 16907 21190 16953 21242
rect 16977 21190 17023 21242
rect 17023 21190 17033 21242
rect 17057 21190 17087 21242
rect 17087 21190 17113 21242
rect 16817 21188 16873 21190
rect 16897 21188 16953 21190
rect 16977 21188 17033 21190
rect 17057 21188 17113 21190
rect 17222 21392 17278 21448
rect 16817 20154 16873 20156
rect 16897 20154 16953 20156
rect 16977 20154 17033 20156
rect 17057 20154 17113 20156
rect 16817 20102 16843 20154
rect 16843 20102 16873 20154
rect 16897 20102 16907 20154
rect 16907 20102 16953 20154
rect 16977 20102 17023 20154
rect 17023 20102 17033 20154
rect 17057 20102 17087 20154
rect 17087 20102 17113 20154
rect 16817 20100 16873 20102
rect 16897 20100 16953 20102
rect 16977 20100 17033 20102
rect 17057 20100 17113 20102
rect 16817 19066 16873 19068
rect 16897 19066 16953 19068
rect 16977 19066 17033 19068
rect 17057 19066 17113 19068
rect 16817 19014 16843 19066
rect 16843 19014 16873 19066
rect 16897 19014 16907 19066
rect 16907 19014 16953 19066
rect 16977 19014 17023 19066
rect 17023 19014 17033 19066
rect 17057 19014 17087 19066
rect 17087 19014 17113 19066
rect 16817 19012 16873 19014
rect 16897 19012 16953 19014
rect 16977 19012 17033 19014
rect 17057 19012 17113 19014
rect 16817 17978 16873 17980
rect 16897 17978 16953 17980
rect 16977 17978 17033 17980
rect 17057 17978 17113 17980
rect 16817 17926 16843 17978
rect 16843 17926 16873 17978
rect 16897 17926 16907 17978
rect 16907 17926 16953 17978
rect 16977 17926 17023 17978
rect 17023 17926 17033 17978
rect 17057 17926 17087 17978
rect 17087 17926 17113 17978
rect 16817 17924 16873 17926
rect 16897 17924 16953 17926
rect 16977 17924 17033 17926
rect 17057 17924 17113 17926
rect 20782 26138 20838 26140
rect 20862 26138 20918 26140
rect 20942 26138 20998 26140
rect 21022 26138 21078 26140
rect 20782 26086 20808 26138
rect 20808 26086 20838 26138
rect 20862 26086 20872 26138
rect 20872 26086 20918 26138
rect 20942 26086 20988 26138
rect 20988 26086 20998 26138
rect 21022 26086 21052 26138
rect 21052 26086 21078 26138
rect 20782 26084 20838 26086
rect 20862 26084 20918 26086
rect 20942 26084 20998 26086
rect 21022 26084 21078 26086
rect 20782 25050 20838 25052
rect 20862 25050 20918 25052
rect 20942 25050 20998 25052
rect 21022 25050 21078 25052
rect 20782 24998 20808 25050
rect 20808 24998 20838 25050
rect 20862 24998 20872 25050
rect 20872 24998 20918 25050
rect 20942 24998 20988 25050
rect 20988 24998 20998 25050
rect 21022 24998 21052 25050
rect 21052 24998 21078 25050
rect 20782 24996 20838 24998
rect 20862 24996 20918 24998
rect 20942 24996 20998 24998
rect 21022 24996 21078 24998
rect 17958 23568 18014 23624
rect 16817 16890 16873 16892
rect 16897 16890 16953 16892
rect 16977 16890 17033 16892
rect 17057 16890 17113 16892
rect 16817 16838 16843 16890
rect 16843 16838 16873 16890
rect 16897 16838 16907 16890
rect 16907 16838 16953 16890
rect 16977 16838 17023 16890
rect 17023 16838 17033 16890
rect 17057 16838 17087 16890
rect 17087 16838 17113 16890
rect 16817 16836 16873 16838
rect 16897 16836 16953 16838
rect 16977 16836 17033 16838
rect 17057 16836 17113 16838
rect 18326 21528 18382 21584
rect 20782 23962 20838 23964
rect 20862 23962 20918 23964
rect 20942 23962 20998 23964
rect 21022 23962 21078 23964
rect 20782 23910 20808 23962
rect 20808 23910 20838 23962
rect 20862 23910 20872 23962
rect 20872 23910 20918 23962
rect 20942 23910 20988 23962
rect 20988 23910 20998 23962
rect 21022 23910 21052 23962
rect 21052 23910 21078 23962
rect 20782 23908 20838 23910
rect 20862 23908 20918 23910
rect 20942 23908 20998 23910
rect 21022 23908 21078 23910
rect 20782 22874 20838 22876
rect 20862 22874 20918 22876
rect 20942 22874 20998 22876
rect 21022 22874 21078 22876
rect 20782 22822 20808 22874
rect 20808 22822 20838 22874
rect 20862 22822 20872 22874
rect 20872 22822 20918 22874
rect 20942 22822 20988 22874
rect 20988 22822 20998 22874
rect 21022 22822 21052 22874
rect 21052 22822 21078 22874
rect 20782 22820 20838 22822
rect 20862 22820 20918 22822
rect 20942 22820 20998 22822
rect 21022 22820 21078 22822
rect 20782 21786 20838 21788
rect 20862 21786 20918 21788
rect 20942 21786 20998 21788
rect 21022 21786 21078 21788
rect 20782 21734 20808 21786
rect 20808 21734 20838 21786
rect 20862 21734 20872 21786
rect 20872 21734 20918 21786
rect 20942 21734 20988 21786
rect 20988 21734 20998 21786
rect 21022 21734 21052 21786
rect 21052 21734 21078 21786
rect 20782 21732 20838 21734
rect 20862 21732 20918 21734
rect 20942 21732 20998 21734
rect 21022 21732 21078 21734
rect 16817 15802 16873 15804
rect 16897 15802 16953 15804
rect 16977 15802 17033 15804
rect 17057 15802 17113 15804
rect 16817 15750 16843 15802
rect 16843 15750 16873 15802
rect 16897 15750 16907 15802
rect 16907 15750 16953 15802
rect 16977 15750 17023 15802
rect 17023 15750 17033 15802
rect 17057 15750 17087 15802
rect 17087 15750 17113 15802
rect 16817 15748 16873 15750
rect 16897 15748 16953 15750
rect 16977 15748 17033 15750
rect 17057 15748 17113 15750
rect 15290 8880 15346 8936
rect 16817 14714 16873 14716
rect 16897 14714 16953 14716
rect 16977 14714 17033 14716
rect 17057 14714 17113 14716
rect 16817 14662 16843 14714
rect 16843 14662 16873 14714
rect 16897 14662 16907 14714
rect 16907 14662 16953 14714
rect 16977 14662 17023 14714
rect 17023 14662 17033 14714
rect 17057 14662 17087 14714
rect 17087 14662 17113 14714
rect 16817 14660 16873 14662
rect 16897 14660 16953 14662
rect 16977 14660 17033 14662
rect 17057 14660 17113 14662
rect 16817 13626 16873 13628
rect 16897 13626 16953 13628
rect 16977 13626 17033 13628
rect 17057 13626 17113 13628
rect 16817 13574 16843 13626
rect 16843 13574 16873 13626
rect 16897 13574 16907 13626
rect 16907 13574 16953 13626
rect 16977 13574 17023 13626
rect 17023 13574 17033 13626
rect 17057 13574 17087 13626
rect 17087 13574 17113 13626
rect 16817 13572 16873 13574
rect 16897 13572 16953 13574
rect 16977 13572 17033 13574
rect 17057 13572 17113 13574
rect 16817 12538 16873 12540
rect 16897 12538 16953 12540
rect 16977 12538 17033 12540
rect 17057 12538 17113 12540
rect 16817 12486 16843 12538
rect 16843 12486 16873 12538
rect 16897 12486 16907 12538
rect 16907 12486 16953 12538
rect 16977 12486 17023 12538
rect 17023 12486 17033 12538
rect 17057 12486 17087 12538
rect 17087 12486 17113 12538
rect 16817 12484 16873 12486
rect 16897 12484 16953 12486
rect 16977 12484 17033 12486
rect 17057 12484 17113 12486
rect 16817 11450 16873 11452
rect 16897 11450 16953 11452
rect 16977 11450 17033 11452
rect 17057 11450 17113 11452
rect 16817 11398 16843 11450
rect 16843 11398 16873 11450
rect 16897 11398 16907 11450
rect 16907 11398 16953 11450
rect 16977 11398 17023 11450
rect 17023 11398 17033 11450
rect 17057 11398 17087 11450
rect 17087 11398 17113 11450
rect 16817 11396 16873 11398
rect 16897 11396 16953 11398
rect 16977 11396 17033 11398
rect 17057 11396 17113 11398
rect 16817 10362 16873 10364
rect 16897 10362 16953 10364
rect 16977 10362 17033 10364
rect 17057 10362 17113 10364
rect 16817 10310 16843 10362
rect 16843 10310 16873 10362
rect 16897 10310 16907 10362
rect 16907 10310 16953 10362
rect 16977 10310 17023 10362
rect 17023 10310 17033 10362
rect 17057 10310 17087 10362
rect 17087 10310 17113 10362
rect 16817 10308 16873 10310
rect 16897 10308 16953 10310
rect 16977 10308 17033 10310
rect 17057 10308 17113 10310
rect 20782 20698 20838 20700
rect 20862 20698 20918 20700
rect 20942 20698 20998 20700
rect 21022 20698 21078 20700
rect 20782 20646 20808 20698
rect 20808 20646 20838 20698
rect 20862 20646 20872 20698
rect 20872 20646 20918 20698
rect 20942 20646 20988 20698
rect 20988 20646 20998 20698
rect 21022 20646 21052 20698
rect 21052 20646 21078 20698
rect 20782 20644 20838 20646
rect 20862 20644 20918 20646
rect 20942 20644 20998 20646
rect 21022 20644 21078 20646
rect 20782 19610 20838 19612
rect 20862 19610 20918 19612
rect 20942 19610 20998 19612
rect 21022 19610 21078 19612
rect 20782 19558 20808 19610
rect 20808 19558 20838 19610
rect 20862 19558 20872 19610
rect 20872 19558 20918 19610
rect 20942 19558 20988 19610
rect 20988 19558 20998 19610
rect 21022 19558 21052 19610
rect 21052 19558 21078 19610
rect 20782 19556 20838 19558
rect 20862 19556 20918 19558
rect 20942 19556 20998 19558
rect 21022 19556 21078 19558
rect 20782 18522 20838 18524
rect 20862 18522 20918 18524
rect 20942 18522 20998 18524
rect 21022 18522 21078 18524
rect 20782 18470 20808 18522
rect 20808 18470 20838 18522
rect 20862 18470 20872 18522
rect 20872 18470 20918 18522
rect 20942 18470 20988 18522
rect 20988 18470 20998 18522
rect 21022 18470 21052 18522
rect 21052 18470 21078 18522
rect 20782 18468 20838 18470
rect 20862 18468 20918 18470
rect 20942 18468 20998 18470
rect 21022 18468 21078 18470
rect 20782 17434 20838 17436
rect 20862 17434 20918 17436
rect 20942 17434 20998 17436
rect 21022 17434 21078 17436
rect 20782 17382 20808 17434
rect 20808 17382 20838 17434
rect 20862 17382 20872 17434
rect 20872 17382 20918 17434
rect 20942 17382 20988 17434
rect 20988 17382 20998 17434
rect 21022 17382 21052 17434
rect 21052 17382 21078 17434
rect 20782 17380 20838 17382
rect 20862 17380 20918 17382
rect 20942 17380 20998 17382
rect 21022 17380 21078 17382
rect 20782 16346 20838 16348
rect 20862 16346 20918 16348
rect 20942 16346 20998 16348
rect 21022 16346 21078 16348
rect 20782 16294 20808 16346
rect 20808 16294 20838 16346
rect 20862 16294 20872 16346
rect 20872 16294 20918 16346
rect 20942 16294 20988 16346
rect 20988 16294 20998 16346
rect 21022 16294 21052 16346
rect 21052 16294 21078 16346
rect 20782 16292 20838 16294
rect 20862 16292 20918 16294
rect 20942 16292 20998 16294
rect 21022 16292 21078 16294
rect 20782 15258 20838 15260
rect 20862 15258 20918 15260
rect 20942 15258 20998 15260
rect 21022 15258 21078 15260
rect 20782 15206 20808 15258
rect 20808 15206 20838 15258
rect 20862 15206 20872 15258
rect 20872 15206 20918 15258
rect 20942 15206 20988 15258
rect 20988 15206 20998 15258
rect 21022 15206 21052 15258
rect 21052 15206 21078 15258
rect 20782 15204 20838 15206
rect 20862 15204 20918 15206
rect 20942 15204 20998 15206
rect 21022 15204 21078 15206
rect 20782 14170 20838 14172
rect 20862 14170 20918 14172
rect 20942 14170 20998 14172
rect 21022 14170 21078 14172
rect 20782 14118 20808 14170
rect 20808 14118 20838 14170
rect 20862 14118 20872 14170
rect 20872 14118 20918 14170
rect 20942 14118 20988 14170
rect 20988 14118 20998 14170
rect 21022 14118 21052 14170
rect 21052 14118 21078 14170
rect 20782 14116 20838 14118
rect 20862 14116 20918 14118
rect 20942 14116 20998 14118
rect 21022 14116 21078 14118
rect 16486 9288 16542 9344
rect 16817 9274 16873 9276
rect 16897 9274 16953 9276
rect 16977 9274 17033 9276
rect 17057 9274 17113 9276
rect 16817 9222 16843 9274
rect 16843 9222 16873 9274
rect 16897 9222 16907 9274
rect 16907 9222 16953 9274
rect 16977 9222 17023 9274
rect 17023 9222 17033 9274
rect 17057 9222 17087 9274
rect 17087 9222 17113 9274
rect 16817 9220 16873 9222
rect 16897 9220 16953 9222
rect 16977 9220 17033 9222
rect 17057 9220 17113 9222
rect 16817 8186 16873 8188
rect 16897 8186 16953 8188
rect 16977 8186 17033 8188
rect 17057 8186 17113 8188
rect 16817 8134 16843 8186
rect 16843 8134 16873 8186
rect 16897 8134 16907 8186
rect 16907 8134 16953 8186
rect 16977 8134 17023 8186
rect 17023 8134 17033 8186
rect 17057 8134 17087 8186
rect 17087 8134 17113 8186
rect 16817 8132 16873 8134
rect 16897 8132 16953 8134
rect 16977 8132 17033 8134
rect 17057 8132 17113 8134
rect 17498 9016 17554 9072
rect 18234 9444 18290 9480
rect 18234 9424 18236 9444
rect 18236 9424 18288 9444
rect 18288 9424 18290 9444
rect 20782 13082 20838 13084
rect 20862 13082 20918 13084
rect 20942 13082 20998 13084
rect 21022 13082 21078 13084
rect 20782 13030 20808 13082
rect 20808 13030 20838 13082
rect 20862 13030 20872 13082
rect 20872 13030 20918 13082
rect 20942 13030 20988 13082
rect 20988 13030 20998 13082
rect 21022 13030 21052 13082
rect 21052 13030 21078 13082
rect 20782 13028 20838 13030
rect 20862 13028 20918 13030
rect 20942 13028 20998 13030
rect 21022 13028 21078 13030
rect 20782 11994 20838 11996
rect 20862 11994 20918 11996
rect 20942 11994 20998 11996
rect 21022 11994 21078 11996
rect 20782 11942 20808 11994
rect 20808 11942 20838 11994
rect 20862 11942 20872 11994
rect 20872 11942 20918 11994
rect 20942 11942 20988 11994
rect 20988 11942 20998 11994
rect 21022 11942 21052 11994
rect 21052 11942 21078 11994
rect 20782 11940 20838 11942
rect 20862 11940 20918 11942
rect 20942 11940 20998 11942
rect 21022 11940 21078 11942
rect 20782 10906 20838 10908
rect 20862 10906 20918 10908
rect 20942 10906 20998 10908
rect 21022 10906 21078 10908
rect 20782 10854 20808 10906
rect 20808 10854 20838 10906
rect 20862 10854 20872 10906
rect 20872 10854 20918 10906
rect 20942 10854 20988 10906
rect 20988 10854 20998 10906
rect 21022 10854 21052 10906
rect 21052 10854 21078 10906
rect 20782 10852 20838 10854
rect 20862 10852 20918 10854
rect 20942 10852 20998 10854
rect 21022 10852 21078 10854
rect 19154 10648 19210 10704
rect 16817 7098 16873 7100
rect 16897 7098 16953 7100
rect 16977 7098 17033 7100
rect 17057 7098 17113 7100
rect 16817 7046 16843 7098
rect 16843 7046 16873 7098
rect 16897 7046 16907 7098
rect 16907 7046 16953 7098
rect 16977 7046 17023 7098
rect 17023 7046 17033 7098
rect 17057 7046 17087 7098
rect 17087 7046 17113 7098
rect 16817 7044 16873 7046
rect 16897 7044 16953 7046
rect 16977 7044 17033 7046
rect 17057 7044 17113 7046
rect 20902 9968 20958 10024
rect 20782 9818 20838 9820
rect 20862 9818 20918 9820
rect 20942 9818 20998 9820
rect 21022 9818 21078 9820
rect 20782 9766 20808 9818
rect 20808 9766 20838 9818
rect 20862 9766 20872 9818
rect 20872 9766 20918 9818
rect 20942 9766 20988 9818
rect 20988 9766 20998 9818
rect 21022 9766 21052 9818
rect 21052 9766 21078 9818
rect 20782 9764 20838 9766
rect 20862 9764 20918 9766
rect 20942 9764 20998 9766
rect 21022 9764 21078 9766
rect 20782 8730 20838 8732
rect 20862 8730 20918 8732
rect 20942 8730 20998 8732
rect 21022 8730 21078 8732
rect 20782 8678 20808 8730
rect 20808 8678 20838 8730
rect 20862 8678 20872 8730
rect 20872 8678 20918 8730
rect 20942 8678 20988 8730
rect 20988 8678 20998 8730
rect 21022 8678 21052 8730
rect 21052 8678 21078 8730
rect 20782 8676 20838 8678
rect 20862 8676 20918 8678
rect 20942 8676 20998 8678
rect 21022 8676 21078 8678
rect 20782 7642 20838 7644
rect 20862 7642 20918 7644
rect 20942 7642 20998 7644
rect 21022 7642 21078 7644
rect 20782 7590 20808 7642
rect 20808 7590 20838 7642
rect 20862 7590 20872 7642
rect 20872 7590 20918 7642
rect 20942 7590 20988 7642
rect 20988 7590 20998 7642
rect 21022 7590 21052 7642
rect 21052 7590 21078 7642
rect 20782 7588 20838 7590
rect 20862 7588 20918 7590
rect 20942 7588 20998 7590
rect 21022 7588 21078 7590
rect 20782 6554 20838 6556
rect 20862 6554 20918 6556
rect 20942 6554 20998 6556
rect 21022 6554 21078 6556
rect 20782 6502 20808 6554
rect 20808 6502 20838 6554
rect 20862 6502 20872 6554
rect 20872 6502 20918 6554
rect 20942 6502 20988 6554
rect 20988 6502 20998 6554
rect 21022 6502 21052 6554
rect 21052 6502 21078 6554
rect 20782 6500 20838 6502
rect 20862 6500 20918 6502
rect 20942 6500 20998 6502
rect 21022 6500 21078 6502
rect 16817 6010 16873 6012
rect 16897 6010 16953 6012
rect 16977 6010 17033 6012
rect 17057 6010 17113 6012
rect 16817 5958 16843 6010
rect 16843 5958 16873 6010
rect 16897 5958 16907 6010
rect 16907 5958 16953 6010
rect 16977 5958 17023 6010
rect 17023 5958 17033 6010
rect 17057 5958 17087 6010
rect 17087 5958 17113 6010
rect 16817 5956 16873 5958
rect 16897 5956 16953 5958
rect 16977 5956 17033 5958
rect 17057 5956 17113 5958
rect 20782 5466 20838 5468
rect 20862 5466 20918 5468
rect 20942 5466 20998 5468
rect 21022 5466 21078 5468
rect 20782 5414 20808 5466
rect 20808 5414 20838 5466
rect 20862 5414 20872 5466
rect 20872 5414 20918 5466
rect 20942 5414 20988 5466
rect 20988 5414 20998 5466
rect 21022 5414 21052 5466
rect 21052 5414 21078 5466
rect 20782 5412 20838 5414
rect 20862 5412 20918 5414
rect 20942 5412 20998 5414
rect 21022 5412 21078 5414
rect 16817 4922 16873 4924
rect 16897 4922 16953 4924
rect 16977 4922 17033 4924
rect 17057 4922 17113 4924
rect 16817 4870 16843 4922
rect 16843 4870 16873 4922
rect 16897 4870 16907 4922
rect 16907 4870 16953 4922
rect 16977 4870 17023 4922
rect 17023 4870 17033 4922
rect 17057 4870 17087 4922
rect 17087 4870 17113 4922
rect 16817 4868 16873 4870
rect 16897 4868 16953 4870
rect 16977 4868 17033 4870
rect 17057 4868 17113 4870
rect 20782 4378 20838 4380
rect 20862 4378 20918 4380
rect 20942 4378 20998 4380
rect 21022 4378 21078 4380
rect 20782 4326 20808 4378
rect 20808 4326 20838 4378
rect 20862 4326 20872 4378
rect 20872 4326 20918 4378
rect 20942 4326 20988 4378
rect 20988 4326 20998 4378
rect 21022 4326 21052 4378
rect 21052 4326 21078 4378
rect 20782 4324 20838 4326
rect 20862 4324 20918 4326
rect 20942 4324 20998 4326
rect 21022 4324 21078 4326
rect 16817 3834 16873 3836
rect 16897 3834 16953 3836
rect 16977 3834 17033 3836
rect 17057 3834 17113 3836
rect 16817 3782 16843 3834
rect 16843 3782 16873 3834
rect 16897 3782 16907 3834
rect 16907 3782 16953 3834
rect 16977 3782 17023 3834
rect 17023 3782 17033 3834
rect 17057 3782 17087 3834
rect 17087 3782 17113 3834
rect 16817 3780 16873 3782
rect 16897 3780 16953 3782
rect 16977 3780 17033 3782
rect 17057 3780 17113 3782
rect 16817 2746 16873 2748
rect 16897 2746 16953 2748
rect 16977 2746 17033 2748
rect 17057 2746 17113 2748
rect 16817 2694 16843 2746
rect 16843 2694 16873 2746
rect 16897 2694 16907 2746
rect 16907 2694 16953 2746
rect 16977 2694 17023 2746
rect 17023 2694 17033 2746
rect 17057 2694 17087 2746
rect 17087 2694 17113 2746
rect 16817 2692 16873 2694
rect 16897 2692 16953 2694
rect 16977 2692 17033 2694
rect 17057 2692 17113 2694
rect 20782 3290 20838 3292
rect 20862 3290 20918 3292
rect 20942 3290 20998 3292
rect 21022 3290 21078 3292
rect 20782 3238 20808 3290
rect 20808 3238 20838 3290
rect 20862 3238 20872 3290
rect 20872 3238 20918 3290
rect 20942 3238 20988 3290
rect 20988 3238 20998 3290
rect 21022 3238 21052 3290
rect 21052 3238 21078 3290
rect 20782 3236 20838 3238
rect 20862 3236 20918 3238
rect 20942 3236 20998 3238
rect 21022 3236 21078 3238
rect 20782 2202 20838 2204
rect 20862 2202 20918 2204
rect 20942 2202 20998 2204
rect 21022 2202 21078 2204
rect 20782 2150 20808 2202
rect 20808 2150 20838 2202
rect 20862 2150 20872 2202
rect 20872 2150 20918 2202
rect 20942 2150 20988 2202
rect 20988 2150 20998 2202
rect 21022 2150 21052 2202
rect 21052 2150 21078 2202
rect 20782 2148 20838 2150
rect 20862 2148 20918 2150
rect 20942 2148 20998 2150
rect 21022 2148 21078 2150
<< metal3 >>
rect 8874 47360 9194 47361
rect 0 47290 800 47320
rect 8874 47296 8882 47360
rect 8946 47296 8962 47360
rect 9026 47296 9042 47360
rect 9106 47296 9122 47360
rect 9186 47296 9194 47360
rect 8874 47295 9194 47296
rect 16805 47360 17125 47361
rect 16805 47296 16813 47360
rect 16877 47296 16893 47360
rect 16957 47296 16973 47360
rect 17037 47296 17053 47360
rect 17117 47296 17125 47360
rect 16805 47295 17125 47296
rect 3049 47290 3115 47293
rect 0 47288 3115 47290
rect 0 47232 3054 47288
rect 3110 47232 3115 47288
rect 0 47230 3115 47232
rect 0 47200 800 47230
rect 3049 47227 3115 47230
rect 4909 46816 5229 46817
rect 4909 46752 4917 46816
rect 4981 46752 4997 46816
rect 5061 46752 5077 46816
rect 5141 46752 5157 46816
rect 5221 46752 5229 46816
rect 4909 46751 5229 46752
rect 12840 46816 13160 46817
rect 12840 46752 12848 46816
rect 12912 46752 12928 46816
rect 12992 46752 13008 46816
rect 13072 46752 13088 46816
rect 13152 46752 13160 46816
rect 12840 46751 13160 46752
rect 20770 46816 21090 46817
rect 20770 46752 20778 46816
rect 20842 46752 20858 46816
rect 20922 46752 20938 46816
rect 21002 46752 21018 46816
rect 21082 46752 21090 46816
rect 20770 46751 21090 46752
rect 8874 46272 9194 46273
rect 8874 46208 8882 46272
rect 8946 46208 8962 46272
rect 9026 46208 9042 46272
rect 9106 46208 9122 46272
rect 9186 46208 9194 46272
rect 8874 46207 9194 46208
rect 16805 46272 17125 46273
rect 16805 46208 16813 46272
rect 16877 46208 16893 46272
rect 16957 46208 16973 46272
rect 17037 46208 17053 46272
rect 17117 46208 17125 46272
rect 16805 46207 17125 46208
rect 4909 45728 5229 45729
rect 4909 45664 4917 45728
rect 4981 45664 4997 45728
rect 5061 45664 5077 45728
rect 5141 45664 5157 45728
rect 5221 45664 5229 45728
rect 4909 45663 5229 45664
rect 12840 45728 13160 45729
rect 12840 45664 12848 45728
rect 12912 45664 12928 45728
rect 12992 45664 13008 45728
rect 13072 45664 13088 45728
rect 13152 45664 13160 45728
rect 12840 45663 13160 45664
rect 20770 45728 21090 45729
rect 20770 45664 20778 45728
rect 20842 45664 20858 45728
rect 20922 45664 20938 45728
rect 21002 45664 21018 45728
rect 21082 45664 21090 45728
rect 20770 45663 21090 45664
rect 8874 45184 9194 45185
rect 8874 45120 8882 45184
rect 8946 45120 8962 45184
rect 9026 45120 9042 45184
rect 9106 45120 9122 45184
rect 9186 45120 9194 45184
rect 8874 45119 9194 45120
rect 16805 45184 17125 45185
rect 16805 45120 16813 45184
rect 16877 45120 16893 45184
rect 16957 45120 16973 45184
rect 17037 45120 17053 45184
rect 17117 45120 17125 45184
rect 16805 45119 17125 45120
rect 4909 44640 5229 44641
rect 4909 44576 4917 44640
rect 4981 44576 4997 44640
rect 5061 44576 5077 44640
rect 5141 44576 5157 44640
rect 5221 44576 5229 44640
rect 4909 44575 5229 44576
rect 12840 44640 13160 44641
rect 12840 44576 12848 44640
rect 12912 44576 12928 44640
rect 12992 44576 13008 44640
rect 13072 44576 13088 44640
rect 13152 44576 13160 44640
rect 12840 44575 13160 44576
rect 20770 44640 21090 44641
rect 20770 44576 20778 44640
rect 20842 44576 20858 44640
rect 20922 44576 20938 44640
rect 21002 44576 21018 44640
rect 21082 44576 21090 44640
rect 20770 44575 21090 44576
rect 8874 44096 9194 44097
rect 8874 44032 8882 44096
rect 8946 44032 8962 44096
rect 9026 44032 9042 44096
rect 9106 44032 9122 44096
rect 9186 44032 9194 44096
rect 8874 44031 9194 44032
rect 16805 44096 17125 44097
rect 16805 44032 16813 44096
rect 16877 44032 16893 44096
rect 16957 44032 16973 44096
rect 17037 44032 17053 44096
rect 17117 44032 17125 44096
rect 16805 44031 17125 44032
rect 4909 43552 5229 43553
rect 4909 43488 4917 43552
rect 4981 43488 4997 43552
rect 5061 43488 5077 43552
rect 5141 43488 5157 43552
rect 5221 43488 5229 43552
rect 4909 43487 5229 43488
rect 12840 43552 13160 43553
rect 12840 43488 12848 43552
rect 12912 43488 12928 43552
rect 12992 43488 13008 43552
rect 13072 43488 13088 43552
rect 13152 43488 13160 43552
rect 12840 43487 13160 43488
rect 20770 43552 21090 43553
rect 20770 43488 20778 43552
rect 20842 43488 20858 43552
rect 20922 43488 20938 43552
rect 21002 43488 21018 43552
rect 21082 43488 21090 43552
rect 20770 43487 21090 43488
rect 8874 43008 9194 43009
rect 8874 42944 8882 43008
rect 8946 42944 8962 43008
rect 9026 42944 9042 43008
rect 9106 42944 9122 43008
rect 9186 42944 9194 43008
rect 8874 42943 9194 42944
rect 16805 43008 17125 43009
rect 16805 42944 16813 43008
rect 16877 42944 16893 43008
rect 16957 42944 16973 43008
rect 17037 42944 17053 43008
rect 17117 42944 17125 43008
rect 16805 42943 17125 42944
rect 4909 42464 5229 42465
rect 4909 42400 4917 42464
rect 4981 42400 4997 42464
rect 5061 42400 5077 42464
rect 5141 42400 5157 42464
rect 5221 42400 5229 42464
rect 4909 42399 5229 42400
rect 12840 42464 13160 42465
rect 12840 42400 12848 42464
rect 12912 42400 12928 42464
rect 12992 42400 13008 42464
rect 13072 42400 13088 42464
rect 13152 42400 13160 42464
rect 12840 42399 13160 42400
rect 20770 42464 21090 42465
rect 20770 42400 20778 42464
rect 20842 42400 20858 42464
rect 20922 42400 20938 42464
rect 21002 42400 21018 42464
rect 21082 42400 21090 42464
rect 20770 42399 21090 42400
rect 8874 41920 9194 41921
rect 8874 41856 8882 41920
rect 8946 41856 8962 41920
rect 9026 41856 9042 41920
rect 9106 41856 9122 41920
rect 9186 41856 9194 41920
rect 8874 41855 9194 41856
rect 16805 41920 17125 41921
rect 16805 41856 16813 41920
rect 16877 41856 16893 41920
rect 16957 41856 16973 41920
rect 17037 41856 17053 41920
rect 17117 41856 17125 41920
rect 16805 41855 17125 41856
rect 0 41714 800 41744
rect 3325 41714 3391 41717
rect 0 41712 3391 41714
rect 0 41656 3330 41712
rect 3386 41656 3391 41712
rect 0 41654 3391 41656
rect 0 41624 800 41654
rect 3325 41651 3391 41654
rect 4909 41376 5229 41377
rect 4909 41312 4917 41376
rect 4981 41312 4997 41376
rect 5061 41312 5077 41376
rect 5141 41312 5157 41376
rect 5221 41312 5229 41376
rect 4909 41311 5229 41312
rect 12840 41376 13160 41377
rect 12840 41312 12848 41376
rect 12912 41312 12928 41376
rect 12992 41312 13008 41376
rect 13072 41312 13088 41376
rect 13152 41312 13160 41376
rect 12840 41311 13160 41312
rect 20770 41376 21090 41377
rect 20770 41312 20778 41376
rect 20842 41312 20858 41376
rect 20922 41312 20938 41376
rect 21002 41312 21018 41376
rect 21082 41312 21090 41376
rect 20770 41311 21090 41312
rect 8874 40832 9194 40833
rect 8874 40768 8882 40832
rect 8946 40768 8962 40832
rect 9026 40768 9042 40832
rect 9106 40768 9122 40832
rect 9186 40768 9194 40832
rect 8874 40767 9194 40768
rect 16805 40832 17125 40833
rect 16805 40768 16813 40832
rect 16877 40768 16893 40832
rect 16957 40768 16973 40832
rect 17037 40768 17053 40832
rect 17117 40768 17125 40832
rect 16805 40767 17125 40768
rect 4909 40288 5229 40289
rect 4909 40224 4917 40288
rect 4981 40224 4997 40288
rect 5061 40224 5077 40288
rect 5141 40224 5157 40288
rect 5221 40224 5229 40288
rect 4909 40223 5229 40224
rect 12840 40288 13160 40289
rect 12840 40224 12848 40288
rect 12912 40224 12928 40288
rect 12992 40224 13008 40288
rect 13072 40224 13088 40288
rect 13152 40224 13160 40288
rect 12840 40223 13160 40224
rect 20770 40288 21090 40289
rect 20770 40224 20778 40288
rect 20842 40224 20858 40288
rect 20922 40224 20938 40288
rect 21002 40224 21018 40288
rect 21082 40224 21090 40288
rect 20770 40223 21090 40224
rect 8874 39744 9194 39745
rect 8874 39680 8882 39744
rect 8946 39680 8962 39744
rect 9026 39680 9042 39744
rect 9106 39680 9122 39744
rect 9186 39680 9194 39744
rect 8874 39679 9194 39680
rect 16805 39744 17125 39745
rect 16805 39680 16813 39744
rect 16877 39680 16893 39744
rect 16957 39680 16973 39744
rect 17037 39680 17053 39744
rect 17117 39680 17125 39744
rect 16805 39679 17125 39680
rect 4909 39200 5229 39201
rect 4909 39136 4917 39200
rect 4981 39136 4997 39200
rect 5061 39136 5077 39200
rect 5141 39136 5157 39200
rect 5221 39136 5229 39200
rect 4909 39135 5229 39136
rect 12840 39200 13160 39201
rect 12840 39136 12848 39200
rect 12912 39136 12928 39200
rect 12992 39136 13008 39200
rect 13072 39136 13088 39200
rect 13152 39136 13160 39200
rect 12840 39135 13160 39136
rect 20770 39200 21090 39201
rect 20770 39136 20778 39200
rect 20842 39136 20858 39200
rect 20922 39136 20938 39200
rect 21002 39136 21018 39200
rect 21082 39136 21090 39200
rect 20770 39135 21090 39136
rect 2405 38994 2471 38997
rect 2957 38994 3023 38997
rect 7925 38994 7991 38997
rect 9581 38994 9647 38997
rect 2405 38992 9647 38994
rect 2405 38936 2410 38992
rect 2466 38936 2962 38992
rect 3018 38936 7930 38992
rect 7986 38936 9586 38992
rect 9642 38936 9647 38992
rect 2405 38934 9647 38936
rect 2405 38931 2471 38934
rect 2957 38931 3023 38934
rect 7925 38931 7991 38934
rect 9581 38931 9647 38934
rect 12065 38994 12131 38997
rect 16665 38994 16731 38997
rect 12065 38992 16731 38994
rect 12065 38936 12070 38992
rect 12126 38936 16670 38992
rect 16726 38936 16731 38992
rect 12065 38934 16731 38936
rect 12065 38931 12131 38934
rect 16665 38931 16731 38934
rect 11329 38858 11395 38861
rect 14089 38858 14155 38861
rect 11329 38856 14155 38858
rect 11329 38800 11334 38856
rect 11390 38800 14094 38856
rect 14150 38800 14155 38856
rect 11329 38798 14155 38800
rect 11329 38795 11395 38798
rect 14089 38795 14155 38798
rect 8874 38656 9194 38657
rect 8874 38592 8882 38656
rect 8946 38592 8962 38656
rect 9026 38592 9042 38656
rect 9106 38592 9122 38656
rect 9186 38592 9194 38656
rect 8874 38591 9194 38592
rect 16805 38656 17125 38657
rect 16805 38592 16813 38656
rect 16877 38592 16893 38656
rect 16957 38592 16973 38656
rect 17037 38592 17053 38656
rect 17117 38592 17125 38656
rect 16805 38591 17125 38592
rect 4909 38112 5229 38113
rect 4909 38048 4917 38112
rect 4981 38048 4997 38112
rect 5061 38048 5077 38112
rect 5141 38048 5157 38112
rect 5221 38048 5229 38112
rect 4909 38047 5229 38048
rect 12840 38112 13160 38113
rect 12840 38048 12848 38112
rect 12912 38048 12928 38112
rect 12992 38048 13008 38112
rect 13072 38048 13088 38112
rect 13152 38048 13160 38112
rect 12840 38047 13160 38048
rect 20770 38112 21090 38113
rect 20770 38048 20778 38112
rect 20842 38048 20858 38112
rect 20922 38048 20938 38112
rect 21002 38048 21018 38112
rect 21082 38048 21090 38112
rect 20770 38047 21090 38048
rect 8874 37568 9194 37569
rect 8874 37504 8882 37568
rect 8946 37504 8962 37568
rect 9026 37504 9042 37568
rect 9106 37504 9122 37568
rect 9186 37504 9194 37568
rect 8874 37503 9194 37504
rect 16805 37568 17125 37569
rect 16805 37504 16813 37568
rect 16877 37504 16893 37568
rect 16957 37504 16973 37568
rect 17037 37504 17053 37568
rect 17117 37504 17125 37568
rect 16805 37503 17125 37504
rect 4909 37024 5229 37025
rect 4909 36960 4917 37024
rect 4981 36960 4997 37024
rect 5061 36960 5077 37024
rect 5141 36960 5157 37024
rect 5221 36960 5229 37024
rect 4909 36959 5229 36960
rect 12840 37024 13160 37025
rect 12840 36960 12848 37024
rect 12912 36960 12928 37024
rect 12992 36960 13008 37024
rect 13072 36960 13088 37024
rect 13152 36960 13160 37024
rect 12840 36959 13160 36960
rect 20770 37024 21090 37025
rect 20770 36960 20778 37024
rect 20842 36960 20858 37024
rect 20922 36960 20938 37024
rect 21002 36960 21018 37024
rect 21082 36960 21090 37024
rect 20770 36959 21090 36960
rect 8874 36480 9194 36481
rect 8874 36416 8882 36480
rect 8946 36416 8962 36480
rect 9026 36416 9042 36480
rect 9106 36416 9122 36480
rect 9186 36416 9194 36480
rect 8874 36415 9194 36416
rect 16805 36480 17125 36481
rect 16805 36416 16813 36480
rect 16877 36416 16893 36480
rect 16957 36416 16973 36480
rect 17037 36416 17053 36480
rect 17117 36416 17125 36480
rect 16805 36415 17125 36416
rect 0 36138 800 36168
rect 3325 36138 3391 36141
rect 0 36136 3391 36138
rect 0 36080 3330 36136
rect 3386 36080 3391 36136
rect 0 36078 3391 36080
rect 0 36048 800 36078
rect 3325 36075 3391 36078
rect 4909 35936 5229 35937
rect 4909 35872 4917 35936
rect 4981 35872 4997 35936
rect 5061 35872 5077 35936
rect 5141 35872 5157 35936
rect 5221 35872 5229 35936
rect 4909 35871 5229 35872
rect 12840 35936 13160 35937
rect 12840 35872 12848 35936
rect 12912 35872 12928 35936
rect 12992 35872 13008 35936
rect 13072 35872 13088 35936
rect 13152 35872 13160 35936
rect 12840 35871 13160 35872
rect 20770 35936 21090 35937
rect 20770 35872 20778 35936
rect 20842 35872 20858 35936
rect 20922 35872 20938 35936
rect 21002 35872 21018 35936
rect 21082 35872 21090 35936
rect 20770 35871 21090 35872
rect 8874 35392 9194 35393
rect 8874 35328 8882 35392
rect 8946 35328 8962 35392
rect 9026 35328 9042 35392
rect 9106 35328 9122 35392
rect 9186 35328 9194 35392
rect 8874 35327 9194 35328
rect 16805 35392 17125 35393
rect 16805 35328 16813 35392
rect 16877 35328 16893 35392
rect 16957 35328 16973 35392
rect 17037 35328 17053 35392
rect 17117 35328 17125 35392
rect 16805 35327 17125 35328
rect 4909 34848 5229 34849
rect 4909 34784 4917 34848
rect 4981 34784 4997 34848
rect 5061 34784 5077 34848
rect 5141 34784 5157 34848
rect 5221 34784 5229 34848
rect 4909 34783 5229 34784
rect 12840 34848 13160 34849
rect 12840 34784 12848 34848
rect 12912 34784 12928 34848
rect 12992 34784 13008 34848
rect 13072 34784 13088 34848
rect 13152 34784 13160 34848
rect 12840 34783 13160 34784
rect 20770 34848 21090 34849
rect 20770 34784 20778 34848
rect 20842 34784 20858 34848
rect 20922 34784 20938 34848
rect 21002 34784 21018 34848
rect 21082 34784 21090 34848
rect 20770 34783 21090 34784
rect 8874 34304 9194 34305
rect 8874 34240 8882 34304
rect 8946 34240 8962 34304
rect 9026 34240 9042 34304
rect 9106 34240 9122 34304
rect 9186 34240 9194 34304
rect 8874 34239 9194 34240
rect 16805 34304 17125 34305
rect 16805 34240 16813 34304
rect 16877 34240 16893 34304
rect 16957 34240 16973 34304
rect 17037 34240 17053 34304
rect 17117 34240 17125 34304
rect 16805 34239 17125 34240
rect 5349 34236 5415 34237
rect 5349 34232 5396 34236
rect 5460 34234 5466 34236
rect 5349 34176 5354 34232
rect 5349 34172 5396 34176
rect 5460 34174 5506 34234
rect 5460 34172 5466 34174
rect 5349 34171 5415 34172
rect 4909 33760 5229 33761
rect 4909 33696 4917 33760
rect 4981 33696 4997 33760
rect 5061 33696 5077 33760
rect 5141 33696 5157 33760
rect 5221 33696 5229 33760
rect 4909 33695 5229 33696
rect 12840 33760 13160 33761
rect 12840 33696 12848 33760
rect 12912 33696 12928 33760
rect 12992 33696 13008 33760
rect 13072 33696 13088 33760
rect 13152 33696 13160 33760
rect 12840 33695 13160 33696
rect 20770 33760 21090 33761
rect 20770 33696 20778 33760
rect 20842 33696 20858 33760
rect 20922 33696 20938 33760
rect 21002 33696 21018 33760
rect 21082 33696 21090 33760
rect 20770 33695 21090 33696
rect 8874 33216 9194 33217
rect 8874 33152 8882 33216
rect 8946 33152 8962 33216
rect 9026 33152 9042 33216
rect 9106 33152 9122 33216
rect 9186 33152 9194 33216
rect 8874 33151 9194 33152
rect 16805 33216 17125 33217
rect 16805 33152 16813 33216
rect 16877 33152 16893 33216
rect 16957 33152 16973 33216
rect 17037 33152 17053 33216
rect 17117 33152 17125 33216
rect 16805 33151 17125 33152
rect 4909 32672 5229 32673
rect 4909 32608 4917 32672
rect 4981 32608 4997 32672
rect 5061 32608 5077 32672
rect 5141 32608 5157 32672
rect 5221 32608 5229 32672
rect 4909 32607 5229 32608
rect 12840 32672 13160 32673
rect 12840 32608 12848 32672
rect 12912 32608 12928 32672
rect 12992 32608 13008 32672
rect 13072 32608 13088 32672
rect 13152 32608 13160 32672
rect 12840 32607 13160 32608
rect 20770 32672 21090 32673
rect 20770 32608 20778 32672
rect 20842 32608 20858 32672
rect 20922 32608 20938 32672
rect 21002 32608 21018 32672
rect 21082 32608 21090 32672
rect 20770 32607 21090 32608
rect 8874 32128 9194 32129
rect 8874 32064 8882 32128
rect 8946 32064 8962 32128
rect 9026 32064 9042 32128
rect 9106 32064 9122 32128
rect 9186 32064 9194 32128
rect 8874 32063 9194 32064
rect 16805 32128 17125 32129
rect 16805 32064 16813 32128
rect 16877 32064 16893 32128
rect 16957 32064 16973 32128
rect 17037 32064 17053 32128
rect 17117 32064 17125 32128
rect 16805 32063 17125 32064
rect 5441 31652 5507 31653
rect 5390 31650 5396 31652
rect 5350 31590 5396 31650
rect 5460 31648 5507 31652
rect 5502 31592 5507 31648
rect 5390 31588 5396 31590
rect 5460 31588 5507 31592
rect 5441 31587 5507 31588
rect 4909 31584 5229 31585
rect 4909 31520 4917 31584
rect 4981 31520 4997 31584
rect 5061 31520 5077 31584
rect 5141 31520 5157 31584
rect 5221 31520 5229 31584
rect 4909 31519 5229 31520
rect 12840 31584 13160 31585
rect 12840 31520 12848 31584
rect 12912 31520 12928 31584
rect 12992 31520 13008 31584
rect 13072 31520 13088 31584
rect 13152 31520 13160 31584
rect 12840 31519 13160 31520
rect 20770 31584 21090 31585
rect 20770 31520 20778 31584
rect 20842 31520 20858 31584
rect 20922 31520 20938 31584
rect 21002 31520 21018 31584
rect 21082 31520 21090 31584
rect 20770 31519 21090 31520
rect 3141 31378 3207 31381
rect 4889 31378 4955 31381
rect 3141 31376 4955 31378
rect 3141 31320 3146 31376
rect 3202 31320 4894 31376
rect 4950 31320 4955 31376
rect 3141 31318 4955 31320
rect 3141 31315 3207 31318
rect 4889 31315 4955 31318
rect 8874 31040 9194 31041
rect 8874 30976 8882 31040
rect 8946 30976 8962 31040
rect 9026 30976 9042 31040
rect 9106 30976 9122 31040
rect 9186 30976 9194 31040
rect 8874 30975 9194 30976
rect 16805 31040 17125 31041
rect 16805 30976 16813 31040
rect 16877 30976 16893 31040
rect 16957 30976 16973 31040
rect 17037 30976 17053 31040
rect 17117 30976 17125 31040
rect 16805 30975 17125 30976
rect 0 30562 800 30592
rect 3509 30562 3575 30565
rect 0 30560 3575 30562
rect 0 30504 3514 30560
rect 3570 30504 3575 30560
rect 0 30502 3575 30504
rect 0 30472 800 30502
rect 3509 30499 3575 30502
rect 4909 30496 5229 30497
rect 4909 30432 4917 30496
rect 4981 30432 4997 30496
rect 5061 30432 5077 30496
rect 5141 30432 5157 30496
rect 5221 30432 5229 30496
rect 4909 30431 5229 30432
rect 12840 30496 13160 30497
rect 12840 30432 12848 30496
rect 12912 30432 12928 30496
rect 12992 30432 13008 30496
rect 13072 30432 13088 30496
rect 13152 30432 13160 30496
rect 12840 30431 13160 30432
rect 20770 30496 21090 30497
rect 20770 30432 20778 30496
rect 20842 30432 20858 30496
rect 20922 30432 20938 30496
rect 21002 30432 21018 30496
rect 21082 30432 21090 30496
rect 20770 30431 21090 30432
rect 8874 29952 9194 29953
rect 8874 29888 8882 29952
rect 8946 29888 8962 29952
rect 9026 29888 9042 29952
rect 9106 29888 9122 29952
rect 9186 29888 9194 29952
rect 8874 29887 9194 29888
rect 16805 29952 17125 29953
rect 16805 29888 16813 29952
rect 16877 29888 16893 29952
rect 16957 29888 16973 29952
rect 17037 29888 17053 29952
rect 17117 29888 17125 29952
rect 16805 29887 17125 29888
rect 4909 29408 5229 29409
rect 4909 29344 4917 29408
rect 4981 29344 4997 29408
rect 5061 29344 5077 29408
rect 5141 29344 5157 29408
rect 5221 29344 5229 29408
rect 4909 29343 5229 29344
rect 12840 29408 13160 29409
rect 12840 29344 12848 29408
rect 12912 29344 12928 29408
rect 12992 29344 13008 29408
rect 13072 29344 13088 29408
rect 13152 29344 13160 29408
rect 12840 29343 13160 29344
rect 20770 29408 21090 29409
rect 20770 29344 20778 29408
rect 20842 29344 20858 29408
rect 20922 29344 20938 29408
rect 21002 29344 21018 29408
rect 21082 29344 21090 29408
rect 20770 29343 21090 29344
rect 8874 28864 9194 28865
rect 8874 28800 8882 28864
rect 8946 28800 8962 28864
rect 9026 28800 9042 28864
rect 9106 28800 9122 28864
rect 9186 28800 9194 28864
rect 8874 28799 9194 28800
rect 16805 28864 17125 28865
rect 16805 28800 16813 28864
rect 16877 28800 16893 28864
rect 16957 28800 16973 28864
rect 17037 28800 17053 28864
rect 17117 28800 17125 28864
rect 16805 28799 17125 28800
rect 4153 28658 4219 28661
rect 4797 28658 4863 28661
rect 4153 28656 4863 28658
rect 4153 28600 4158 28656
rect 4214 28600 4802 28656
rect 4858 28600 4863 28656
rect 4153 28598 4863 28600
rect 4153 28595 4219 28598
rect 4478 28389 4538 28598
rect 4797 28595 4863 28598
rect 4797 28522 4863 28525
rect 4662 28520 4863 28522
rect 4662 28464 4802 28520
rect 4858 28464 4863 28520
rect 4662 28462 4863 28464
rect 4478 28384 4587 28389
rect 4478 28328 4526 28384
rect 4582 28328 4587 28384
rect 4478 28326 4587 28328
rect 4521 28323 4587 28326
rect 4662 28114 4722 28462
rect 4797 28459 4863 28462
rect 5073 28522 5139 28525
rect 8293 28524 8359 28525
rect 5390 28522 5396 28524
rect 5073 28520 5396 28522
rect 5073 28464 5078 28520
rect 5134 28464 5396 28520
rect 5073 28462 5396 28464
rect 5073 28459 5139 28462
rect 5390 28460 5396 28462
rect 5460 28460 5466 28524
rect 8293 28522 8340 28524
rect 8248 28520 8340 28522
rect 8248 28464 8298 28520
rect 8248 28462 8340 28464
rect 8293 28460 8340 28462
rect 8404 28460 8410 28524
rect 8293 28459 8359 28460
rect 4909 28320 5229 28321
rect 4909 28256 4917 28320
rect 4981 28256 4997 28320
rect 5061 28256 5077 28320
rect 5141 28256 5157 28320
rect 5221 28256 5229 28320
rect 4909 28255 5229 28256
rect 12840 28320 13160 28321
rect 12840 28256 12848 28320
rect 12912 28256 12928 28320
rect 12992 28256 13008 28320
rect 13072 28256 13088 28320
rect 13152 28256 13160 28320
rect 12840 28255 13160 28256
rect 20770 28320 21090 28321
rect 20770 28256 20778 28320
rect 20842 28256 20858 28320
rect 20922 28256 20938 28320
rect 21002 28256 21018 28320
rect 21082 28256 21090 28320
rect 20770 28255 21090 28256
rect 4889 28114 4955 28117
rect 4662 28112 4955 28114
rect 4662 28056 4894 28112
rect 4950 28056 4955 28112
rect 4662 28054 4955 28056
rect 4889 28051 4955 28054
rect 8874 27776 9194 27777
rect 8874 27712 8882 27776
rect 8946 27712 8962 27776
rect 9026 27712 9042 27776
rect 9106 27712 9122 27776
rect 9186 27712 9194 27776
rect 8874 27711 9194 27712
rect 16805 27776 17125 27777
rect 16805 27712 16813 27776
rect 16877 27712 16893 27776
rect 16957 27712 16973 27776
rect 17037 27712 17053 27776
rect 17117 27712 17125 27776
rect 16805 27711 17125 27712
rect 8477 27298 8543 27301
rect 9622 27298 9628 27300
rect 8477 27296 9628 27298
rect 8477 27240 8482 27296
rect 8538 27240 9628 27296
rect 8477 27238 9628 27240
rect 8477 27235 8543 27238
rect 9622 27236 9628 27238
rect 9692 27236 9698 27300
rect 4909 27232 5229 27233
rect 4909 27168 4917 27232
rect 4981 27168 4997 27232
rect 5061 27168 5077 27232
rect 5141 27168 5157 27232
rect 5221 27168 5229 27232
rect 4909 27167 5229 27168
rect 12840 27232 13160 27233
rect 12840 27168 12848 27232
rect 12912 27168 12928 27232
rect 12992 27168 13008 27232
rect 13072 27168 13088 27232
rect 13152 27168 13160 27232
rect 12840 27167 13160 27168
rect 20770 27232 21090 27233
rect 20770 27168 20778 27232
rect 20842 27168 20858 27232
rect 20922 27168 20938 27232
rect 21002 27168 21018 27232
rect 21082 27168 21090 27232
rect 20770 27167 21090 27168
rect 8293 27026 8359 27029
rect 8293 27024 8402 27026
rect 8293 26968 8298 27024
rect 8354 26968 8402 27024
rect 8293 26963 8402 26968
rect 8518 26964 8524 27028
rect 8588 27026 8594 27028
rect 8661 27026 8727 27029
rect 8588 27024 8727 27026
rect 8588 26968 8666 27024
rect 8722 26968 8727 27024
rect 8588 26966 8727 26968
rect 8588 26964 8594 26966
rect 8661 26963 8727 26966
rect 10174 26964 10180 27028
rect 10244 27026 10250 27028
rect 10777 27026 10843 27029
rect 10244 27024 10843 27026
rect 10244 26968 10782 27024
rect 10838 26968 10843 27024
rect 10244 26966 10843 26968
rect 10244 26964 10250 26966
rect 10777 26963 10843 26966
rect 8342 26890 8402 26963
rect 9673 26890 9739 26893
rect 8342 26888 9739 26890
rect 8342 26832 9678 26888
rect 9734 26832 9739 26888
rect 8342 26830 9739 26832
rect 9673 26827 9739 26830
rect 8293 26754 8359 26757
rect 8661 26756 8727 26757
rect 8661 26754 8708 26756
rect 8293 26752 8708 26754
rect 8293 26696 8298 26752
rect 8354 26696 8666 26752
rect 8293 26694 8708 26696
rect 8293 26691 8359 26694
rect 8661 26692 8708 26694
rect 8772 26692 8778 26756
rect 8661 26691 8727 26692
rect 8874 26688 9194 26689
rect 8874 26624 8882 26688
rect 8946 26624 8962 26688
rect 9026 26624 9042 26688
rect 9106 26624 9122 26688
rect 9186 26624 9194 26688
rect 8874 26623 9194 26624
rect 16805 26688 17125 26689
rect 16805 26624 16813 26688
rect 16877 26624 16893 26688
rect 16957 26624 16973 26688
rect 17037 26624 17053 26688
rect 17117 26624 17125 26688
rect 16805 26623 17125 26624
rect 2589 26482 2655 26485
rect 3785 26482 3851 26485
rect 2589 26480 3851 26482
rect 2589 26424 2594 26480
rect 2650 26424 3790 26480
rect 3846 26424 3851 26480
rect 2589 26422 3851 26424
rect 2589 26419 2655 26422
rect 3785 26419 3851 26422
rect 4909 26144 5229 26145
rect 4909 26080 4917 26144
rect 4981 26080 4997 26144
rect 5061 26080 5077 26144
rect 5141 26080 5157 26144
rect 5221 26080 5229 26144
rect 4909 26079 5229 26080
rect 12840 26144 13160 26145
rect 12840 26080 12848 26144
rect 12912 26080 12928 26144
rect 12992 26080 13008 26144
rect 13072 26080 13088 26144
rect 13152 26080 13160 26144
rect 12840 26079 13160 26080
rect 20770 26144 21090 26145
rect 20770 26080 20778 26144
rect 20842 26080 20858 26144
rect 20922 26080 20938 26144
rect 21002 26080 21018 26144
rect 21082 26080 21090 26144
rect 20770 26079 21090 26080
rect 9489 26076 9555 26077
rect 9438 26074 9444 26076
rect 9398 26014 9444 26074
rect 9508 26072 9555 26076
rect 9550 26016 9555 26072
rect 9438 26012 9444 26014
rect 9508 26012 9555 26016
rect 9489 26011 9555 26012
rect 8874 25600 9194 25601
rect 8874 25536 8882 25600
rect 8946 25536 8962 25600
rect 9026 25536 9042 25600
rect 9106 25536 9122 25600
rect 9186 25536 9194 25600
rect 8874 25535 9194 25536
rect 16805 25600 17125 25601
rect 16805 25536 16813 25600
rect 16877 25536 16893 25600
rect 16957 25536 16973 25600
rect 17037 25536 17053 25600
rect 17117 25536 17125 25600
rect 16805 25535 17125 25536
rect 4909 25056 5229 25057
rect 0 24986 800 25016
rect 4909 24992 4917 25056
rect 4981 24992 4997 25056
rect 5061 24992 5077 25056
rect 5141 24992 5157 25056
rect 5221 24992 5229 25056
rect 4909 24991 5229 24992
rect 12840 25056 13160 25057
rect 12840 24992 12848 25056
rect 12912 24992 12928 25056
rect 12992 24992 13008 25056
rect 13072 24992 13088 25056
rect 13152 24992 13160 25056
rect 12840 24991 13160 24992
rect 20770 25056 21090 25057
rect 20770 24992 20778 25056
rect 20842 24992 20858 25056
rect 20922 24992 20938 25056
rect 21002 24992 21018 25056
rect 21082 24992 21090 25056
rect 20770 24991 21090 24992
rect 4061 24986 4127 24989
rect 0 24984 4127 24986
rect 0 24928 4066 24984
rect 4122 24928 4127 24984
rect 0 24926 4127 24928
rect 0 24896 800 24926
rect 4061 24923 4127 24926
rect 9213 24852 9279 24853
rect 9213 24848 9260 24852
rect 9324 24850 9330 24852
rect 9213 24792 9218 24848
rect 9213 24788 9260 24792
rect 9324 24790 9370 24850
rect 9324 24788 9330 24790
rect 9213 24787 9279 24788
rect 9489 24714 9555 24717
rect 12617 24714 12683 24717
rect 9489 24712 12683 24714
rect 9489 24656 9494 24712
rect 9550 24656 12622 24712
rect 12678 24656 12683 24712
rect 9489 24654 12683 24656
rect 9489 24651 9555 24654
rect 12617 24651 12683 24654
rect 8874 24512 9194 24513
rect 8874 24448 8882 24512
rect 8946 24448 8962 24512
rect 9026 24448 9042 24512
rect 9106 24448 9122 24512
rect 9186 24448 9194 24512
rect 8874 24447 9194 24448
rect 16805 24512 17125 24513
rect 16805 24448 16813 24512
rect 16877 24448 16893 24512
rect 16957 24448 16973 24512
rect 17037 24448 17053 24512
rect 17117 24448 17125 24512
rect 16805 24447 17125 24448
rect 10133 24442 10199 24445
rect 11421 24442 11487 24445
rect 10133 24440 11487 24442
rect 10133 24384 10138 24440
rect 10194 24384 11426 24440
rect 11482 24384 11487 24440
rect 10133 24382 11487 24384
rect 10133 24379 10199 24382
rect 11421 24379 11487 24382
rect 8518 24244 8524 24308
rect 8588 24306 8594 24308
rect 10685 24306 10751 24309
rect 8588 24304 10751 24306
rect 8588 24248 10690 24304
rect 10746 24248 10751 24304
rect 8588 24246 10751 24248
rect 8588 24244 8594 24246
rect 10685 24243 10751 24246
rect 9765 24170 9831 24173
rect 10133 24170 10199 24173
rect 9765 24168 10199 24170
rect 9765 24112 9770 24168
rect 9826 24112 10138 24168
rect 10194 24112 10199 24168
rect 9765 24110 10199 24112
rect 9765 24107 9831 24110
rect 10133 24107 10199 24110
rect 9673 24034 9739 24037
rect 12617 24034 12683 24037
rect 9673 24032 12683 24034
rect 9673 23976 9678 24032
rect 9734 23976 12622 24032
rect 12678 23976 12683 24032
rect 9673 23974 12683 23976
rect 9673 23971 9739 23974
rect 12617 23971 12683 23974
rect 4909 23968 5229 23969
rect 4909 23904 4917 23968
rect 4981 23904 4997 23968
rect 5061 23904 5077 23968
rect 5141 23904 5157 23968
rect 5221 23904 5229 23968
rect 4909 23903 5229 23904
rect 12840 23968 13160 23969
rect 12840 23904 12848 23968
rect 12912 23904 12928 23968
rect 12992 23904 13008 23968
rect 13072 23904 13088 23968
rect 13152 23904 13160 23968
rect 12840 23903 13160 23904
rect 20770 23968 21090 23969
rect 20770 23904 20778 23968
rect 20842 23904 20858 23968
rect 20922 23904 20938 23968
rect 21002 23904 21018 23968
rect 21082 23904 21090 23968
rect 20770 23903 21090 23904
rect 9673 23762 9739 23765
rect 12433 23762 12499 23765
rect 9673 23760 14658 23762
rect 9673 23704 9678 23760
rect 9734 23704 12438 23760
rect 12494 23704 14658 23760
rect 9673 23702 14658 23704
rect 9673 23699 9739 23702
rect 12433 23699 12499 23702
rect 14598 23629 14658 23702
rect 14598 23626 14707 23629
rect 17953 23626 18019 23629
rect 14598 23624 18019 23626
rect 14598 23568 14646 23624
rect 14702 23568 17958 23624
rect 18014 23568 18019 23624
rect 14598 23566 18019 23568
rect 14641 23563 14707 23566
rect 17953 23563 18019 23566
rect 8874 23424 9194 23425
rect 8874 23360 8882 23424
rect 8946 23360 8962 23424
rect 9026 23360 9042 23424
rect 9106 23360 9122 23424
rect 9186 23360 9194 23424
rect 8874 23359 9194 23360
rect 16805 23424 17125 23425
rect 16805 23360 16813 23424
rect 16877 23360 16893 23424
rect 16957 23360 16973 23424
rect 17037 23360 17053 23424
rect 17117 23360 17125 23424
rect 16805 23359 17125 23360
rect 11237 23354 11303 23357
rect 12249 23354 12315 23357
rect 11237 23352 12315 23354
rect 11237 23296 11242 23352
rect 11298 23296 12254 23352
rect 12310 23296 12315 23352
rect 11237 23294 12315 23296
rect 11237 23291 11303 23294
rect 12249 23291 12315 23294
rect 11881 23218 11947 23221
rect 12065 23218 12131 23221
rect 12525 23218 12591 23221
rect 11881 23216 12591 23218
rect 11881 23160 11886 23216
rect 11942 23160 12070 23216
rect 12126 23160 12530 23216
rect 12586 23160 12591 23216
rect 11881 23158 12591 23160
rect 11881 23155 11947 23158
rect 12065 23155 12131 23158
rect 12525 23155 12591 23158
rect 5349 23084 5415 23085
rect 5349 23080 5396 23084
rect 5460 23082 5466 23084
rect 11421 23082 11487 23085
rect 12249 23082 12315 23085
rect 5349 23024 5354 23080
rect 5349 23020 5396 23024
rect 5460 23022 5506 23082
rect 11421 23080 12315 23082
rect 11421 23024 11426 23080
rect 11482 23024 12254 23080
rect 12310 23024 12315 23080
rect 11421 23022 12315 23024
rect 5460 23020 5466 23022
rect 5349 23019 5415 23020
rect 11421 23019 11487 23022
rect 12249 23019 12315 23022
rect 4909 22880 5229 22881
rect 4909 22816 4917 22880
rect 4981 22816 4997 22880
rect 5061 22816 5077 22880
rect 5141 22816 5157 22880
rect 5221 22816 5229 22880
rect 4909 22815 5229 22816
rect 12840 22880 13160 22881
rect 12840 22816 12848 22880
rect 12912 22816 12928 22880
rect 12992 22816 13008 22880
rect 13072 22816 13088 22880
rect 13152 22816 13160 22880
rect 12840 22815 13160 22816
rect 20770 22880 21090 22881
rect 20770 22816 20778 22880
rect 20842 22816 20858 22880
rect 20922 22816 20938 22880
rect 21002 22816 21018 22880
rect 21082 22816 21090 22880
rect 20770 22815 21090 22816
rect 7557 22810 7623 22813
rect 7925 22812 7991 22813
rect 7925 22810 7972 22812
rect 7557 22808 7972 22810
rect 8036 22810 8042 22812
rect 7557 22752 7562 22808
rect 7618 22752 7930 22808
rect 7557 22750 7972 22752
rect 7557 22747 7623 22750
rect 7925 22748 7972 22750
rect 8036 22750 8082 22810
rect 8036 22748 8042 22750
rect 7925 22747 7991 22748
rect 8477 22676 8543 22677
rect 8477 22674 8524 22676
rect 8432 22672 8524 22674
rect 8432 22616 8482 22672
rect 8432 22614 8524 22616
rect 8477 22612 8524 22614
rect 8588 22612 8594 22676
rect 8477 22611 8543 22612
rect 1669 22538 1735 22541
rect 8334 22538 8340 22540
rect 1669 22536 8340 22538
rect 1669 22480 1674 22536
rect 1730 22480 8340 22536
rect 1669 22478 8340 22480
rect 1669 22475 1735 22478
rect 8334 22476 8340 22478
rect 8404 22476 8410 22540
rect 6821 22402 6887 22405
rect 7189 22402 7255 22405
rect 6821 22400 7255 22402
rect 6821 22344 6826 22400
rect 6882 22344 7194 22400
rect 7250 22344 7255 22400
rect 6821 22342 7255 22344
rect 6821 22339 6887 22342
rect 7189 22339 7255 22342
rect 8874 22336 9194 22337
rect 8874 22272 8882 22336
rect 8946 22272 8962 22336
rect 9026 22272 9042 22336
rect 9106 22272 9122 22336
rect 9186 22272 9194 22336
rect 8874 22271 9194 22272
rect 16805 22336 17125 22337
rect 16805 22272 16813 22336
rect 16877 22272 16893 22336
rect 16957 22272 16973 22336
rect 17037 22272 17053 22336
rect 17117 22272 17125 22336
rect 16805 22271 17125 22272
rect 8201 22130 8267 22133
rect 11329 22130 11395 22133
rect 8201 22128 11395 22130
rect 8201 22072 8206 22128
rect 8262 22072 11334 22128
rect 11390 22072 11395 22128
rect 8201 22070 11395 22072
rect 8201 22067 8267 22070
rect 11329 22067 11395 22070
rect 7046 21932 7052 21996
rect 7116 21994 7122 21996
rect 7465 21994 7531 21997
rect 9489 21996 9555 21997
rect 9438 21994 9444 21996
rect 7116 21992 7531 21994
rect 7116 21936 7470 21992
rect 7526 21936 7531 21992
rect 7116 21934 7531 21936
rect 9398 21934 9444 21994
rect 9508 21992 9555 21996
rect 9550 21936 9555 21992
rect 7116 21932 7122 21934
rect 7465 21931 7531 21934
rect 9438 21932 9444 21934
rect 9508 21932 9555 21936
rect 9489 21931 9555 21932
rect 7465 21858 7531 21861
rect 7966 21858 7972 21860
rect 7465 21856 7972 21858
rect 7465 21800 7470 21856
rect 7526 21800 7972 21856
rect 7465 21798 7972 21800
rect 7465 21795 7531 21798
rect 7966 21796 7972 21798
rect 8036 21796 8042 21860
rect 4909 21792 5229 21793
rect 4909 21728 4917 21792
rect 4981 21728 4997 21792
rect 5061 21728 5077 21792
rect 5141 21728 5157 21792
rect 5221 21728 5229 21792
rect 4909 21727 5229 21728
rect 12840 21792 13160 21793
rect 12840 21728 12848 21792
rect 12912 21728 12928 21792
rect 12992 21728 13008 21792
rect 13072 21728 13088 21792
rect 13152 21728 13160 21792
rect 12840 21727 13160 21728
rect 20770 21792 21090 21793
rect 20770 21728 20778 21792
rect 20842 21728 20858 21792
rect 20922 21728 20938 21792
rect 21002 21728 21018 21792
rect 21082 21728 21090 21792
rect 20770 21727 21090 21728
rect 7414 21660 7420 21724
rect 7484 21722 7490 21724
rect 7557 21722 7623 21725
rect 7484 21720 7623 21722
rect 7484 21664 7562 21720
rect 7618 21664 7623 21720
rect 7484 21662 7623 21664
rect 7484 21660 7490 21662
rect 7557 21659 7623 21662
rect 4245 21586 4311 21589
rect 6545 21586 6611 21589
rect 4245 21584 4354 21586
rect 4245 21528 4250 21584
rect 4306 21528 4354 21584
rect 4245 21523 4354 21528
rect 6545 21584 6746 21586
rect 6545 21528 6550 21584
rect 6606 21528 6746 21584
rect 6545 21526 6746 21528
rect 6545 21523 6611 21526
rect 4294 20909 4354 21523
rect 4294 20904 4403 20909
rect 4294 20848 4342 20904
rect 4398 20848 4403 20904
rect 4294 20846 4403 20848
rect 4337 20843 4403 20846
rect 6686 20770 6746 21526
rect 6862 21524 6868 21588
rect 6932 21586 6938 21588
rect 7741 21586 7807 21589
rect 9581 21586 9647 21589
rect 6932 21584 7807 21586
rect 6932 21528 7746 21584
rect 7802 21528 7807 21584
rect 6932 21526 7807 21528
rect 6932 21524 6938 21526
rect 7741 21523 7807 21526
rect 9262 21584 9647 21586
rect 9262 21528 9586 21584
rect 9642 21528 9647 21584
rect 9262 21526 9647 21528
rect 9262 21453 9322 21526
rect 9581 21523 9647 21526
rect 11145 21586 11211 21589
rect 18321 21586 18387 21589
rect 11145 21584 18387 21586
rect 11145 21528 11150 21584
rect 11206 21528 18326 21584
rect 18382 21528 18387 21584
rect 11145 21526 18387 21528
rect 11145 21523 11211 21526
rect 18321 21523 18387 21526
rect 9213 21448 9322 21453
rect 9213 21392 9218 21448
rect 9274 21392 9322 21448
rect 9213 21390 9322 21392
rect 11145 21450 11211 21453
rect 14089 21450 14155 21453
rect 17217 21450 17283 21453
rect 11145 21448 17283 21450
rect 11145 21392 11150 21448
rect 11206 21392 14094 21448
rect 14150 21392 17222 21448
rect 17278 21392 17283 21448
rect 11145 21390 17283 21392
rect 9213 21387 9279 21390
rect 11145 21387 11211 21390
rect 14089 21387 14155 21390
rect 17217 21387 17283 21390
rect 8874 21248 9194 21249
rect 8874 21184 8882 21248
rect 8946 21184 8962 21248
rect 9026 21184 9042 21248
rect 9106 21184 9122 21248
rect 9186 21184 9194 21248
rect 8874 21183 9194 21184
rect 16805 21248 17125 21249
rect 16805 21184 16813 21248
rect 16877 21184 16893 21248
rect 16957 21184 16973 21248
rect 17037 21184 17053 21248
rect 17117 21184 17125 21248
rect 16805 21183 17125 21184
rect 8702 20980 8708 21044
rect 8772 21042 8778 21044
rect 9121 21042 9187 21045
rect 8772 21040 9187 21042
rect 8772 20984 9126 21040
rect 9182 20984 9187 21040
rect 8772 20982 9187 20984
rect 8772 20980 8778 20982
rect 9121 20979 9187 20982
rect 6821 20770 6887 20773
rect 8385 20772 8451 20773
rect 8334 20770 8340 20772
rect 6686 20768 6887 20770
rect 6686 20712 6826 20768
rect 6882 20712 6887 20768
rect 6686 20710 6887 20712
rect 8294 20710 8340 20770
rect 8404 20768 8451 20772
rect 8446 20712 8451 20768
rect 6821 20707 6887 20710
rect 8334 20708 8340 20710
rect 8404 20708 8451 20712
rect 8385 20707 8451 20708
rect 4909 20704 5229 20705
rect 4909 20640 4917 20704
rect 4981 20640 4997 20704
rect 5061 20640 5077 20704
rect 5141 20640 5157 20704
rect 5221 20640 5229 20704
rect 4909 20639 5229 20640
rect 12840 20704 13160 20705
rect 12840 20640 12848 20704
rect 12912 20640 12928 20704
rect 12992 20640 13008 20704
rect 13072 20640 13088 20704
rect 13152 20640 13160 20704
rect 12840 20639 13160 20640
rect 20770 20704 21090 20705
rect 20770 20640 20778 20704
rect 20842 20640 20858 20704
rect 20922 20640 20938 20704
rect 21002 20640 21018 20704
rect 21082 20640 21090 20704
rect 20770 20639 21090 20640
rect 8845 20498 8911 20501
rect 9254 20498 9260 20500
rect 8845 20496 9260 20498
rect 8845 20440 8850 20496
rect 8906 20440 9260 20496
rect 8845 20438 9260 20440
rect 8845 20435 8911 20438
rect 9254 20436 9260 20438
rect 9324 20436 9330 20500
rect 8874 20160 9194 20161
rect 8874 20096 8882 20160
rect 8946 20096 8962 20160
rect 9026 20096 9042 20160
rect 9106 20096 9122 20160
rect 9186 20096 9194 20160
rect 8874 20095 9194 20096
rect 16805 20160 17125 20161
rect 16805 20096 16813 20160
rect 16877 20096 16893 20160
rect 16957 20096 16973 20160
rect 17037 20096 17053 20160
rect 17117 20096 17125 20160
rect 16805 20095 17125 20096
rect 6913 19954 6979 19957
rect 7046 19954 7052 19956
rect 6913 19952 7052 19954
rect 6913 19896 6918 19952
rect 6974 19896 7052 19952
rect 6913 19894 7052 19896
rect 6913 19891 6979 19894
rect 7046 19892 7052 19894
rect 7116 19892 7122 19956
rect 8385 19818 8451 19821
rect 9622 19818 9628 19820
rect 8385 19816 9628 19818
rect 8385 19760 8390 19816
rect 8446 19760 9628 19816
rect 8385 19758 9628 19760
rect 8385 19755 8451 19758
rect 9622 19756 9628 19758
rect 9692 19756 9698 19820
rect 4909 19616 5229 19617
rect 4909 19552 4917 19616
rect 4981 19552 4997 19616
rect 5061 19552 5077 19616
rect 5141 19552 5157 19616
rect 5221 19552 5229 19616
rect 4909 19551 5229 19552
rect 12840 19616 13160 19617
rect 12840 19552 12848 19616
rect 12912 19552 12928 19616
rect 12992 19552 13008 19616
rect 13072 19552 13088 19616
rect 13152 19552 13160 19616
rect 12840 19551 13160 19552
rect 20770 19616 21090 19617
rect 20770 19552 20778 19616
rect 20842 19552 20858 19616
rect 20922 19552 20938 19616
rect 21002 19552 21018 19616
rect 21082 19552 21090 19616
rect 20770 19551 21090 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 3417 19410 3483 19413
rect 4981 19410 5047 19413
rect 6862 19410 6868 19412
rect 3417 19408 6868 19410
rect 3417 19352 3422 19408
rect 3478 19352 4986 19408
rect 5042 19352 6868 19408
rect 3417 19350 6868 19352
rect 3417 19347 3483 19350
rect 4981 19347 5047 19350
rect 6862 19348 6868 19350
rect 6932 19348 6938 19412
rect 9949 19138 10015 19141
rect 10174 19138 10180 19140
rect 9949 19136 10180 19138
rect 9949 19080 9954 19136
rect 10010 19080 10180 19136
rect 9949 19078 10180 19080
rect 9949 19075 10015 19078
rect 10174 19076 10180 19078
rect 10244 19076 10250 19140
rect 8874 19072 9194 19073
rect 8874 19008 8882 19072
rect 8946 19008 8962 19072
rect 9026 19008 9042 19072
rect 9106 19008 9122 19072
rect 9186 19008 9194 19072
rect 8874 19007 9194 19008
rect 16805 19072 17125 19073
rect 16805 19008 16813 19072
rect 16877 19008 16893 19072
rect 16957 19008 16973 19072
rect 17037 19008 17053 19072
rect 17117 19008 17125 19072
rect 16805 19007 17125 19008
rect 7373 19004 7439 19005
rect 7373 19000 7420 19004
rect 7484 19002 7490 19004
rect 7373 18944 7378 19000
rect 7373 18940 7420 18944
rect 7484 18942 7530 19002
rect 7484 18940 7490 18942
rect 7373 18939 7439 18940
rect 4981 18730 5047 18733
rect 5390 18730 5396 18732
rect 4981 18728 5396 18730
rect 4981 18672 4986 18728
rect 5042 18672 5396 18728
rect 4981 18670 5396 18672
rect 4981 18667 5047 18670
rect 5390 18668 5396 18670
rect 5460 18668 5466 18732
rect 4909 18528 5229 18529
rect 4909 18464 4917 18528
rect 4981 18464 4997 18528
rect 5061 18464 5077 18528
rect 5141 18464 5157 18528
rect 5221 18464 5229 18528
rect 4909 18463 5229 18464
rect 12840 18528 13160 18529
rect 12840 18464 12848 18528
rect 12912 18464 12928 18528
rect 12992 18464 13008 18528
rect 13072 18464 13088 18528
rect 13152 18464 13160 18528
rect 12840 18463 13160 18464
rect 20770 18528 21090 18529
rect 20770 18464 20778 18528
rect 20842 18464 20858 18528
rect 20922 18464 20938 18528
rect 21002 18464 21018 18528
rect 21082 18464 21090 18528
rect 20770 18463 21090 18464
rect 8874 17984 9194 17985
rect 8874 17920 8882 17984
rect 8946 17920 8962 17984
rect 9026 17920 9042 17984
rect 9106 17920 9122 17984
rect 9186 17920 9194 17984
rect 8874 17919 9194 17920
rect 16805 17984 17125 17985
rect 16805 17920 16813 17984
rect 16877 17920 16893 17984
rect 16957 17920 16973 17984
rect 17037 17920 17053 17984
rect 17117 17920 17125 17984
rect 16805 17919 17125 17920
rect 4909 17440 5229 17441
rect 4909 17376 4917 17440
rect 4981 17376 4997 17440
rect 5061 17376 5077 17440
rect 5141 17376 5157 17440
rect 5221 17376 5229 17440
rect 4909 17375 5229 17376
rect 12840 17440 13160 17441
rect 12840 17376 12848 17440
rect 12912 17376 12928 17440
rect 12992 17376 13008 17440
rect 13072 17376 13088 17440
rect 13152 17376 13160 17440
rect 12840 17375 13160 17376
rect 20770 17440 21090 17441
rect 20770 17376 20778 17440
rect 20842 17376 20858 17440
rect 20922 17376 20938 17440
rect 21002 17376 21018 17440
rect 21082 17376 21090 17440
rect 20770 17375 21090 17376
rect 8874 16896 9194 16897
rect 8874 16832 8882 16896
rect 8946 16832 8962 16896
rect 9026 16832 9042 16896
rect 9106 16832 9122 16896
rect 9186 16832 9194 16896
rect 8874 16831 9194 16832
rect 16805 16896 17125 16897
rect 16805 16832 16813 16896
rect 16877 16832 16893 16896
rect 16957 16832 16973 16896
rect 17037 16832 17053 16896
rect 17117 16832 17125 16896
rect 16805 16831 17125 16832
rect 10133 16690 10199 16693
rect 15561 16690 15627 16693
rect 10133 16688 15627 16690
rect 10133 16632 10138 16688
rect 10194 16632 15566 16688
rect 15622 16632 15627 16688
rect 10133 16630 15627 16632
rect 10133 16627 10199 16630
rect 15561 16627 15627 16630
rect 4909 16352 5229 16353
rect 4909 16288 4917 16352
rect 4981 16288 4997 16352
rect 5061 16288 5077 16352
rect 5141 16288 5157 16352
rect 5221 16288 5229 16352
rect 4909 16287 5229 16288
rect 12840 16352 13160 16353
rect 12840 16288 12848 16352
rect 12912 16288 12928 16352
rect 12992 16288 13008 16352
rect 13072 16288 13088 16352
rect 13152 16288 13160 16352
rect 12840 16287 13160 16288
rect 20770 16352 21090 16353
rect 20770 16288 20778 16352
rect 20842 16288 20858 16352
rect 20922 16288 20938 16352
rect 21002 16288 21018 16352
rect 21082 16288 21090 16352
rect 20770 16287 21090 16288
rect 8874 15808 9194 15809
rect 8874 15744 8882 15808
rect 8946 15744 8962 15808
rect 9026 15744 9042 15808
rect 9106 15744 9122 15808
rect 9186 15744 9194 15808
rect 8874 15743 9194 15744
rect 16805 15808 17125 15809
rect 16805 15744 16813 15808
rect 16877 15744 16893 15808
rect 16957 15744 16973 15808
rect 17037 15744 17053 15808
rect 17117 15744 17125 15808
rect 16805 15743 17125 15744
rect 4909 15264 5229 15265
rect 4909 15200 4917 15264
rect 4981 15200 4997 15264
rect 5061 15200 5077 15264
rect 5141 15200 5157 15264
rect 5221 15200 5229 15264
rect 4909 15199 5229 15200
rect 12840 15264 13160 15265
rect 12840 15200 12848 15264
rect 12912 15200 12928 15264
rect 12992 15200 13008 15264
rect 13072 15200 13088 15264
rect 13152 15200 13160 15264
rect 12840 15199 13160 15200
rect 20770 15264 21090 15265
rect 20770 15200 20778 15264
rect 20842 15200 20858 15264
rect 20922 15200 20938 15264
rect 21002 15200 21018 15264
rect 21082 15200 21090 15264
rect 20770 15199 21090 15200
rect 8874 14720 9194 14721
rect 8874 14656 8882 14720
rect 8946 14656 8962 14720
rect 9026 14656 9042 14720
rect 9106 14656 9122 14720
rect 9186 14656 9194 14720
rect 8874 14655 9194 14656
rect 16805 14720 17125 14721
rect 16805 14656 16813 14720
rect 16877 14656 16893 14720
rect 16957 14656 16973 14720
rect 17037 14656 17053 14720
rect 17117 14656 17125 14720
rect 16805 14655 17125 14656
rect 4909 14176 5229 14177
rect 4909 14112 4917 14176
rect 4981 14112 4997 14176
rect 5061 14112 5077 14176
rect 5141 14112 5157 14176
rect 5221 14112 5229 14176
rect 4909 14111 5229 14112
rect 12840 14176 13160 14177
rect 12840 14112 12848 14176
rect 12912 14112 12928 14176
rect 12992 14112 13008 14176
rect 13072 14112 13088 14176
rect 13152 14112 13160 14176
rect 12840 14111 13160 14112
rect 20770 14176 21090 14177
rect 20770 14112 20778 14176
rect 20842 14112 20858 14176
rect 20922 14112 20938 14176
rect 21002 14112 21018 14176
rect 21082 14112 21090 14176
rect 20770 14111 21090 14112
rect 0 13834 800 13864
rect 5441 13834 5507 13837
rect 0 13832 5507 13834
rect 0 13776 5446 13832
rect 5502 13776 5507 13832
rect 0 13774 5507 13776
rect 0 13744 800 13774
rect 5441 13771 5507 13774
rect 8874 13632 9194 13633
rect 8874 13568 8882 13632
rect 8946 13568 8962 13632
rect 9026 13568 9042 13632
rect 9106 13568 9122 13632
rect 9186 13568 9194 13632
rect 8874 13567 9194 13568
rect 16805 13632 17125 13633
rect 16805 13568 16813 13632
rect 16877 13568 16893 13632
rect 16957 13568 16973 13632
rect 17037 13568 17053 13632
rect 17117 13568 17125 13632
rect 16805 13567 17125 13568
rect 9397 13156 9463 13157
rect 9397 13154 9444 13156
rect 9352 13152 9444 13154
rect 9352 13096 9402 13152
rect 9352 13094 9444 13096
rect 9397 13092 9444 13094
rect 9508 13092 9514 13156
rect 9397 13091 9463 13092
rect 4909 13088 5229 13089
rect 4909 13024 4917 13088
rect 4981 13024 4997 13088
rect 5061 13024 5077 13088
rect 5141 13024 5157 13088
rect 5221 13024 5229 13088
rect 4909 13023 5229 13024
rect 12840 13088 13160 13089
rect 12840 13024 12848 13088
rect 12912 13024 12928 13088
rect 12992 13024 13008 13088
rect 13072 13024 13088 13088
rect 13152 13024 13160 13088
rect 12840 13023 13160 13024
rect 20770 13088 21090 13089
rect 20770 13024 20778 13088
rect 20842 13024 20858 13088
rect 20922 13024 20938 13088
rect 21002 13024 21018 13088
rect 21082 13024 21090 13088
rect 20770 13023 21090 13024
rect 5165 12882 5231 12885
rect 5390 12882 5396 12884
rect 5165 12880 5396 12882
rect 5165 12824 5170 12880
rect 5226 12824 5396 12880
rect 5165 12822 5396 12824
rect 5165 12819 5231 12822
rect 5390 12820 5396 12822
rect 5460 12820 5466 12884
rect 8874 12544 9194 12545
rect 8874 12480 8882 12544
rect 8946 12480 8962 12544
rect 9026 12480 9042 12544
rect 9106 12480 9122 12544
rect 9186 12480 9194 12544
rect 8874 12479 9194 12480
rect 16805 12544 17125 12545
rect 16805 12480 16813 12544
rect 16877 12480 16893 12544
rect 16957 12480 16973 12544
rect 17037 12480 17053 12544
rect 17117 12480 17125 12544
rect 16805 12479 17125 12480
rect 8201 12474 8267 12477
rect 8158 12472 8267 12474
rect 8158 12416 8206 12472
rect 8262 12416 8267 12472
rect 8158 12411 8267 12416
rect 8158 12341 8218 12411
rect 8158 12336 8267 12341
rect 8158 12280 8206 12336
rect 8262 12280 8267 12336
rect 8158 12278 8267 12280
rect 8201 12275 8267 12278
rect 4909 12000 5229 12001
rect 4909 11936 4917 12000
rect 4981 11936 4997 12000
rect 5061 11936 5077 12000
rect 5141 11936 5157 12000
rect 5221 11936 5229 12000
rect 4909 11935 5229 11936
rect 12840 12000 13160 12001
rect 12840 11936 12848 12000
rect 12912 11936 12928 12000
rect 12992 11936 13008 12000
rect 13072 11936 13088 12000
rect 13152 11936 13160 12000
rect 12840 11935 13160 11936
rect 20770 12000 21090 12001
rect 20770 11936 20778 12000
rect 20842 11936 20858 12000
rect 20922 11936 20938 12000
rect 21002 11936 21018 12000
rect 21082 11936 21090 12000
rect 20770 11935 21090 11936
rect 8874 11456 9194 11457
rect 8874 11392 8882 11456
rect 8946 11392 8962 11456
rect 9026 11392 9042 11456
rect 9106 11392 9122 11456
rect 9186 11392 9194 11456
rect 8874 11391 9194 11392
rect 16805 11456 17125 11457
rect 16805 11392 16813 11456
rect 16877 11392 16893 11456
rect 16957 11392 16973 11456
rect 17037 11392 17053 11456
rect 17117 11392 17125 11456
rect 16805 11391 17125 11392
rect 12709 11250 12775 11253
rect 12436 11248 12775 11250
rect 12436 11192 12714 11248
rect 12770 11192 12775 11248
rect 12436 11190 12775 11192
rect 12436 10981 12496 11190
rect 12709 11187 12775 11190
rect 12433 10976 12499 10981
rect 12433 10920 12438 10976
rect 12494 10920 12499 10976
rect 12433 10915 12499 10920
rect 4909 10912 5229 10913
rect 4909 10848 4917 10912
rect 4981 10848 4997 10912
rect 5061 10848 5077 10912
rect 5141 10848 5157 10912
rect 5221 10848 5229 10912
rect 4909 10847 5229 10848
rect 12840 10912 13160 10913
rect 12840 10848 12848 10912
rect 12912 10848 12928 10912
rect 12992 10848 13008 10912
rect 13072 10848 13088 10912
rect 13152 10848 13160 10912
rect 12840 10847 13160 10848
rect 20770 10912 21090 10913
rect 20770 10848 20778 10912
rect 20842 10848 20858 10912
rect 20922 10848 20938 10912
rect 21002 10848 21018 10912
rect 21082 10848 21090 10912
rect 20770 10847 21090 10848
rect 12341 10706 12407 10709
rect 19149 10706 19215 10709
rect 12341 10704 19215 10706
rect 12341 10648 12346 10704
rect 12402 10648 19154 10704
rect 19210 10648 19215 10704
rect 12341 10646 19215 10648
rect 12341 10643 12407 10646
rect 19149 10643 19215 10646
rect 8874 10368 9194 10369
rect 8874 10304 8882 10368
rect 8946 10304 8962 10368
rect 9026 10304 9042 10368
rect 9106 10304 9122 10368
rect 9186 10304 9194 10368
rect 8874 10303 9194 10304
rect 16805 10368 17125 10369
rect 16805 10304 16813 10368
rect 16877 10304 16893 10368
rect 16957 10304 16973 10368
rect 17037 10304 17053 10368
rect 17117 10304 17125 10368
rect 16805 10303 17125 10304
rect 7097 10298 7163 10301
rect 7230 10298 7236 10300
rect 7097 10296 7236 10298
rect 7097 10240 7102 10296
rect 7158 10240 7236 10296
rect 7097 10238 7236 10240
rect 7097 10235 7163 10238
rect 7230 10236 7236 10238
rect 7300 10236 7306 10300
rect 2037 10026 2103 10029
rect 20897 10026 20963 10029
rect 2037 10024 20963 10026
rect 2037 9968 2042 10024
rect 2098 9968 20902 10024
rect 20958 9968 20963 10024
rect 2037 9966 20963 9968
rect 2037 9963 2103 9966
rect 20897 9963 20963 9966
rect 12198 9828 12204 9892
rect 12268 9890 12274 9892
rect 12433 9890 12499 9893
rect 12268 9888 12499 9890
rect 12268 9832 12438 9888
rect 12494 9832 12499 9888
rect 12268 9830 12499 9832
rect 12268 9828 12274 9830
rect 12433 9827 12499 9830
rect 4909 9824 5229 9825
rect 4909 9760 4917 9824
rect 4981 9760 4997 9824
rect 5061 9760 5077 9824
rect 5141 9760 5157 9824
rect 5221 9760 5229 9824
rect 4909 9759 5229 9760
rect 12840 9824 13160 9825
rect 12840 9760 12848 9824
rect 12912 9760 12928 9824
rect 12992 9760 13008 9824
rect 13072 9760 13088 9824
rect 13152 9760 13160 9824
rect 12840 9759 13160 9760
rect 20770 9824 21090 9825
rect 20770 9760 20778 9824
rect 20842 9760 20858 9824
rect 20922 9760 20938 9824
rect 21002 9760 21018 9824
rect 21082 9760 21090 9824
rect 20770 9759 21090 9760
rect 4889 9618 4955 9621
rect 5901 9618 5967 9621
rect 4889 9616 5967 9618
rect 4889 9560 4894 9616
rect 4950 9560 5906 9616
rect 5962 9560 5967 9616
rect 4889 9558 5967 9560
rect 4889 9555 4955 9558
rect 5901 9555 5967 9558
rect 6085 9618 6151 9621
rect 10961 9618 11027 9621
rect 6085 9616 11027 9618
rect 6085 9560 6090 9616
rect 6146 9560 10966 9616
rect 11022 9560 11027 9616
rect 6085 9558 11027 9560
rect 6085 9555 6151 9558
rect 10961 9555 11027 9558
rect 5165 9482 5231 9485
rect 5625 9482 5691 9485
rect 5165 9480 5691 9482
rect 5165 9424 5170 9480
rect 5226 9424 5630 9480
rect 5686 9424 5691 9480
rect 5165 9422 5691 9424
rect 5165 9419 5231 9422
rect 5625 9419 5691 9422
rect 10961 9482 11027 9485
rect 18229 9482 18295 9485
rect 10961 9480 18295 9482
rect 10961 9424 10966 9480
rect 11022 9424 18234 9480
rect 18290 9424 18295 9480
rect 10961 9422 18295 9424
rect 10961 9419 11027 9422
rect 18229 9419 18295 9422
rect 11513 9346 11579 9349
rect 12893 9346 12959 9349
rect 13302 9346 13308 9348
rect 11513 9344 13308 9346
rect 11513 9288 11518 9344
rect 11574 9288 12898 9344
rect 12954 9288 13308 9344
rect 11513 9286 13308 9288
rect 11513 9283 11579 9286
rect 12893 9283 12959 9286
rect 13302 9284 13308 9286
rect 13372 9346 13378 9348
rect 16481 9346 16547 9349
rect 13372 9344 16547 9346
rect 13372 9288 16486 9344
rect 16542 9288 16547 9344
rect 13372 9286 16547 9288
rect 13372 9284 13378 9286
rect 16481 9283 16547 9286
rect 8874 9280 9194 9281
rect 8874 9216 8882 9280
rect 8946 9216 8962 9280
rect 9026 9216 9042 9280
rect 9106 9216 9122 9280
rect 9186 9216 9194 9280
rect 8874 9215 9194 9216
rect 16805 9280 17125 9281
rect 16805 9216 16813 9280
rect 16877 9216 16893 9280
rect 16957 9216 16973 9280
rect 17037 9216 17053 9280
rect 17117 9216 17125 9280
rect 16805 9215 17125 9216
rect 10777 9210 10843 9213
rect 14733 9210 14799 9213
rect 10777 9208 14799 9210
rect 10777 9152 10782 9208
rect 10838 9152 14738 9208
rect 14794 9152 14799 9208
rect 10777 9150 14799 9152
rect 10777 9147 10843 9150
rect 14733 9147 14799 9150
rect 4429 9074 4495 9077
rect 5390 9074 5396 9076
rect 4429 9072 5396 9074
rect 4429 9016 4434 9072
rect 4490 9016 5396 9072
rect 4429 9014 5396 9016
rect 4429 9011 4495 9014
rect 5390 9012 5396 9014
rect 5460 9012 5466 9076
rect 8293 9074 8359 9077
rect 12433 9074 12499 9077
rect 8293 9072 12499 9074
rect 8293 9016 8298 9072
rect 8354 9016 12438 9072
rect 12494 9016 12499 9072
rect 8293 9014 12499 9016
rect 8293 9011 8359 9014
rect 12433 9011 12499 9014
rect 12566 9012 12572 9076
rect 12636 9074 12642 9076
rect 17493 9074 17559 9077
rect 12636 9072 17559 9074
rect 12636 9016 17498 9072
rect 17554 9016 17559 9072
rect 12636 9014 17559 9016
rect 12636 9012 12642 9014
rect 17493 9011 17559 9014
rect 10961 8938 11027 8941
rect 12249 8938 12315 8941
rect 15285 8938 15351 8941
rect 10961 8936 15351 8938
rect 10961 8880 10966 8936
rect 11022 8880 12254 8936
rect 12310 8880 15290 8936
rect 15346 8880 15351 8936
rect 10961 8878 15351 8880
rect 10961 8875 11027 8878
rect 12249 8875 12315 8878
rect 15285 8875 15351 8878
rect 4909 8736 5229 8737
rect 4909 8672 4917 8736
rect 4981 8672 4997 8736
rect 5061 8672 5077 8736
rect 5141 8672 5157 8736
rect 5221 8672 5229 8736
rect 4909 8671 5229 8672
rect 12840 8736 13160 8737
rect 12840 8672 12848 8736
rect 12912 8672 12928 8736
rect 12992 8672 13008 8736
rect 13072 8672 13088 8736
rect 13152 8672 13160 8736
rect 12840 8671 13160 8672
rect 20770 8736 21090 8737
rect 20770 8672 20778 8736
rect 20842 8672 20858 8736
rect 20922 8672 20938 8736
rect 21002 8672 21018 8736
rect 21082 8672 21090 8736
rect 20770 8671 21090 8672
rect 4429 8530 4495 8533
rect 12566 8530 12572 8532
rect 4429 8528 12572 8530
rect 4429 8472 4434 8528
rect 4490 8472 12572 8528
rect 4429 8470 12572 8472
rect 4429 8467 4495 8470
rect 12566 8468 12572 8470
rect 12636 8468 12642 8532
rect 10409 8394 10475 8397
rect 12433 8394 12499 8397
rect 10409 8392 12499 8394
rect 10409 8336 10414 8392
rect 10470 8336 12438 8392
rect 12494 8336 12499 8392
rect 10409 8334 12499 8336
rect 10409 8331 10475 8334
rect 12433 8331 12499 8334
rect 13077 8394 13143 8397
rect 13302 8394 13308 8396
rect 13077 8392 13308 8394
rect 13077 8336 13082 8392
rect 13138 8336 13308 8392
rect 13077 8334 13308 8336
rect 13077 8331 13143 8334
rect 13302 8332 13308 8334
rect 13372 8332 13378 8396
rect 0 8258 800 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 800 8198
rect 4061 8195 4127 8198
rect 13169 8258 13235 8261
rect 13486 8258 13492 8260
rect 13169 8256 13492 8258
rect 13169 8200 13174 8256
rect 13230 8200 13492 8256
rect 13169 8198 13492 8200
rect 13169 8195 13235 8198
rect 13486 8196 13492 8198
rect 13556 8196 13562 8260
rect 8874 8192 9194 8193
rect 8874 8128 8882 8192
rect 8946 8128 8962 8192
rect 9026 8128 9042 8192
rect 9106 8128 9122 8192
rect 9186 8128 9194 8192
rect 8874 8127 9194 8128
rect 16805 8192 17125 8193
rect 16805 8128 16813 8192
rect 16877 8128 16893 8192
rect 16957 8128 16973 8192
rect 17037 8128 17053 8192
rect 17117 8128 17125 8192
rect 16805 8127 17125 8128
rect 12893 8122 12959 8125
rect 13445 8122 13511 8125
rect 12893 8120 13511 8122
rect 12893 8064 12898 8120
rect 12954 8064 13450 8120
rect 13506 8064 13511 8120
rect 12893 8062 13511 8064
rect 12893 8059 12959 8062
rect 13445 8059 13511 8062
rect 10961 7986 11027 7989
rect 14365 7986 14431 7989
rect 10961 7984 14431 7986
rect 10961 7928 10966 7984
rect 11022 7928 14370 7984
rect 14426 7928 14431 7984
rect 10961 7926 14431 7928
rect 10961 7923 11027 7926
rect 14365 7923 14431 7926
rect 7281 7852 7347 7853
rect 7230 7788 7236 7852
rect 7300 7850 7347 7852
rect 12157 7850 12223 7853
rect 14457 7850 14523 7853
rect 7300 7848 7392 7850
rect 7342 7792 7392 7848
rect 7300 7790 7392 7792
rect 12157 7848 14523 7850
rect 12157 7792 12162 7848
rect 12218 7792 14462 7848
rect 14518 7792 14523 7848
rect 12157 7790 14523 7792
rect 7300 7788 7347 7790
rect 7281 7787 7347 7788
rect 12157 7787 12223 7790
rect 14457 7787 14523 7790
rect 4909 7648 5229 7649
rect 4909 7584 4917 7648
rect 4981 7584 4997 7648
rect 5061 7584 5077 7648
rect 5141 7584 5157 7648
rect 5221 7584 5229 7648
rect 4909 7583 5229 7584
rect 12840 7648 13160 7649
rect 12840 7584 12848 7648
rect 12912 7584 12928 7648
rect 12992 7584 13008 7648
rect 13072 7584 13088 7648
rect 13152 7584 13160 7648
rect 12840 7583 13160 7584
rect 20770 7648 21090 7649
rect 20770 7584 20778 7648
rect 20842 7584 20858 7648
rect 20922 7584 20938 7648
rect 21002 7584 21018 7648
rect 21082 7584 21090 7648
rect 20770 7583 21090 7584
rect 8874 7104 9194 7105
rect 8874 7040 8882 7104
rect 8946 7040 8962 7104
rect 9026 7040 9042 7104
rect 9106 7040 9122 7104
rect 9186 7040 9194 7104
rect 8874 7039 9194 7040
rect 16805 7104 17125 7105
rect 16805 7040 16813 7104
rect 16877 7040 16893 7104
rect 16957 7040 16973 7104
rect 17037 7040 17053 7104
rect 17117 7040 17125 7104
rect 16805 7039 17125 7040
rect 4909 6560 5229 6561
rect 4909 6496 4917 6560
rect 4981 6496 4997 6560
rect 5061 6496 5077 6560
rect 5141 6496 5157 6560
rect 5221 6496 5229 6560
rect 4909 6495 5229 6496
rect 12840 6560 13160 6561
rect 12840 6496 12848 6560
rect 12912 6496 12928 6560
rect 12992 6496 13008 6560
rect 13072 6496 13088 6560
rect 13152 6496 13160 6560
rect 12840 6495 13160 6496
rect 20770 6560 21090 6561
rect 20770 6496 20778 6560
rect 20842 6496 20858 6560
rect 20922 6496 20938 6560
rect 21002 6496 21018 6560
rect 21082 6496 21090 6560
rect 20770 6495 21090 6496
rect 8874 6016 9194 6017
rect 8874 5952 8882 6016
rect 8946 5952 8962 6016
rect 9026 5952 9042 6016
rect 9106 5952 9122 6016
rect 9186 5952 9194 6016
rect 8874 5951 9194 5952
rect 16805 6016 17125 6017
rect 16805 5952 16813 6016
rect 16877 5952 16893 6016
rect 16957 5952 16973 6016
rect 17037 5952 17053 6016
rect 17117 5952 17125 6016
rect 16805 5951 17125 5952
rect 4909 5472 5229 5473
rect 4909 5408 4917 5472
rect 4981 5408 4997 5472
rect 5061 5408 5077 5472
rect 5141 5408 5157 5472
rect 5221 5408 5229 5472
rect 4909 5407 5229 5408
rect 12840 5472 13160 5473
rect 12840 5408 12848 5472
rect 12912 5408 12928 5472
rect 12992 5408 13008 5472
rect 13072 5408 13088 5472
rect 13152 5408 13160 5472
rect 12840 5407 13160 5408
rect 20770 5472 21090 5473
rect 20770 5408 20778 5472
rect 20842 5408 20858 5472
rect 20922 5408 20938 5472
rect 21002 5408 21018 5472
rect 21082 5408 21090 5472
rect 20770 5407 21090 5408
rect 2957 4994 3023 4997
rect 6821 4994 6887 4997
rect 2957 4992 6887 4994
rect 2957 4936 2962 4992
rect 3018 4936 6826 4992
rect 6882 4936 6887 4992
rect 2957 4934 6887 4936
rect 2957 4931 3023 4934
rect 6821 4931 6887 4934
rect 8874 4928 9194 4929
rect 8874 4864 8882 4928
rect 8946 4864 8962 4928
rect 9026 4864 9042 4928
rect 9106 4864 9122 4928
rect 9186 4864 9194 4928
rect 8874 4863 9194 4864
rect 16805 4928 17125 4929
rect 16805 4864 16813 4928
rect 16877 4864 16893 4928
rect 16957 4864 16973 4928
rect 17037 4864 17053 4928
rect 17117 4864 17125 4928
rect 16805 4863 17125 4864
rect 12157 4452 12223 4453
rect 12157 4450 12204 4452
rect 12112 4448 12204 4450
rect 12112 4392 12162 4448
rect 12112 4390 12204 4392
rect 12157 4388 12204 4390
rect 12268 4388 12274 4452
rect 12157 4387 12223 4388
rect 4909 4384 5229 4385
rect 4909 4320 4917 4384
rect 4981 4320 4997 4384
rect 5061 4320 5077 4384
rect 5141 4320 5157 4384
rect 5221 4320 5229 4384
rect 4909 4319 5229 4320
rect 12840 4384 13160 4385
rect 12840 4320 12848 4384
rect 12912 4320 12928 4384
rect 12992 4320 13008 4384
rect 13072 4320 13088 4384
rect 13152 4320 13160 4384
rect 12840 4319 13160 4320
rect 20770 4384 21090 4385
rect 20770 4320 20778 4384
rect 20842 4320 20858 4384
rect 20922 4320 20938 4384
rect 21002 4320 21018 4384
rect 21082 4320 21090 4384
rect 20770 4319 21090 4320
rect 13486 4116 13492 4180
rect 13556 4178 13562 4180
rect 13629 4178 13695 4181
rect 13556 4176 13695 4178
rect 13556 4120 13634 4176
rect 13690 4120 13695 4176
rect 13556 4118 13695 4120
rect 13556 4116 13562 4118
rect 13629 4115 13695 4118
rect 8874 3840 9194 3841
rect 8874 3776 8882 3840
rect 8946 3776 8962 3840
rect 9026 3776 9042 3840
rect 9106 3776 9122 3840
rect 9186 3776 9194 3840
rect 8874 3775 9194 3776
rect 16805 3840 17125 3841
rect 16805 3776 16813 3840
rect 16877 3776 16893 3840
rect 16957 3776 16973 3840
rect 17037 3776 17053 3840
rect 17117 3776 17125 3840
rect 16805 3775 17125 3776
rect 4909 3296 5229 3297
rect 4909 3232 4917 3296
rect 4981 3232 4997 3296
rect 5061 3232 5077 3296
rect 5141 3232 5157 3296
rect 5221 3232 5229 3296
rect 4909 3231 5229 3232
rect 12840 3296 13160 3297
rect 12840 3232 12848 3296
rect 12912 3232 12928 3296
rect 12992 3232 13008 3296
rect 13072 3232 13088 3296
rect 13152 3232 13160 3296
rect 12840 3231 13160 3232
rect 20770 3296 21090 3297
rect 20770 3232 20778 3296
rect 20842 3232 20858 3296
rect 20922 3232 20938 3296
rect 21002 3232 21018 3296
rect 21082 3232 21090 3296
rect 20770 3231 21090 3232
rect 9305 3226 9371 3229
rect 9438 3226 9444 3228
rect 9305 3224 9444 3226
rect 9305 3168 9310 3224
rect 9366 3168 9444 3224
rect 9305 3166 9444 3168
rect 9305 3163 9371 3166
rect 9438 3164 9444 3166
rect 9508 3164 9514 3228
rect 0 2818 800 2848
rect 2405 2818 2471 2821
rect 0 2816 2471 2818
rect 0 2760 2410 2816
rect 2466 2760 2471 2816
rect 0 2758 2471 2760
rect 0 2728 800 2758
rect 2405 2755 2471 2758
rect 8874 2752 9194 2753
rect 8874 2688 8882 2752
rect 8946 2688 8962 2752
rect 9026 2688 9042 2752
rect 9106 2688 9122 2752
rect 9186 2688 9194 2752
rect 8874 2687 9194 2688
rect 16805 2752 17125 2753
rect 16805 2688 16813 2752
rect 16877 2688 16893 2752
rect 16957 2688 16973 2752
rect 17037 2688 17053 2752
rect 17117 2688 17125 2752
rect 16805 2687 17125 2688
rect 4909 2208 5229 2209
rect 4909 2144 4917 2208
rect 4981 2144 4997 2208
rect 5061 2144 5077 2208
rect 5141 2144 5157 2208
rect 5221 2144 5229 2208
rect 4909 2143 5229 2144
rect 12840 2208 13160 2209
rect 12840 2144 12848 2208
rect 12912 2144 12928 2208
rect 12992 2144 13008 2208
rect 13072 2144 13088 2208
rect 13152 2144 13160 2208
rect 12840 2143 13160 2144
rect 20770 2208 21090 2209
rect 20770 2144 20778 2208
rect 20842 2144 20858 2208
rect 20922 2144 20938 2208
rect 21002 2144 21018 2208
rect 21082 2144 21090 2208
rect 20770 2143 21090 2144
rect 5441 1868 5507 1869
rect 5390 1804 5396 1868
rect 5460 1866 5507 1868
rect 5460 1864 5552 1866
rect 5502 1808 5552 1864
rect 5460 1806 5552 1808
rect 5460 1804 5507 1806
rect 5441 1803 5507 1804
<< via3 >>
rect 8882 47356 8946 47360
rect 8882 47300 8886 47356
rect 8886 47300 8942 47356
rect 8942 47300 8946 47356
rect 8882 47296 8946 47300
rect 8962 47356 9026 47360
rect 8962 47300 8966 47356
rect 8966 47300 9022 47356
rect 9022 47300 9026 47356
rect 8962 47296 9026 47300
rect 9042 47356 9106 47360
rect 9042 47300 9046 47356
rect 9046 47300 9102 47356
rect 9102 47300 9106 47356
rect 9042 47296 9106 47300
rect 9122 47356 9186 47360
rect 9122 47300 9126 47356
rect 9126 47300 9182 47356
rect 9182 47300 9186 47356
rect 9122 47296 9186 47300
rect 16813 47356 16877 47360
rect 16813 47300 16817 47356
rect 16817 47300 16873 47356
rect 16873 47300 16877 47356
rect 16813 47296 16877 47300
rect 16893 47356 16957 47360
rect 16893 47300 16897 47356
rect 16897 47300 16953 47356
rect 16953 47300 16957 47356
rect 16893 47296 16957 47300
rect 16973 47356 17037 47360
rect 16973 47300 16977 47356
rect 16977 47300 17033 47356
rect 17033 47300 17037 47356
rect 16973 47296 17037 47300
rect 17053 47356 17117 47360
rect 17053 47300 17057 47356
rect 17057 47300 17113 47356
rect 17113 47300 17117 47356
rect 17053 47296 17117 47300
rect 4917 46812 4981 46816
rect 4917 46756 4921 46812
rect 4921 46756 4977 46812
rect 4977 46756 4981 46812
rect 4917 46752 4981 46756
rect 4997 46812 5061 46816
rect 4997 46756 5001 46812
rect 5001 46756 5057 46812
rect 5057 46756 5061 46812
rect 4997 46752 5061 46756
rect 5077 46812 5141 46816
rect 5077 46756 5081 46812
rect 5081 46756 5137 46812
rect 5137 46756 5141 46812
rect 5077 46752 5141 46756
rect 5157 46812 5221 46816
rect 5157 46756 5161 46812
rect 5161 46756 5217 46812
rect 5217 46756 5221 46812
rect 5157 46752 5221 46756
rect 12848 46812 12912 46816
rect 12848 46756 12852 46812
rect 12852 46756 12908 46812
rect 12908 46756 12912 46812
rect 12848 46752 12912 46756
rect 12928 46812 12992 46816
rect 12928 46756 12932 46812
rect 12932 46756 12988 46812
rect 12988 46756 12992 46812
rect 12928 46752 12992 46756
rect 13008 46812 13072 46816
rect 13008 46756 13012 46812
rect 13012 46756 13068 46812
rect 13068 46756 13072 46812
rect 13008 46752 13072 46756
rect 13088 46812 13152 46816
rect 13088 46756 13092 46812
rect 13092 46756 13148 46812
rect 13148 46756 13152 46812
rect 13088 46752 13152 46756
rect 20778 46812 20842 46816
rect 20778 46756 20782 46812
rect 20782 46756 20838 46812
rect 20838 46756 20842 46812
rect 20778 46752 20842 46756
rect 20858 46812 20922 46816
rect 20858 46756 20862 46812
rect 20862 46756 20918 46812
rect 20918 46756 20922 46812
rect 20858 46752 20922 46756
rect 20938 46812 21002 46816
rect 20938 46756 20942 46812
rect 20942 46756 20998 46812
rect 20998 46756 21002 46812
rect 20938 46752 21002 46756
rect 21018 46812 21082 46816
rect 21018 46756 21022 46812
rect 21022 46756 21078 46812
rect 21078 46756 21082 46812
rect 21018 46752 21082 46756
rect 8882 46268 8946 46272
rect 8882 46212 8886 46268
rect 8886 46212 8942 46268
rect 8942 46212 8946 46268
rect 8882 46208 8946 46212
rect 8962 46268 9026 46272
rect 8962 46212 8966 46268
rect 8966 46212 9022 46268
rect 9022 46212 9026 46268
rect 8962 46208 9026 46212
rect 9042 46268 9106 46272
rect 9042 46212 9046 46268
rect 9046 46212 9102 46268
rect 9102 46212 9106 46268
rect 9042 46208 9106 46212
rect 9122 46268 9186 46272
rect 9122 46212 9126 46268
rect 9126 46212 9182 46268
rect 9182 46212 9186 46268
rect 9122 46208 9186 46212
rect 16813 46268 16877 46272
rect 16813 46212 16817 46268
rect 16817 46212 16873 46268
rect 16873 46212 16877 46268
rect 16813 46208 16877 46212
rect 16893 46268 16957 46272
rect 16893 46212 16897 46268
rect 16897 46212 16953 46268
rect 16953 46212 16957 46268
rect 16893 46208 16957 46212
rect 16973 46268 17037 46272
rect 16973 46212 16977 46268
rect 16977 46212 17033 46268
rect 17033 46212 17037 46268
rect 16973 46208 17037 46212
rect 17053 46268 17117 46272
rect 17053 46212 17057 46268
rect 17057 46212 17113 46268
rect 17113 46212 17117 46268
rect 17053 46208 17117 46212
rect 4917 45724 4981 45728
rect 4917 45668 4921 45724
rect 4921 45668 4977 45724
rect 4977 45668 4981 45724
rect 4917 45664 4981 45668
rect 4997 45724 5061 45728
rect 4997 45668 5001 45724
rect 5001 45668 5057 45724
rect 5057 45668 5061 45724
rect 4997 45664 5061 45668
rect 5077 45724 5141 45728
rect 5077 45668 5081 45724
rect 5081 45668 5137 45724
rect 5137 45668 5141 45724
rect 5077 45664 5141 45668
rect 5157 45724 5221 45728
rect 5157 45668 5161 45724
rect 5161 45668 5217 45724
rect 5217 45668 5221 45724
rect 5157 45664 5221 45668
rect 12848 45724 12912 45728
rect 12848 45668 12852 45724
rect 12852 45668 12908 45724
rect 12908 45668 12912 45724
rect 12848 45664 12912 45668
rect 12928 45724 12992 45728
rect 12928 45668 12932 45724
rect 12932 45668 12988 45724
rect 12988 45668 12992 45724
rect 12928 45664 12992 45668
rect 13008 45724 13072 45728
rect 13008 45668 13012 45724
rect 13012 45668 13068 45724
rect 13068 45668 13072 45724
rect 13008 45664 13072 45668
rect 13088 45724 13152 45728
rect 13088 45668 13092 45724
rect 13092 45668 13148 45724
rect 13148 45668 13152 45724
rect 13088 45664 13152 45668
rect 20778 45724 20842 45728
rect 20778 45668 20782 45724
rect 20782 45668 20838 45724
rect 20838 45668 20842 45724
rect 20778 45664 20842 45668
rect 20858 45724 20922 45728
rect 20858 45668 20862 45724
rect 20862 45668 20918 45724
rect 20918 45668 20922 45724
rect 20858 45664 20922 45668
rect 20938 45724 21002 45728
rect 20938 45668 20942 45724
rect 20942 45668 20998 45724
rect 20998 45668 21002 45724
rect 20938 45664 21002 45668
rect 21018 45724 21082 45728
rect 21018 45668 21022 45724
rect 21022 45668 21078 45724
rect 21078 45668 21082 45724
rect 21018 45664 21082 45668
rect 8882 45180 8946 45184
rect 8882 45124 8886 45180
rect 8886 45124 8942 45180
rect 8942 45124 8946 45180
rect 8882 45120 8946 45124
rect 8962 45180 9026 45184
rect 8962 45124 8966 45180
rect 8966 45124 9022 45180
rect 9022 45124 9026 45180
rect 8962 45120 9026 45124
rect 9042 45180 9106 45184
rect 9042 45124 9046 45180
rect 9046 45124 9102 45180
rect 9102 45124 9106 45180
rect 9042 45120 9106 45124
rect 9122 45180 9186 45184
rect 9122 45124 9126 45180
rect 9126 45124 9182 45180
rect 9182 45124 9186 45180
rect 9122 45120 9186 45124
rect 16813 45180 16877 45184
rect 16813 45124 16817 45180
rect 16817 45124 16873 45180
rect 16873 45124 16877 45180
rect 16813 45120 16877 45124
rect 16893 45180 16957 45184
rect 16893 45124 16897 45180
rect 16897 45124 16953 45180
rect 16953 45124 16957 45180
rect 16893 45120 16957 45124
rect 16973 45180 17037 45184
rect 16973 45124 16977 45180
rect 16977 45124 17033 45180
rect 17033 45124 17037 45180
rect 16973 45120 17037 45124
rect 17053 45180 17117 45184
rect 17053 45124 17057 45180
rect 17057 45124 17113 45180
rect 17113 45124 17117 45180
rect 17053 45120 17117 45124
rect 4917 44636 4981 44640
rect 4917 44580 4921 44636
rect 4921 44580 4977 44636
rect 4977 44580 4981 44636
rect 4917 44576 4981 44580
rect 4997 44636 5061 44640
rect 4997 44580 5001 44636
rect 5001 44580 5057 44636
rect 5057 44580 5061 44636
rect 4997 44576 5061 44580
rect 5077 44636 5141 44640
rect 5077 44580 5081 44636
rect 5081 44580 5137 44636
rect 5137 44580 5141 44636
rect 5077 44576 5141 44580
rect 5157 44636 5221 44640
rect 5157 44580 5161 44636
rect 5161 44580 5217 44636
rect 5217 44580 5221 44636
rect 5157 44576 5221 44580
rect 12848 44636 12912 44640
rect 12848 44580 12852 44636
rect 12852 44580 12908 44636
rect 12908 44580 12912 44636
rect 12848 44576 12912 44580
rect 12928 44636 12992 44640
rect 12928 44580 12932 44636
rect 12932 44580 12988 44636
rect 12988 44580 12992 44636
rect 12928 44576 12992 44580
rect 13008 44636 13072 44640
rect 13008 44580 13012 44636
rect 13012 44580 13068 44636
rect 13068 44580 13072 44636
rect 13008 44576 13072 44580
rect 13088 44636 13152 44640
rect 13088 44580 13092 44636
rect 13092 44580 13148 44636
rect 13148 44580 13152 44636
rect 13088 44576 13152 44580
rect 20778 44636 20842 44640
rect 20778 44580 20782 44636
rect 20782 44580 20838 44636
rect 20838 44580 20842 44636
rect 20778 44576 20842 44580
rect 20858 44636 20922 44640
rect 20858 44580 20862 44636
rect 20862 44580 20918 44636
rect 20918 44580 20922 44636
rect 20858 44576 20922 44580
rect 20938 44636 21002 44640
rect 20938 44580 20942 44636
rect 20942 44580 20998 44636
rect 20998 44580 21002 44636
rect 20938 44576 21002 44580
rect 21018 44636 21082 44640
rect 21018 44580 21022 44636
rect 21022 44580 21078 44636
rect 21078 44580 21082 44636
rect 21018 44576 21082 44580
rect 8882 44092 8946 44096
rect 8882 44036 8886 44092
rect 8886 44036 8942 44092
rect 8942 44036 8946 44092
rect 8882 44032 8946 44036
rect 8962 44092 9026 44096
rect 8962 44036 8966 44092
rect 8966 44036 9022 44092
rect 9022 44036 9026 44092
rect 8962 44032 9026 44036
rect 9042 44092 9106 44096
rect 9042 44036 9046 44092
rect 9046 44036 9102 44092
rect 9102 44036 9106 44092
rect 9042 44032 9106 44036
rect 9122 44092 9186 44096
rect 9122 44036 9126 44092
rect 9126 44036 9182 44092
rect 9182 44036 9186 44092
rect 9122 44032 9186 44036
rect 16813 44092 16877 44096
rect 16813 44036 16817 44092
rect 16817 44036 16873 44092
rect 16873 44036 16877 44092
rect 16813 44032 16877 44036
rect 16893 44092 16957 44096
rect 16893 44036 16897 44092
rect 16897 44036 16953 44092
rect 16953 44036 16957 44092
rect 16893 44032 16957 44036
rect 16973 44092 17037 44096
rect 16973 44036 16977 44092
rect 16977 44036 17033 44092
rect 17033 44036 17037 44092
rect 16973 44032 17037 44036
rect 17053 44092 17117 44096
rect 17053 44036 17057 44092
rect 17057 44036 17113 44092
rect 17113 44036 17117 44092
rect 17053 44032 17117 44036
rect 4917 43548 4981 43552
rect 4917 43492 4921 43548
rect 4921 43492 4977 43548
rect 4977 43492 4981 43548
rect 4917 43488 4981 43492
rect 4997 43548 5061 43552
rect 4997 43492 5001 43548
rect 5001 43492 5057 43548
rect 5057 43492 5061 43548
rect 4997 43488 5061 43492
rect 5077 43548 5141 43552
rect 5077 43492 5081 43548
rect 5081 43492 5137 43548
rect 5137 43492 5141 43548
rect 5077 43488 5141 43492
rect 5157 43548 5221 43552
rect 5157 43492 5161 43548
rect 5161 43492 5217 43548
rect 5217 43492 5221 43548
rect 5157 43488 5221 43492
rect 12848 43548 12912 43552
rect 12848 43492 12852 43548
rect 12852 43492 12908 43548
rect 12908 43492 12912 43548
rect 12848 43488 12912 43492
rect 12928 43548 12992 43552
rect 12928 43492 12932 43548
rect 12932 43492 12988 43548
rect 12988 43492 12992 43548
rect 12928 43488 12992 43492
rect 13008 43548 13072 43552
rect 13008 43492 13012 43548
rect 13012 43492 13068 43548
rect 13068 43492 13072 43548
rect 13008 43488 13072 43492
rect 13088 43548 13152 43552
rect 13088 43492 13092 43548
rect 13092 43492 13148 43548
rect 13148 43492 13152 43548
rect 13088 43488 13152 43492
rect 20778 43548 20842 43552
rect 20778 43492 20782 43548
rect 20782 43492 20838 43548
rect 20838 43492 20842 43548
rect 20778 43488 20842 43492
rect 20858 43548 20922 43552
rect 20858 43492 20862 43548
rect 20862 43492 20918 43548
rect 20918 43492 20922 43548
rect 20858 43488 20922 43492
rect 20938 43548 21002 43552
rect 20938 43492 20942 43548
rect 20942 43492 20998 43548
rect 20998 43492 21002 43548
rect 20938 43488 21002 43492
rect 21018 43548 21082 43552
rect 21018 43492 21022 43548
rect 21022 43492 21078 43548
rect 21078 43492 21082 43548
rect 21018 43488 21082 43492
rect 8882 43004 8946 43008
rect 8882 42948 8886 43004
rect 8886 42948 8942 43004
rect 8942 42948 8946 43004
rect 8882 42944 8946 42948
rect 8962 43004 9026 43008
rect 8962 42948 8966 43004
rect 8966 42948 9022 43004
rect 9022 42948 9026 43004
rect 8962 42944 9026 42948
rect 9042 43004 9106 43008
rect 9042 42948 9046 43004
rect 9046 42948 9102 43004
rect 9102 42948 9106 43004
rect 9042 42944 9106 42948
rect 9122 43004 9186 43008
rect 9122 42948 9126 43004
rect 9126 42948 9182 43004
rect 9182 42948 9186 43004
rect 9122 42944 9186 42948
rect 16813 43004 16877 43008
rect 16813 42948 16817 43004
rect 16817 42948 16873 43004
rect 16873 42948 16877 43004
rect 16813 42944 16877 42948
rect 16893 43004 16957 43008
rect 16893 42948 16897 43004
rect 16897 42948 16953 43004
rect 16953 42948 16957 43004
rect 16893 42944 16957 42948
rect 16973 43004 17037 43008
rect 16973 42948 16977 43004
rect 16977 42948 17033 43004
rect 17033 42948 17037 43004
rect 16973 42944 17037 42948
rect 17053 43004 17117 43008
rect 17053 42948 17057 43004
rect 17057 42948 17113 43004
rect 17113 42948 17117 43004
rect 17053 42944 17117 42948
rect 4917 42460 4981 42464
rect 4917 42404 4921 42460
rect 4921 42404 4977 42460
rect 4977 42404 4981 42460
rect 4917 42400 4981 42404
rect 4997 42460 5061 42464
rect 4997 42404 5001 42460
rect 5001 42404 5057 42460
rect 5057 42404 5061 42460
rect 4997 42400 5061 42404
rect 5077 42460 5141 42464
rect 5077 42404 5081 42460
rect 5081 42404 5137 42460
rect 5137 42404 5141 42460
rect 5077 42400 5141 42404
rect 5157 42460 5221 42464
rect 5157 42404 5161 42460
rect 5161 42404 5217 42460
rect 5217 42404 5221 42460
rect 5157 42400 5221 42404
rect 12848 42460 12912 42464
rect 12848 42404 12852 42460
rect 12852 42404 12908 42460
rect 12908 42404 12912 42460
rect 12848 42400 12912 42404
rect 12928 42460 12992 42464
rect 12928 42404 12932 42460
rect 12932 42404 12988 42460
rect 12988 42404 12992 42460
rect 12928 42400 12992 42404
rect 13008 42460 13072 42464
rect 13008 42404 13012 42460
rect 13012 42404 13068 42460
rect 13068 42404 13072 42460
rect 13008 42400 13072 42404
rect 13088 42460 13152 42464
rect 13088 42404 13092 42460
rect 13092 42404 13148 42460
rect 13148 42404 13152 42460
rect 13088 42400 13152 42404
rect 20778 42460 20842 42464
rect 20778 42404 20782 42460
rect 20782 42404 20838 42460
rect 20838 42404 20842 42460
rect 20778 42400 20842 42404
rect 20858 42460 20922 42464
rect 20858 42404 20862 42460
rect 20862 42404 20918 42460
rect 20918 42404 20922 42460
rect 20858 42400 20922 42404
rect 20938 42460 21002 42464
rect 20938 42404 20942 42460
rect 20942 42404 20998 42460
rect 20998 42404 21002 42460
rect 20938 42400 21002 42404
rect 21018 42460 21082 42464
rect 21018 42404 21022 42460
rect 21022 42404 21078 42460
rect 21078 42404 21082 42460
rect 21018 42400 21082 42404
rect 8882 41916 8946 41920
rect 8882 41860 8886 41916
rect 8886 41860 8942 41916
rect 8942 41860 8946 41916
rect 8882 41856 8946 41860
rect 8962 41916 9026 41920
rect 8962 41860 8966 41916
rect 8966 41860 9022 41916
rect 9022 41860 9026 41916
rect 8962 41856 9026 41860
rect 9042 41916 9106 41920
rect 9042 41860 9046 41916
rect 9046 41860 9102 41916
rect 9102 41860 9106 41916
rect 9042 41856 9106 41860
rect 9122 41916 9186 41920
rect 9122 41860 9126 41916
rect 9126 41860 9182 41916
rect 9182 41860 9186 41916
rect 9122 41856 9186 41860
rect 16813 41916 16877 41920
rect 16813 41860 16817 41916
rect 16817 41860 16873 41916
rect 16873 41860 16877 41916
rect 16813 41856 16877 41860
rect 16893 41916 16957 41920
rect 16893 41860 16897 41916
rect 16897 41860 16953 41916
rect 16953 41860 16957 41916
rect 16893 41856 16957 41860
rect 16973 41916 17037 41920
rect 16973 41860 16977 41916
rect 16977 41860 17033 41916
rect 17033 41860 17037 41916
rect 16973 41856 17037 41860
rect 17053 41916 17117 41920
rect 17053 41860 17057 41916
rect 17057 41860 17113 41916
rect 17113 41860 17117 41916
rect 17053 41856 17117 41860
rect 4917 41372 4981 41376
rect 4917 41316 4921 41372
rect 4921 41316 4977 41372
rect 4977 41316 4981 41372
rect 4917 41312 4981 41316
rect 4997 41372 5061 41376
rect 4997 41316 5001 41372
rect 5001 41316 5057 41372
rect 5057 41316 5061 41372
rect 4997 41312 5061 41316
rect 5077 41372 5141 41376
rect 5077 41316 5081 41372
rect 5081 41316 5137 41372
rect 5137 41316 5141 41372
rect 5077 41312 5141 41316
rect 5157 41372 5221 41376
rect 5157 41316 5161 41372
rect 5161 41316 5217 41372
rect 5217 41316 5221 41372
rect 5157 41312 5221 41316
rect 12848 41372 12912 41376
rect 12848 41316 12852 41372
rect 12852 41316 12908 41372
rect 12908 41316 12912 41372
rect 12848 41312 12912 41316
rect 12928 41372 12992 41376
rect 12928 41316 12932 41372
rect 12932 41316 12988 41372
rect 12988 41316 12992 41372
rect 12928 41312 12992 41316
rect 13008 41372 13072 41376
rect 13008 41316 13012 41372
rect 13012 41316 13068 41372
rect 13068 41316 13072 41372
rect 13008 41312 13072 41316
rect 13088 41372 13152 41376
rect 13088 41316 13092 41372
rect 13092 41316 13148 41372
rect 13148 41316 13152 41372
rect 13088 41312 13152 41316
rect 20778 41372 20842 41376
rect 20778 41316 20782 41372
rect 20782 41316 20838 41372
rect 20838 41316 20842 41372
rect 20778 41312 20842 41316
rect 20858 41372 20922 41376
rect 20858 41316 20862 41372
rect 20862 41316 20918 41372
rect 20918 41316 20922 41372
rect 20858 41312 20922 41316
rect 20938 41372 21002 41376
rect 20938 41316 20942 41372
rect 20942 41316 20998 41372
rect 20998 41316 21002 41372
rect 20938 41312 21002 41316
rect 21018 41372 21082 41376
rect 21018 41316 21022 41372
rect 21022 41316 21078 41372
rect 21078 41316 21082 41372
rect 21018 41312 21082 41316
rect 8882 40828 8946 40832
rect 8882 40772 8886 40828
rect 8886 40772 8942 40828
rect 8942 40772 8946 40828
rect 8882 40768 8946 40772
rect 8962 40828 9026 40832
rect 8962 40772 8966 40828
rect 8966 40772 9022 40828
rect 9022 40772 9026 40828
rect 8962 40768 9026 40772
rect 9042 40828 9106 40832
rect 9042 40772 9046 40828
rect 9046 40772 9102 40828
rect 9102 40772 9106 40828
rect 9042 40768 9106 40772
rect 9122 40828 9186 40832
rect 9122 40772 9126 40828
rect 9126 40772 9182 40828
rect 9182 40772 9186 40828
rect 9122 40768 9186 40772
rect 16813 40828 16877 40832
rect 16813 40772 16817 40828
rect 16817 40772 16873 40828
rect 16873 40772 16877 40828
rect 16813 40768 16877 40772
rect 16893 40828 16957 40832
rect 16893 40772 16897 40828
rect 16897 40772 16953 40828
rect 16953 40772 16957 40828
rect 16893 40768 16957 40772
rect 16973 40828 17037 40832
rect 16973 40772 16977 40828
rect 16977 40772 17033 40828
rect 17033 40772 17037 40828
rect 16973 40768 17037 40772
rect 17053 40828 17117 40832
rect 17053 40772 17057 40828
rect 17057 40772 17113 40828
rect 17113 40772 17117 40828
rect 17053 40768 17117 40772
rect 4917 40284 4981 40288
rect 4917 40228 4921 40284
rect 4921 40228 4977 40284
rect 4977 40228 4981 40284
rect 4917 40224 4981 40228
rect 4997 40284 5061 40288
rect 4997 40228 5001 40284
rect 5001 40228 5057 40284
rect 5057 40228 5061 40284
rect 4997 40224 5061 40228
rect 5077 40284 5141 40288
rect 5077 40228 5081 40284
rect 5081 40228 5137 40284
rect 5137 40228 5141 40284
rect 5077 40224 5141 40228
rect 5157 40284 5221 40288
rect 5157 40228 5161 40284
rect 5161 40228 5217 40284
rect 5217 40228 5221 40284
rect 5157 40224 5221 40228
rect 12848 40284 12912 40288
rect 12848 40228 12852 40284
rect 12852 40228 12908 40284
rect 12908 40228 12912 40284
rect 12848 40224 12912 40228
rect 12928 40284 12992 40288
rect 12928 40228 12932 40284
rect 12932 40228 12988 40284
rect 12988 40228 12992 40284
rect 12928 40224 12992 40228
rect 13008 40284 13072 40288
rect 13008 40228 13012 40284
rect 13012 40228 13068 40284
rect 13068 40228 13072 40284
rect 13008 40224 13072 40228
rect 13088 40284 13152 40288
rect 13088 40228 13092 40284
rect 13092 40228 13148 40284
rect 13148 40228 13152 40284
rect 13088 40224 13152 40228
rect 20778 40284 20842 40288
rect 20778 40228 20782 40284
rect 20782 40228 20838 40284
rect 20838 40228 20842 40284
rect 20778 40224 20842 40228
rect 20858 40284 20922 40288
rect 20858 40228 20862 40284
rect 20862 40228 20918 40284
rect 20918 40228 20922 40284
rect 20858 40224 20922 40228
rect 20938 40284 21002 40288
rect 20938 40228 20942 40284
rect 20942 40228 20998 40284
rect 20998 40228 21002 40284
rect 20938 40224 21002 40228
rect 21018 40284 21082 40288
rect 21018 40228 21022 40284
rect 21022 40228 21078 40284
rect 21078 40228 21082 40284
rect 21018 40224 21082 40228
rect 8882 39740 8946 39744
rect 8882 39684 8886 39740
rect 8886 39684 8942 39740
rect 8942 39684 8946 39740
rect 8882 39680 8946 39684
rect 8962 39740 9026 39744
rect 8962 39684 8966 39740
rect 8966 39684 9022 39740
rect 9022 39684 9026 39740
rect 8962 39680 9026 39684
rect 9042 39740 9106 39744
rect 9042 39684 9046 39740
rect 9046 39684 9102 39740
rect 9102 39684 9106 39740
rect 9042 39680 9106 39684
rect 9122 39740 9186 39744
rect 9122 39684 9126 39740
rect 9126 39684 9182 39740
rect 9182 39684 9186 39740
rect 9122 39680 9186 39684
rect 16813 39740 16877 39744
rect 16813 39684 16817 39740
rect 16817 39684 16873 39740
rect 16873 39684 16877 39740
rect 16813 39680 16877 39684
rect 16893 39740 16957 39744
rect 16893 39684 16897 39740
rect 16897 39684 16953 39740
rect 16953 39684 16957 39740
rect 16893 39680 16957 39684
rect 16973 39740 17037 39744
rect 16973 39684 16977 39740
rect 16977 39684 17033 39740
rect 17033 39684 17037 39740
rect 16973 39680 17037 39684
rect 17053 39740 17117 39744
rect 17053 39684 17057 39740
rect 17057 39684 17113 39740
rect 17113 39684 17117 39740
rect 17053 39680 17117 39684
rect 4917 39196 4981 39200
rect 4917 39140 4921 39196
rect 4921 39140 4977 39196
rect 4977 39140 4981 39196
rect 4917 39136 4981 39140
rect 4997 39196 5061 39200
rect 4997 39140 5001 39196
rect 5001 39140 5057 39196
rect 5057 39140 5061 39196
rect 4997 39136 5061 39140
rect 5077 39196 5141 39200
rect 5077 39140 5081 39196
rect 5081 39140 5137 39196
rect 5137 39140 5141 39196
rect 5077 39136 5141 39140
rect 5157 39196 5221 39200
rect 5157 39140 5161 39196
rect 5161 39140 5217 39196
rect 5217 39140 5221 39196
rect 5157 39136 5221 39140
rect 12848 39196 12912 39200
rect 12848 39140 12852 39196
rect 12852 39140 12908 39196
rect 12908 39140 12912 39196
rect 12848 39136 12912 39140
rect 12928 39196 12992 39200
rect 12928 39140 12932 39196
rect 12932 39140 12988 39196
rect 12988 39140 12992 39196
rect 12928 39136 12992 39140
rect 13008 39196 13072 39200
rect 13008 39140 13012 39196
rect 13012 39140 13068 39196
rect 13068 39140 13072 39196
rect 13008 39136 13072 39140
rect 13088 39196 13152 39200
rect 13088 39140 13092 39196
rect 13092 39140 13148 39196
rect 13148 39140 13152 39196
rect 13088 39136 13152 39140
rect 20778 39196 20842 39200
rect 20778 39140 20782 39196
rect 20782 39140 20838 39196
rect 20838 39140 20842 39196
rect 20778 39136 20842 39140
rect 20858 39196 20922 39200
rect 20858 39140 20862 39196
rect 20862 39140 20918 39196
rect 20918 39140 20922 39196
rect 20858 39136 20922 39140
rect 20938 39196 21002 39200
rect 20938 39140 20942 39196
rect 20942 39140 20998 39196
rect 20998 39140 21002 39196
rect 20938 39136 21002 39140
rect 21018 39196 21082 39200
rect 21018 39140 21022 39196
rect 21022 39140 21078 39196
rect 21078 39140 21082 39196
rect 21018 39136 21082 39140
rect 8882 38652 8946 38656
rect 8882 38596 8886 38652
rect 8886 38596 8942 38652
rect 8942 38596 8946 38652
rect 8882 38592 8946 38596
rect 8962 38652 9026 38656
rect 8962 38596 8966 38652
rect 8966 38596 9022 38652
rect 9022 38596 9026 38652
rect 8962 38592 9026 38596
rect 9042 38652 9106 38656
rect 9042 38596 9046 38652
rect 9046 38596 9102 38652
rect 9102 38596 9106 38652
rect 9042 38592 9106 38596
rect 9122 38652 9186 38656
rect 9122 38596 9126 38652
rect 9126 38596 9182 38652
rect 9182 38596 9186 38652
rect 9122 38592 9186 38596
rect 16813 38652 16877 38656
rect 16813 38596 16817 38652
rect 16817 38596 16873 38652
rect 16873 38596 16877 38652
rect 16813 38592 16877 38596
rect 16893 38652 16957 38656
rect 16893 38596 16897 38652
rect 16897 38596 16953 38652
rect 16953 38596 16957 38652
rect 16893 38592 16957 38596
rect 16973 38652 17037 38656
rect 16973 38596 16977 38652
rect 16977 38596 17033 38652
rect 17033 38596 17037 38652
rect 16973 38592 17037 38596
rect 17053 38652 17117 38656
rect 17053 38596 17057 38652
rect 17057 38596 17113 38652
rect 17113 38596 17117 38652
rect 17053 38592 17117 38596
rect 4917 38108 4981 38112
rect 4917 38052 4921 38108
rect 4921 38052 4977 38108
rect 4977 38052 4981 38108
rect 4917 38048 4981 38052
rect 4997 38108 5061 38112
rect 4997 38052 5001 38108
rect 5001 38052 5057 38108
rect 5057 38052 5061 38108
rect 4997 38048 5061 38052
rect 5077 38108 5141 38112
rect 5077 38052 5081 38108
rect 5081 38052 5137 38108
rect 5137 38052 5141 38108
rect 5077 38048 5141 38052
rect 5157 38108 5221 38112
rect 5157 38052 5161 38108
rect 5161 38052 5217 38108
rect 5217 38052 5221 38108
rect 5157 38048 5221 38052
rect 12848 38108 12912 38112
rect 12848 38052 12852 38108
rect 12852 38052 12908 38108
rect 12908 38052 12912 38108
rect 12848 38048 12912 38052
rect 12928 38108 12992 38112
rect 12928 38052 12932 38108
rect 12932 38052 12988 38108
rect 12988 38052 12992 38108
rect 12928 38048 12992 38052
rect 13008 38108 13072 38112
rect 13008 38052 13012 38108
rect 13012 38052 13068 38108
rect 13068 38052 13072 38108
rect 13008 38048 13072 38052
rect 13088 38108 13152 38112
rect 13088 38052 13092 38108
rect 13092 38052 13148 38108
rect 13148 38052 13152 38108
rect 13088 38048 13152 38052
rect 20778 38108 20842 38112
rect 20778 38052 20782 38108
rect 20782 38052 20838 38108
rect 20838 38052 20842 38108
rect 20778 38048 20842 38052
rect 20858 38108 20922 38112
rect 20858 38052 20862 38108
rect 20862 38052 20918 38108
rect 20918 38052 20922 38108
rect 20858 38048 20922 38052
rect 20938 38108 21002 38112
rect 20938 38052 20942 38108
rect 20942 38052 20998 38108
rect 20998 38052 21002 38108
rect 20938 38048 21002 38052
rect 21018 38108 21082 38112
rect 21018 38052 21022 38108
rect 21022 38052 21078 38108
rect 21078 38052 21082 38108
rect 21018 38048 21082 38052
rect 8882 37564 8946 37568
rect 8882 37508 8886 37564
rect 8886 37508 8942 37564
rect 8942 37508 8946 37564
rect 8882 37504 8946 37508
rect 8962 37564 9026 37568
rect 8962 37508 8966 37564
rect 8966 37508 9022 37564
rect 9022 37508 9026 37564
rect 8962 37504 9026 37508
rect 9042 37564 9106 37568
rect 9042 37508 9046 37564
rect 9046 37508 9102 37564
rect 9102 37508 9106 37564
rect 9042 37504 9106 37508
rect 9122 37564 9186 37568
rect 9122 37508 9126 37564
rect 9126 37508 9182 37564
rect 9182 37508 9186 37564
rect 9122 37504 9186 37508
rect 16813 37564 16877 37568
rect 16813 37508 16817 37564
rect 16817 37508 16873 37564
rect 16873 37508 16877 37564
rect 16813 37504 16877 37508
rect 16893 37564 16957 37568
rect 16893 37508 16897 37564
rect 16897 37508 16953 37564
rect 16953 37508 16957 37564
rect 16893 37504 16957 37508
rect 16973 37564 17037 37568
rect 16973 37508 16977 37564
rect 16977 37508 17033 37564
rect 17033 37508 17037 37564
rect 16973 37504 17037 37508
rect 17053 37564 17117 37568
rect 17053 37508 17057 37564
rect 17057 37508 17113 37564
rect 17113 37508 17117 37564
rect 17053 37504 17117 37508
rect 4917 37020 4981 37024
rect 4917 36964 4921 37020
rect 4921 36964 4977 37020
rect 4977 36964 4981 37020
rect 4917 36960 4981 36964
rect 4997 37020 5061 37024
rect 4997 36964 5001 37020
rect 5001 36964 5057 37020
rect 5057 36964 5061 37020
rect 4997 36960 5061 36964
rect 5077 37020 5141 37024
rect 5077 36964 5081 37020
rect 5081 36964 5137 37020
rect 5137 36964 5141 37020
rect 5077 36960 5141 36964
rect 5157 37020 5221 37024
rect 5157 36964 5161 37020
rect 5161 36964 5217 37020
rect 5217 36964 5221 37020
rect 5157 36960 5221 36964
rect 12848 37020 12912 37024
rect 12848 36964 12852 37020
rect 12852 36964 12908 37020
rect 12908 36964 12912 37020
rect 12848 36960 12912 36964
rect 12928 37020 12992 37024
rect 12928 36964 12932 37020
rect 12932 36964 12988 37020
rect 12988 36964 12992 37020
rect 12928 36960 12992 36964
rect 13008 37020 13072 37024
rect 13008 36964 13012 37020
rect 13012 36964 13068 37020
rect 13068 36964 13072 37020
rect 13008 36960 13072 36964
rect 13088 37020 13152 37024
rect 13088 36964 13092 37020
rect 13092 36964 13148 37020
rect 13148 36964 13152 37020
rect 13088 36960 13152 36964
rect 20778 37020 20842 37024
rect 20778 36964 20782 37020
rect 20782 36964 20838 37020
rect 20838 36964 20842 37020
rect 20778 36960 20842 36964
rect 20858 37020 20922 37024
rect 20858 36964 20862 37020
rect 20862 36964 20918 37020
rect 20918 36964 20922 37020
rect 20858 36960 20922 36964
rect 20938 37020 21002 37024
rect 20938 36964 20942 37020
rect 20942 36964 20998 37020
rect 20998 36964 21002 37020
rect 20938 36960 21002 36964
rect 21018 37020 21082 37024
rect 21018 36964 21022 37020
rect 21022 36964 21078 37020
rect 21078 36964 21082 37020
rect 21018 36960 21082 36964
rect 8882 36476 8946 36480
rect 8882 36420 8886 36476
rect 8886 36420 8942 36476
rect 8942 36420 8946 36476
rect 8882 36416 8946 36420
rect 8962 36476 9026 36480
rect 8962 36420 8966 36476
rect 8966 36420 9022 36476
rect 9022 36420 9026 36476
rect 8962 36416 9026 36420
rect 9042 36476 9106 36480
rect 9042 36420 9046 36476
rect 9046 36420 9102 36476
rect 9102 36420 9106 36476
rect 9042 36416 9106 36420
rect 9122 36476 9186 36480
rect 9122 36420 9126 36476
rect 9126 36420 9182 36476
rect 9182 36420 9186 36476
rect 9122 36416 9186 36420
rect 16813 36476 16877 36480
rect 16813 36420 16817 36476
rect 16817 36420 16873 36476
rect 16873 36420 16877 36476
rect 16813 36416 16877 36420
rect 16893 36476 16957 36480
rect 16893 36420 16897 36476
rect 16897 36420 16953 36476
rect 16953 36420 16957 36476
rect 16893 36416 16957 36420
rect 16973 36476 17037 36480
rect 16973 36420 16977 36476
rect 16977 36420 17033 36476
rect 17033 36420 17037 36476
rect 16973 36416 17037 36420
rect 17053 36476 17117 36480
rect 17053 36420 17057 36476
rect 17057 36420 17113 36476
rect 17113 36420 17117 36476
rect 17053 36416 17117 36420
rect 4917 35932 4981 35936
rect 4917 35876 4921 35932
rect 4921 35876 4977 35932
rect 4977 35876 4981 35932
rect 4917 35872 4981 35876
rect 4997 35932 5061 35936
rect 4997 35876 5001 35932
rect 5001 35876 5057 35932
rect 5057 35876 5061 35932
rect 4997 35872 5061 35876
rect 5077 35932 5141 35936
rect 5077 35876 5081 35932
rect 5081 35876 5137 35932
rect 5137 35876 5141 35932
rect 5077 35872 5141 35876
rect 5157 35932 5221 35936
rect 5157 35876 5161 35932
rect 5161 35876 5217 35932
rect 5217 35876 5221 35932
rect 5157 35872 5221 35876
rect 12848 35932 12912 35936
rect 12848 35876 12852 35932
rect 12852 35876 12908 35932
rect 12908 35876 12912 35932
rect 12848 35872 12912 35876
rect 12928 35932 12992 35936
rect 12928 35876 12932 35932
rect 12932 35876 12988 35932
rect 12988 35876 12992 35932
rect 12928 35872 12992 35876
rect 13008 35932 13072 35936
rect 13008 35876 13012 35932
rect 13012 35876 13068 35932
rect 13068 35876 13072 35932
rect 13008 35872 13072 35876
rect 13088 35932 13152 35936
rect 13088 35876 13092 35932
rect 13092 35876 13148 35932
rect 13148 35876 13152 35932
rect 13088 35872 13152 35876
rect 20778 35932 20842 35936
rect 20778 35876 20782 35932
rect 20782 35876 20838 35932
rect 20838 35876 20842 35932
rect 20778 35872 20842 35876
rect 20858 35932 20922 35936
rect 20858 35876 20862 35932
rect 20862 35876 20918 35932
rect 20918 35876 20922 35932
rect 20858 35872 20922 35876
rect 20938 35932 21002 35936
rect 20938 35876 20942 35932
rect 20942 35876 20998 35932
rect 20998 35876 21002 35932
rect 20938 35872 21002 35876
rect 21018 35932 21082 35936
rect 21018 35876 21022 35932
rect 21022 35876 21078 35932
rect 21078 35876 21082 35932
rect 21018 35872 21082 35876
rect 8882 35388 8946 35392
rect 8882 35332 8886 35388
rect 8886 35332 8942 35388
rect 8942 35332 8946 35388
rect 8882 35328 8946 35332
rect 8962 35388 9026 35392
rect 8962 35332 8966 35388
rect 8966 35332 9022 35388
rect 9022 35332 9026 35388
rect 8962 35328 9026 35332
rect 9042 35388 9106 35392
rect 9042 35332 9046 35388
rect 9046 35332 9102 35388
rect 9102 35332 9106 35388
rect 9042 35328 9106 35332
rect 9122 35388 9186 35392
rect 9122 35332 9126 35388
rect 9126 35332 9182 35388
rect 9182 35332 9186 35388
rect 9122 35328 9186 35332
rect 16813 35388 16877 35392
rect 16813 35332 16817 35388
rect 16817 35332 16873 35388
rect 16873 35332 16877 35388
rect 16813 35328 16877 35332
rect 16893 35388 16957 35392
rect 16893 35332 16897 35388
rect 16897 35332 16953 35388
rect 16953 35332 16957 35388
rect 16893 35328 16957 35332
rect 16973 35388 17037 35392
rect 16973 35332 16977 35388
rect 16977 35332 17033 35388
rect 17033 35332 17037 35388
rect 16973 35328 17037 35332
rect 17053 35388 17117 35392
rect 17053 35332 17057 35388
rect 17057 35332 17113 35388
rect 17113 35332 17117 35388
rect 17053 35328 17117 35332
rect 4917 34844 4981 34848
rect 4917 34788 4921 34844
rect 4921 34788 4977 34844
rect 4977 34788 4981 34844
rect 4917 34784 4981 34788
rect 4997 34844 5061 34848
rect 4997 34788 5001 34844
rect 5001 34788 5057 34844
rect 5057 34788 5061 34844
rect 4997 34784 5061 34788
rect 5077 34844 5141 34848
rect 5077 34788 5081 34844
rect 5081 34788 5137 34844
rect 5137 34788 5141 34844
rect 5077 34784 5141 34788
rect 5157 34844 5221 34848
rect 5157 34788 5161 34844
rect 5161 34788 5217 34844
rect 5217 34788 5221 34844
rect 5157 34784 5221 34788
rect 12848 34844 12912 34848
rect 12848 34788 12852 34844
rect 12852 34788 12908 34844
rect 12908 34788 12912 34844
rect 12848 34784 12912 34788
rect 12928 34844 12992 34848
rect 12928 34788 12932 34844
rect 12932 34788 12988 34844
rect 12988 34788 12992 34844
rect 12928 34784 12992 34788
rect 13008 34844 13072 34848
rect 13008 34788 13012 34844
rect 13012 34788 13068 34844
rect 13068 34788 13072 34844
rect 13008 34784 13072 34788
rect 13088 34844 13152 34848
rect 13088 34788 13092 34844
rect 13092 34788 13148 34844
rect 13148 34788 13152 34844
rect 13088 34784 13152 34788
rect 20778 34844 20842 34848
rect 20778 34788 20782 34844
rect 20782 34788 20838 34844
rect 20838 34788 20842 34844
rect 20778 34784 20842 34788
rect 20858 34844 20922 34848
rect 20858 34788 20862 34844
rect 20862 34788 20918 34844
rect 20918 34788 20922 34844
rect 20858 34784 20922 34788
rect 20938 34844 21002 34848
rect 20938 34788 20942 34844
rect 20942 34788 20998 34844
rect 20998 34788 21002 34844
rect 20938 34784 21002 34788
rect 21018 34844 21082 34848
rect 21018 34788 21022 34844
rect 21022 34788 21078 34844
rect 21078 34788 21082 34844
rect 21018 34784 21082 34788
rect 8882 34300 8946 34304
rect 8882 34244 8886 34300
rect 8886 34244 8942 34300
rect 8942 34244 8946 34300
rect 8882 34240 8946 34244
rect 8962 34300 9026 34304
rect 8962 34244 8966 34300
rect 8966 34244 9022 34300
rect 9022 34244 9026 34300
rect 8962 34240 9026 34244
rect 9042 34300 9106 34304
rect 9042 34244 9046 34300
rect 9046 34244 9102 34300
rect 9102 34244 9106 34300
rect 9042 34240 9106 34244
rect 9122 34300 9186 34304
rect 9122 34244 9126 34300
rect 9126 34244 9182 34300
rect 9182 34244 9186 34300
rect 9122 34240 9186 34244
rect 16813 34300 16877 34304
rect 16813 34244 16817 34300
rect 16817 34244 16873 34300
rect 16873 34244 16877 34300
rect 16813 34240 16877 34244
rect 16893 34300 16957 34304
rect 16893 34244 16897 34300
rect 16897 34244 16953 34300
rect 16953 34244 16957 34300
rect 16893 34240 16957 34244
rect 16973 34300 17037 34304
rect 16973 34244 16977 34300
rect 16977 34244 17033 34300
rect 17033 34244 17037 34300
rect 16973 34240 17037 34244
rect 17053 34300 17117 34304
rect 17053 34244 17057 34300
rect 17057 34244 17113 34300
rect 17113 34244 17117 34300
rect 17053 34240 17117 34244
rect 5396 34232 5460 34236
rect 5396 34176 5410 34232
rect 5410 34176 5460 34232
rect 5396 34172 5460 34176
rect 4917 33756 4981 33760
rect 4917 33700 4921 33756
rect 4921 33700 4977 33756
rect 4977 33700 4981 33756
rect 4917 33696 4981 33700
rect 4997 33756 5061 33760
rect 4997 33700 5001 33756
rect 5001 33700 5057 33756
rect 5057 33700 5061 33756
rect 4997 33696 5061 33700
rect 5077 33756 5141 33760
rect 5077 33700 5081 33756
rect 5081 33700 5137 33756
rect 5137 33700 5141 33756
rect 5077 33696 5141 33700
rect 5157 33756 5221 33760
rect 5157 33700 5161 33756
rect 5161 33700 5217 33756
rect 5217 33700 5221 33756
rect 5157 33696 5221 33700
rect 12848 33756 12912 33760
rect 12848 33700 12852 33756
rect 12852 33700 12908 33756
rect 12908 33700 12912 33756
rect 12848 33696 12912 33700
rect 12928 33756 12992 33760
rect 12928 33700 12932 33756
rect 12932 33700 12988 33756
rect 12988 33700 12992 33756
rect 12928 33696 12992 33700
rect 13008 33756 13072 33760
rect 13008 33700 13012 33756
rect 13012 33700 13068 33756
rect 13068 33700 13072 33756
rect 13008 33696 13072 33700
rect 13088 33756 13152 33760
rect 13088 33700 13092 33756
rect 13092 33700 13148 33756
rect 13148 33700 13152 33756
rect 13088 33696 13152 33700
rect 20778 33756 20842 33760
rect 20778 33700 20782 33756
rect 20782 33700 20838 33756
rect 20838 33700 20842 33756
rect 20778 33696 20842 33700
rect 20858 33756 20922 33760
rect 20858 33700 20862 33756
rect 20862 33700 20918 33756
rect 20918 33700 20922 33756
rect 20858 33696 20922 33700
rect 20938 33756 21002 33760
rect 20938 33700 20942 33756
rect 20942 33700 20998 33756
rect 20998 33700 21002 33756
rect 20938 33696 21002 33700
rect 21018 33756 21082 33760
rect 21018 33700 21022 33756
rect 21022 33700 21078 33756
rect 21078 33700 21082 33756
rect 21018 33696 21082 33700
rect 8882 33212 8946 33216
rect 8882 33156 8886 33212
rect 8886 33156 8942 33212
rect 8942 33156 8946 33212
rect 8882 33152 8946 33156
rect 8962 33212 9026 33216
rect 8962 33156 8966 33212
rect 8966 33156 9022 33212
rect 9022 33156 9026 33212
rect 8962 33152 9026 33156
rect 9042 33212 9106 33216
rect 9042 33156 9046 33212
rect 9046 33156 9102 33212
rect 9102 33156 9106 33212
rect 9042 33152 9106 33156
rect 9122 33212 9186 33216
rect 9122 33156 9126 33212
rect 9126 33156 9182 33212
rect 9182 33156 9186 33212
rect 9122 33152 9186 33156
rect 16813 33212 16877 33216
rect 16813 33156 16817 33212
rect 16817 33156 16873 33212
rect 16873 33156 16877 33212
rect 16813 33152 16877 33156
rect 16893 33212 16957 33216
rect 16893 33156 16897 33212
rect 16897 33156 16953 33212
rect 16953 33156 16957 33212
rect 16893 33152 16957 33156
rect 16973 33212 17037 33216
rect 16973 33156 16977 33212
rect 16977 33156 17033 33212
rect 17033 33156 17037 33212
rect 16973 33152 17037 33156
rect 17053 33212 17117 33216
rect 17053 33156 17057 33212
rect 17057 33156 17113 33212
rect 17113 33156 17117 33212
rect 17053 33152 17117 33156
rect 4917 32668 4981 32672
rect 4917 32612 4921 32668
rect 4921 32612 4977 32668
rect 4977 32612 4981 32668
rect 4917 32608 4981 32612
rect 4997 32668 5061 32672
rect 4997 32612 5001 32668
rect 5001 32612 5057 32668
rect 5057 32612 5061 32668
rect 4997 32608 5061 32612
rect 5077 32668 5141 32672
rect 5077 32612 5081 32668
rect 5081 32612 5137 32668
rect 5137 32612 5141 32668
rect 5077 32608 5141 32612
rect 5157 32668 5221 32672
rect 5157 32612 5161 32668
rect 5161 32612 5217 32668
rect 5217 32612 5221 32668
rect 5157 32608 5221 32612
rect 12848 32668 12912 32672
rect 12848 32612 12852 32668
rect 12852 32612 12908 32668
rect 12908 32612 12912 32668
rect 12848 32608 12912 32612
rect 12928 32668 12992 32672
rect 12928 32612 12932 32668
rect 12932 32612 12988 32668
rect 12988 32612 12992 32668
rect 12928 32608 12992 32612
rect 13008 32668 13072 32672
rect 13008 32612 13012 32668
rect 13012 32612 13068 32668
rect 13068 32612 13072 32668
rect 13008 32608 13072 32612
rect 13088 32668 13152 32672
rect 13088 32612 13092 32668
rect 13092 32612 13148 32668
rect 13148 32612 13152 32668
rect 13088 32608 13152 32612
rect 20778 32668 20842 32672
rect 20778 32612 20782 32668
rect 20782 32612 20838 32668
rect 20838 32612 20842 32668
rect 20778 32608 20842 32612
rect 20858 32668 20922 32672
rect 20858 32612 20862 32668
rect 20862 32612 20918 32668
rect 20918 32612 20922 32668
rect 20858 32608 20922 32612
rect 20938 32668 21002 32672
rect 20938 32612 20942 32668
rect 20942 32612 20998 32668
rect 20998 32612 21002 32668
rect 20938 32608 21002 32612
rect 21018 32668 21082 32672
rect 21018 32612 21022 32668
rect 21022 32612 21078 32668
rect 21078 32612 21082 32668
rect 21018 32608 21082 32612
rect 8882 32124 8946 32128
rect 8882 32068 8886 32124
rect 8886 32068 8942 32124
rect 8942 32068 8946 32124
rect 8882 32064 8946 32068
rect 8962 32124 9026 32128
rect 8962 32068 8966 32124
rect 8966 32068 9022 32124
rect 9022 32068 9026 32124
rect 8962 32064 9026 32068
rect 9042 32124 9106 32128
rect 9042 32068 9046 32124
rect 9046 32068 9102 32124
rect 9102 32068 9106 32124
rect 9042 32064 9106 32068
rect 9122 32124 9186 32128
rect 9122 32068 9126 32124
rect 9126 32068 9182 32124
rect 9182 32068 9186 32124
rect 9122 32064 9186 32068
rect 16813 32124 16877 32128
rect 16813 32068 16817 32124
rect 16817 32068 16873 32124
rect 16873 32068 16877 32124
rect 16813 32064 16877 32068
rect 16893 32124 16957 32128
rect 16893 32068 16897 32124
rect 16897 32068 16953 32124
rect 16953 32068 16957 32124
rect 16893 32064 16957 32068
rect 16973 32124 17037 32128
rect 16973 32068 16977 32124
rect 16977 32068 17033 32124
rect 17033 32068 17037 32124
rect 16973 32064 17037 32068
rect 17053 32124 17117 32128
rect 17053 32068 17057 32124
rect 17057 32068 17113 32124
rect 17113 32068 17117 32124
rect 17053 32064 17117 32068
rect 5396 31648 5460 31652
rect 5396 31592 5446 31648
rect 5446 31592 5460 31648
rect 5396 31588 5460 31592
rect 4917 31580 4981 31584
rect 4917 31524 4921 31580
rect 4921 31524 4977 31580
rect 4977 31524 4981 31580
rect 4917 31520 4981 31524
rect 4997 31580 5061 31584
rect 4997 31524 5001 31580
rect 5001 31524 5057 31580
rect 5057 31524 5061 31580
rect 4997 31520 5061 31524
rect 5077 31580 5141 31584
rect 5077 31524 5081 31580
rect 5081 31524 5137 31580
rect 5137 31524 5141 31580
rect 5077 31520 5141 31524
rect 5157 31580 5221 31584
rect 5157 31524 5161 31580
rect 5161 31524 5217 31580
rect 5217 31524 5221 31580
rect 5157 31520 5221 31524
rect 12848 31580 12912 31584
rect 12848 31524 12852 31580
rect 12852 31524 12908 31580
rect 12908 31524 12912 31580
rect 12848 31520 12912 31524
rect 12928 31580 12992 31584
rect 12928 31524 12932 31580
rect 12932 31524 12988 31580
rect 12988 31524 12992 31580
rect 12928 31520 12992 31524
rect 13008 31580 13072 31584
rect 13008 31524 13012 31580
rect 13012 31524 13068 31580
rect 13068 31524 13072 31580
rect 13008 31520 13072 31524
rect 13088 31580 13152 31584
rect 13088 31524 13092 31580
rect 13092 31524 13148 31580
rect 13148 31524 13152 31580
rect 13088 31520 13152 31524
rect 20778 31580 20842 31584
rect 20778 31524 20782 31580
rect 20782 31524 20838 31580
rect 20838 31524 20842 31580
rect 20778 31520 20842 31524
rect 20858 31580 20922 31584
rect 20858 31524 20862 31580
rect 20862 31524 20918 31580
rect 20918 31524 20922 31580
rect 20858 31520 20922 31524
rect 20938 31580 21002 31584
rect 20938 31524 20942 31580
rect 20942 31524 20998 31580
rect 20998 31524 21002 31580
rect 20938 31520 21002 31524
rect 21018 31580 21082 31584
rect 21018 31524 21022 31580
rect 21022 31524 21078 31580
rect 21078 31524 21082 31580
rect 21018 31520 21082 31524
rect 8882 31036 8946 31040
rect 8882 30980 8886 31036
rect 8886 30980 8942 31036
rect 8942 30980 8946 31036
rect 8882 30976 8946 30980
rect 8962 31036 9026 31040
rect 8962 30980 8966 31036
rect 8966 30980 9022 31036
rect 9022 30980 9026 31036
rect 8962 30976 9026 30980
rect 9042 31036 9106 31040
rect 9042 30980 9046 31036
rect 9046 30980 9102 31036
rect 9102 30980 9106 31036
rect 9042 30976 9106 30980
rect 9122 31036 9186 31040
rect 9122 30980 9126 31036
rect 9126 30980 9182 31036
rect 9182 30980 9186 31036
rect 9122 30976 9186 30980
rect 16813 31036 16877 31040
rect 16813 30980 16817 31036
rect 16817 30980 16873 31036
rect 16873 30980 16877 31036
rect 16813 30976 16877 30980
rect 16893 31036 16957 31040
rect 16893 30980 16897 31036
rect 16897 30980 16953 31036
rect 16953 30980 16957 31036
rect 16893 30976 16957 30980
rect 16973 31036 17037 31040
rect 16973 30980 16977 31036
rect 16977 30980 17033 31036
rect 17033 30980 17037 31036
rect 16973 30976 17037 30980
rect 17053 31036 17117 31040
rect 17053 30980 17057 31036
rect 17057 30980 17113 31036
rect 17113 30980 17117 31036
rect 17053 30976 17117 30980
rect 4917 30492 4981 30496
rect 4917 30436 4921 30492
rect 4921 30436 4977 30492
rect 4977 30436 4981 30492
rect 4917 30432 4981 30436
rect 4997 30492 5061 30496
rect 4997 30436 5001 30492
rect 5001 30436 5057 30492
rect 5057 30436 5061 30492
rect 4997 30432 5061 30436
rect 5077 30492 5141 30496
rect 5077 30436 5081 30492
rect 5081 30436 5137 30492
rect 5137 30436 5141 30492
rect 5077 30432 5141 30436
rect 5157 30492 5221 30496
rect 5157 30436 5161 30492
rect 5161 30436 5217 30492
rect 5217 30436 5221 30492
rect 5157 30432 5221 30436
rect 12848 30492 12912 30496
rect 12848 30436 12852 30492
rect 12852 30436 12908 30492
rect 12908 30436 12912 30492
rect 12848 30432 12912 30436
rect 12928 30492 12992 30496
rect 12928 30436 12932 30492
rect 12932 30436 12988 30492
rect 12988 30436 12992 30492
rect 12928 30432 12992 30436
rect 13008 30492 13072 30496
rect 13008 30436 13012 30492
rect 13012 30436 13068 30492
rect 13068 30436 13072 30492
rect 13008 30432 13072 30436
rect 13088 30492 13152 30496
rect 13088 30436 13092 30492
rect 13092 30436 13148 30492
rect 13148 30436 13152 30492
rect 13088 30432 13152 30436
rect 20778 30492 20842 30496
rect 20778 30436 20782 30492
rect 20782 30436 20838 30492
rect 20838 30436 20842 30492
rect 20778 30432 20842 30436
rect 20858 30492 20922 30496
rect 20858 30436 20862 30492
rect 20862 30436 20918 30492
rect 20918 30436 20922 30492
rect 20858 30432 20922 30436
rect 20938 30492 21002 30496
rect 20938 30436 20942 30492
rect 20942 30436 20998 30492
rect 20998 30436 21002 30492
rect 20938 30432 21002 30436
rect 21018 30492 21082 30496
rect 21018 30436 21022 30492
rect 21022 30436 21078 30492
rect 21078 30436 21082 30492
rect 21018 30432 21082 30436
rect 8882 29948 8946 29952
rect 8882 29892 8886 29948
rect 8886 29892 8942 29948
rect 8942 29892 8946 29948
rect 8882 29888 8946 29892
rect 8962 29948 9026 29952
rect 8962 29892 8966 29948
rect 8966 29892 9022 29948
rect 9022 29892 9026 29948
rect 8962 29888 9026 29892
rect 9042 29948 9106 29952
rect 9042 29892 9046 29948
rect 9046 29892 9102 29948
rect 9102 29892 9106 29948
rect 9042 29888 9106 29892
rect 9122 29948 9186 29952
rect 9122 29892 9126 29948
rect 9126 29892 9182 29948
rect 9182 29892 9186 29948
rect 9122 29888 9186 29892
rect 16813 29948 16877 29952
rect 16813 29892 16817 29948
rect 16817 29892 16873 29948
rect 16873 29892 16877 29948
rect 16813 29888 16877 29892
rect 16893 29948 16957 29952
rect 16893 29892 16897 29948
rect 16897 29892 16953 29948
rect 16953 29892 16957 29948
rect 16893 29888 16957 29892
rect 16973 29948 17037 29952
rect 16973 29892 16977 29948
rect 16977 29892 17033 29948
rect 17033 29892 17037 29948
rect 16973 29888 17037 29892
rect 17053 29948 17117 29952
rect 17053 29892 17057 29948
rect 17057 29892 17113 29948
rect 17113 29892 17117 29948
rect 17053 29888 17117 29892
rect 4917 29404 4981 29408
rect 4917 29348 4921 29404
rect 4921 29348 4977 29404
rect 4977 29348 4981 29404
rect 4917 29344 4981 29348
rect 4997 29404 5061 29408
rect 4997 29348 5001 29404
rect 5001 29348 5057 29404
rect 5057 29348 5061 29404
rect 4997 29344 5061 29348
rect 5077 29404 5141 29408
rect 5077 29348 5081 29404
rect 5081 29348 5137 29404
rect 5137 29348 5141 29404
rect 5077 29344 5141 29348
rect 5157 29404 5221 29408
rect 5157 29348 5161 29404
rect 5161 29348 5217 29404
rect 5217 29348 5221 29404
rect 5157 29344 5221 29348
rect 12848 29404 12912 29408
rect 12848 29348 12852 29404
rect 12852 29348 12908 29404
rect 12908 29348 12912 29404
rect 12848 29344 12912 29348
rect 12928 29404 12992 29408
rect 12928 29348 12932 29404
rect 12932 29348 12988 29404
rect 12988 29348 12992 29404
rect 12928 29344 12992 29348
rect 13008 29404 13072 29408
rect 13008 29348 13012 29404
rect 13012 29348 13068 29404
rect 13068 29348 13072 29404
rect 13008 29344 13072 29348
rect 13088 29404 13152 29408
rect 13088 29348 13092 29404
rect 13092 29348 13148 29404
rect 13148 29348 13152 29404
rect 13088 29344 13152 29348
rect 20778 29404 20842 29408
rect 20778 29348 20782 29404
rect 20782 29348 20838 29404
rect 20838 29348 20842 29404
rect 20778 29344 20842 29348
rect 20858 29404 20922 29408
rect 20858 29348 20862 29404
rect 20862 29348 20918 29404
rect 20918 29348 20922 29404
rect 20858 29344 20922 29348
rect 20938 29404 21002 29408
rect 20938 29348 20942 29404
rect 20942 29348 20998 29404
rect 20998 29348 21002 29404
rect 20938 29344 21002 29348
rect 21018 29404 21082 29408
rect 21018 29348 21022 29404
rect 21022 29348 21078 29404
rect 21078 29348 21082 29404
rect 21018 29344 21082 29348
rect 8882 28860 8946 28864
rect 8882 28804 8886 28860
rect 8886 28804 8942 28860
rect 8942 28804 8946 28860
rect 8882 28800 8946 28804
rect 8962 28860 9026 28864
rect 8962 28804 8966 28860
rect 8966 28804 9022 28860
rect 9022 28804 9026 28860
rect 8962 28800 9026 28804
rect 9042 28860 9106 28864
rect 9042 28804 9046 28860
rect 9046 28804 9102 28860
rect 9102 28804 9106 28860
rect 9042 28800 9106 28804
rect 9122 28860 9186 28864
rect 9122 28804 9126 28860
rect 9126 28804 9182 28860
rect 9182 28804 9186 28860
rect 9122 28800 9186 28804
rect 16813 28860 16877 28864
rect 16813 28804 16817 28860
rect 16817 28804 16873 28860
rect 16873 28804 16877 28860
rect 16813 28800 16877 28804
rect 16893 28860 16957 28864
rect 16893 28804 16897 28860
rect 16897 28804 16953 28860
rect 16953 28804 16957 28860
rect 16893 28800 16957 28804
rect 16973 28860 17037 28864
rect 16973 28804 16977 28860
rect 16977 28804 17033 28860
rect 17033 28804 17037 28860
rect 16973 28800 17037 28804
rect 17053 28860 17117 28864
rect 17053 28804 17057 28860
rect 17057 28804 17113 28860
rect 17113 28804 17117 28860
rect 17053 28800 17117 28804
rect 5396 28460 5460 28524
rect 8340 28520 8404 28524
rect 8340 28464 8354 28520
rect 8354 28464 8404 28520
rect 8340 28460 8404 28464
rect 4917 28316 4981 28320
rect 4917 28260 4921 28316
rect 4921 28260 4977 28316
rect 4977 28260 4981 28316
rect 4917 28256 4981 28260
rect 4997 28316 5061 28320
rect 4997 28260 5001 28316
rect 5001 28260 5057 28316
rect 5057 28260 5061 28316
rect 4997 28256 5061 28260
rect 5077 28316 5141 28320
rect 5077 28260 5081 28316
rect 5081 28260 5137 28316
rect 5137 28260 5141 28316
rect 5077 28256 5141 28260
rect 5157 28316 5221 28320
rect 5157 28260 5161 28316
rect 5161 28260 5217 28316
rect 5217 28260 5221 28316
rect 5157 28256 5221 28260
rect 12848 28316 12912 28320
rect 12848 28260 12852 28316
rect 12852 28260 12908 28316
rect 12908 28260 12912 28316
rect 12848 28256 12912 28260
rect 12928 28316 12992 28320
rect 12928 28260 12932 28316
rect 12932 28260 12988 28316
rect 12988 28260 12992 28316
rect 12928 28256 12992 28260
rect 13008 28316 13072 28320
rect 13008 28260 13012 28316
rect 13012 28260 13068 28316
rect 13068 28260 13072 28316
rect 13008 28256 13072 28260
rect 13088 28316 13152 28320
rect 13088 28260 13092 28316
rect 13092 28260 13148 28316
rect 13148 28260 13152 28316
rect 13088 28256 13152 28260
rect 20778 28316 20842 28320
rect 20778 28260 20782 28316
rect 20782 28260 20838 28316
rect 20838 28260 20842 28316
rect 20778 28256 20842 28260
rect 20858 28316 20922 28320
rect 20858 28260 20862 28316
rect 20862 28260 20918 28316
rect 20918 28260 20922 28316
rect 20858 28256 20922 28260
rect 20938 28316 21002 28320
rect 20938 28260 20942 28316
rect 20942 28260 20998 28316
rect 20998 28260 21002 28316
rect 20938 28256 21002 28260
rect 21018 28316 21082 28320
rect 21018 28260 21022 28316
rect 21022 28260 21078 28316
rect 21078 28260 21082 28316
rect 21018 28256 21082 28260
rect 8882 27772 8946 27776
rect 8882 27716 8886 27772
rect 8886 27716 8942 27772
rect 8942 27716 8946 27772
rect 8882 27712 8946 27716
rect 8962 27772 9026 27776
rect 8962 27716 8966 27772
rect 8966 27716 9022 27772
rect 9022 27716 9026 27772
rect 8962 27712 9026 27716
rect 9042 27772 9106 27776
rect 9042 27716 9046 27772
rect 9046 27716 9102 27772
rect 9102 27716 9106 27772
rect 9042 27712 9106 27716
rect 9122 27772 9186 27776
rect 9122 27716 9126 27772
rect 9126 27716 9182 27772
rect 9182 27716 9186 27772
rect 9122 27712 9186 27716
rect 16813 27772 16877 27776
rect 16813 27716 16817 27772
rect 16817 27716 16873 27772
rect 16873 27716 16877 27772
rect 16813 27712 16877 27716
rect 16893 27772 16957 27776
rect 16893 27716 16897 27772
rect 16897 27716 16953 27772
rect 16953 27716 16957 27772
rect 16893 27712 16957 27716
rect 16973 27772 17037 27776
rect 16973 27716 16977 27772
rect 16977 27716 17033 27772
rect 17033 27716 17037 27772
rect 16973 27712 17037 27716
rect 17053 27772 17117 27776
rect 17053 27716 17057 27772
rect 17057 27716 17113 27772
rect 17113 27716 17117 27772
rect 17053 27712 17117 27716
rect 9628 27236 9692 27300
rect 4917 27228 4981 27232
rect 4917 27172 4921 27228
rect 4921 27172 4977 27228
rect 4977 27172 4981 27228
rect 4917 27168 4981 27172
rect 4997 27228 5061 27232
rect 4997 27172 5001 27228
rect 5001 27172 5057 27228
rect 5057 27172 5061 27228
rect 4997 27168 5061 27172
rect 5077 27228 5141 27232
rect 5077 27172 5081 27228
rect 5081 27172 5137 27228
rect 5137 27172 5141 27228
rect 5077 27168 5141 27172
rect 5157 27228 5221 27232
rect 5157 27172 5161 27228
rect 5161 27172 5217 27228
rect 5217 27172 5221 27228
rect 5157 27168 5221 27172
rect 12848 27228 12912 27232
rect 12848 27172 12852 27228
rect 12852 27172 12908 27228
rect 12908 27172 12912 27228
rect 12848 27168 12912 27172
rect 12928 27228 12992 27232
rect 12928 27172 12932 27228
rect 12932 27172 12988 27228
rect 12988 27172 12992 27228
rect 12928 27168 12992 27172
rect 13008 27228 13072 27232
rect 13008 27172 13012 27228
rect 13012 27172 13068 27228
rect 13068 27172 13072 27228
rect 13008 27168 13072 27172
rect 13088 27228 13152 27232
rect 13088 27172 13092 27228
rect 13092 27172 13148 27228
rect 13148 27172 13152 27228
rect 13088 27168 13152 27172
rect 20778 27228 20842 27232
rect 20778 27172 20782 27228
rect 20782 27172 20838 27228
rect 20838 27172 20842 27228
rect 20778 27168 20842 27172
rect 20858 27228 20922 27232
rect 20858 27172 20862 27228
rect 20862 27172 20918 27228
rect 20918 27172 20922 27228
rect 20858 27168 20922 27172
rect 20938 27228 21002 27232
rect 20938 27172 20942 27228
rect 20942 27172 20998 27228
rect 20998 27172 21002 27228
rect 20938 27168 21002 27172
rect 21018 27228 21082 27232
rect 21018 27172 21022 27228
rect 21022 27172 21078 27228
rect 21078 27172 21082 27228
rect 21018 27168 21082 27172
rect 8524 26964 8588 27028
rect 10180 26964 10244 27028
rect 8708 26752 8772 26756
rect 8708 26696 8722 26752
rect 8722 26696 8772 26752
rect 8708 26692 8772 26696
rect 8882 26684 8946 26688
rect 8882 26628 8886 26684
rect 8886 26628 8942 26684
rect 8942 26628 8946 26684
rect 8882 26624 8946 26628
rect 8962 26684 9026 26688
rect 8962 26628 8966 26684
rect 8966 26628 9022 26684
rect 9022 26628 9026 26684
rect 8962 26624 9026 26628
rect 9042 26684 9106 26688
rect 9042 26628 9046 26684
rect 9046 26628 9102 26684
rect 9102 26628 9106 26684
rect 9042 26624 9106 26628
rect 9122 26684 9186 26688
rect 9122 26628 9126 26684
rect 9126 26628 9182 26684
rect 9182 26628 9186 26684
rect 9122 26624 9186 26628
rect 16813 26684 16877 26688
rect 16813 26628 16817 26684
rect 16817 26628 16873 26684
rect 16873 26628 16877 26684
rect 16813 26624 16877 26628
rect 16893 26684 16957 26688
rect 16893 26628 16897 26684
rect 16897 26628 16953 26684
rect 16953 26628 16957 26684
rect 16893 26624 16957 26628
rect 16973 26684 17037 26688
rect 16973 26628 16977 26684
rect 16977 26628 17033 26684
rect 17033 26628 17037 26684
rect 16973 26624 17037 26628
rect 17053 26684 17117 26688
rect 17053 26628 17057 26684
rect 17057 26628 17113 26684
rect 17113 26628 17117 26684
rect 17053 26624 17117 26628
rect 4917 26140 4981 26144
rect 4917 26084 4921 26140
rect 4921 26084 4977 26140
rect 4977 26084 4981 26140
rect 4917 26080 4981 26084
rect 4997 26140 5061 26144
rect 4997 26084 5001 26140
rect 5001 26084 5057 26140
rect 5057 26084 5061 26140
rect 4997 26080 5061 26084
rect 5077 26140 5141 26144
rect 5077 26084 5081 26140
rect 5081 26084 5137 26140
rect 5137 26084 5141 26140
rect 5077 26080 5141 26084
rect 5157 26140 5221 26144
rect 5157 26084 5161 26140
rect 5161 26084 5217 26140
rect 5217 26084 5221 26140
rect 5157 26080 5221 26084
rect 12848 26140 12912 26144
rect 12848 26084 12852 26140
rect 12852 26084 12908 26140
rect 12908 26084 12912 26140
rect 12848 26080 12912 26084
rect 12928 26140 12992 26144
rect 12928 26084 12932 26140
rect 12932 26084 12988 26140
rect 12988 26084 12992 26140
rect 12928 26080 12992 26084
rect 13008 26140 13072 26144
rect 13008 26084 13012 26140
rect 13012 26084 13068 26140
rect 13068 26084 13072 26140
rect 13008 26080 13072 26084
rect 13088 26140 13152 26144
rect 13088 26084 13092 26140
rect 13092 26084 13148 26140
rect 13148 26084 13152 26140
rect 13088 26080 13152 26084
rect 20778 26140 20842 26144
rect 20778 26084 20782 26140
rect 20782 26084 20838 26140
rect 20838 26084 20842 26140
rect 20778 26080 20842 26084
rect 20858 26140 20922 26144
rect 20858 26084 20862 26140
rect 20862 26084 20918 26140
rect 20918 26084 20922 26140
rect 20858 26080 20922 26084
rect 20938 26140 21002 26144
rect 20938 26084 20942 26140
rect 20942 26084 20998 26140
rect 20998 26084 21002 26140
rect 20938 26080 21002 26084
rect 21018 26140 21082 26144
rect 21018 26084 21022 26140
rect 21022 26084 21078 26140
rect 21078 26084 21082 26140
rect 21018 26080 21082 26084
rect 9444 26072 9508 26076
rect 9444 26016 9494 26072
rect 9494 26016 9508 26072
rect 9444 26012 9508 26016
rect 8882 25596 8946 25600
rect 8882 25540 8886 25596
rect 8886 25540 8942 25596
rect 8942 25540 8946 25596
rect 8882 25536 8946 25540
rect 8962 25596 9026 25600
rect 8962 25540 8966 25596
rect 8966 25540 9022 25596
rect 9022 25540 9026 25596
rect 8962 25536 9026 25540
rect 9042 25596 9106 25600
rect 9042 25540 9046 25596
rect 9046 25540 9102 25596
rect 9102 25540 9106 25596
rect 9042 25536 9106 25540
rect 9122 25596 9186 25600
rect 9122 25540 9126 25596
rect 9126 25540 9182 25596
rect 9182 25540 9186 25596
rect 9122 25536 9186 25540
rect 16813 25596 16877 25600
rect 16813 25540 16817 25596
rect 16817 25540 16873 25596
rect 16873 25540 16877 25596
rect 16813 25536 16877 25540
rect 16893 25596 16957 25600
rect 16893 25540 16897 25596
rect 16897 25540 16953 25596
rect 16953 25540 16957 25596
rect 16893 25536 16957 25540
rect 16973 25596 17037 25600
rect 16973 25540 16977 25596
rect 16977 25540 17033 25596
rect 17033 25540 17037 25596
rect 16973 25536 17037 25540
rect 17053 25596 17117 25600
rect 17053 25540 17057 25596
rect 17057 25540 17113 25596
rect 17113 25540 17117 25596
rect 17053 25536 17117 25540
rect 4917 25052 4981 25056
rect 4917 24996 4921 25052
rect 4921 24996 4977 25052
rect 4977 24996 4981 25052
rect 4917 24992 4981 24996
rect 4997 25052 5061 25056
rect 4997 24996 5001 25052
rect 5001 24996 5057 25052
rect 5057 24996 5061 25052
rect 4997 24992 5061 24996
rect 5077 25052 5141 25056
rect 5077 24996 5081 25052
rect 5081 24996 5137 25052
rect 5137 24996 5141 25052
rect 5077 24992 5141 24996
rect 5157 25052 5221 25056
rect 5157 24996 5161 25052
rect 5161 24996 5217 25052
rect 5217 24996 5221 25052
rect 5157 24992 5221 24996
rect 12848 25052 12912 25056
rect 12848 24996 12852 25052
rect 12852 24996 12908 25052
rect 12908 24996 12912 25052
rect 12848 24992 12912 24996
rect 12928 25052 12992 25056
rect 12928 24996 12932 25052
rect 12932 24996 12988 25052
rect 12988 24996 12992 25052
rect 12928 24992 12992 24996
rect 13008 25052 13072 25056
rect 13008 24996 13012 25052
rect 13012 24996 13068 25052
rect 13068 24996 13072 25052
rect 13008 24992 13072 24996
rect 13088 25052 13152 25056
rect 13088 24996 13092 25052
rect 13092 24996 13148 25052
rect 13148 24996 13152 25052
rect 13088 24992 13152 24996
rect 20778 25052 20842 25056
rect 20778 24996 20782 25052
rect 20782 24996 20838 25052
rect 20838 24996 20842 25052
rect 20778 24992 20842 24996
rect 20858 25052 20922 25056
rect 20858 24996 20862 25052
rect 20862 24996 20918 25052
rect 20918 24996 20922 25052
rect 20858 24992 20922 24996
rect 20938 25052 21002 25056
rect 20938 24996 20942 25052
rect 20942 24996 20998 25052
rect 20998 24996 21002 25052
rect 20938 24992 21002 24996
rect 21018 25052 21082 25056
rect 21018 24996 21022 25052
rect 21022 24996 21078 25052
rect 21078 24996 21082 25052
rect 21018 24992 21082 24996
rect 9260 24848 9324 24852
rect 9260 24792 9274 24848
rect 9274 24792 9324 24848
rect 9260 24788 9324 24792
rect 8882 24508 8946 24512
rect 8882 24452 8886 24508
rect 8886 24452 8942 24508
rect 8942 24452 8946 24508
rect 8882 24448 8946 24452
rect 8962 24508 9026 24512
rect 8962 24452 8966 24508
rect 8966 24452 9022 24508
rect 9022 24452 9026 24508
rect 8962 24448 9026 24452
rect 9042 24508 9106 24512
rect 9042 24452 9046 24508
rect 9046 24452 9102 24508
rect 9102 24452 9106 24508
rect 9042 24448 9106 24452
rect 9122 24508 9186 24512
rect 9122 24452 9126 24508
rect 9126 24452 9182 24508
rect 9182 24452 9186 24508
rect 9122 24448 9186 24452
rect 16813 24508 16877 24512
rect 16813 24452 16817 24508
rect 16817 24452 16873 24508
rect 16873 24452 16877 24508
rect 16813 24448 16877 24452
rect 16893 24508 16957 24512
rect 16893 24452 16897 24508
rect 16897 24452 16953 24508
rect 16953 24452 16957 24508
rect 16893 24448 16957 24452
rect 16973 24508 17037 24512
rect 16973 24452 16977 24508
rect 16977 24452 17033 24508
rect 17033 24452 17037 24508
rect 16973 24448 17037 24452
rect 17053 24508 17117 24512
rect 17053 24452 17057 24508
rect 17057 24452 17113 24508
rect 17113 24452 17117 24508
rect 17053 24448 17117 24452
rect 8524 24244 8588 24308
rect 4917 23964 4981 23968
rect 4917 23908 4921 23964
rect 4921 23908 4977 23964
rect 4977 23908 4981 23964
rect 4917 23904 4981 23908
rect 4997 23964 5061 23968
rect 4997 23908 5001 23964
rect 5001 23908 5057 23964
rect 5057 23908 5061 23964
rect 4997 23904 5061 23908
rect 5077 23964 5141 23968
rect 5077 23908 5081 23964
rect 5081 23908 5137 23964
rect 5137 23908 5141 23964
rect 5077 23904 5141 23908
rect 5157 23964 5221 23968
rect 5157 23908 5161 23964
rect 5161 23908 5217 23964
rect 5217 23908 5221 23964
rect 5157 23904 5221 23908
rect 12848 23964 12912 23968
rect 12848 23908 12852 23964
rect 12852 23908 12908 23964
rect 12908 23908 12912 23964
rect 12848 23904 12912 23908
rect 12928 23964 12992 23968
rect 12928 23908 12932 23964
rect 12932 23908 12988 23964
rect 12988 23908 12992 23964
rect 12928 23904 12992 23908
rect 13008 23964 13072 23968
rect 13008 23908 13012 23964
rect 13012 23908 13068 23964
rect 13068 23908 13072 23964
rect 13008 23904 13072 23908
rect 13088 23964 13152 23968
rect 13088 23908 13092 23964
rect 13092 23908 13148 23964
rect 13148 23908 13152 23964
rect 13088 23904 13152 23908
rect 20778 23964 20842 23968
rect 20778 23908 20782 23964
rect 20782 23908 20838 23964
rect 20838 23908 20842 23964
rect 20778 23904 20842 23908
rect 20858 23964 20922 23968
rect 20858 23908 20862 23964
rect 20862 23908 20918 23964
rect 20918 23908 20922 23964
rect 20858 23904 20922 23908
rect 20938 23964 21002 23968
rect 20938 23908 20942 23964
rect 20942 23908 20998 23964
rect 20998 23908 21002 23964
rect 20938 23904 21002 23908
rect 21018 23964 21082 23968
rect 21018 23908 21022 23964
rect 21022 23908 21078 23964
rect 21078 23908 21082 23964
rect 21018 23904 21082 23908
rect 8882 23420 8946 23424
rect 8882 23364 8886 23420
rect 8886 23364 8942 23420
rect 8942 23364 8946 23420
rect 8882 23360 8946 23364
rect 8962 23420 9026 23424
rect 8962 23364 8966 23420
rect 8966 23364 9022 23420
rect 9022 23364 9026 23420
rect 8962 23360 9026 23364
rect 9042 23420 9106 23424
rect 9042 23364 9046 23420
rect 9046 23364 9102 23420
rect 9102 23364 9106 23420
rect 9042 23360 9106 23364
rect 9122 23420 9186 23424
rect 9122 23364 9126 23420
rect 9126 23364 9182 23420
rect 9182 23364 9186 23420
rect 9122 23360 9186 23364
rect 16813 23420 16877 23424
rect 16813 23364 16817 23420
rect 16817 23364 16873 23420
rect 16873 23364 16877 23420
rect 16813 23360 16877 23364
rect 16893 23420 16957 23424
rect 16893 23364 16897 23420
rect 16897 23364 16953 23420
rect 16953 23364 16957 23420
rect 16893 23360 16957 23364
rect 16973 23420 17037 23424
rect 16973 23364 16977 23420
rect 16977 23364 17033 23420
rect 17033 23364 17037 23420
rect 16973 23360 17037 23364
rect 17053 23420 17117 23424
rect 17053 23364 17057 23420
rect 17057 23364 17113 23420
rect 17113 23364 17117 23420
rect 17053 23360 17117 23364
rect 5396 23080 5460 23084
rect 5396 23024 5410 23080
rect 5410 23024 5460 23080
rect 5396 23020 5460 23024
rect 4917 22876 4981 22880
rect 4917 22820 4921 22876
rect 4921 22820 4977 22876
rect 4977 22820 4981 22876
rect 4917 22816 4981 22820
rect 4997 22876 5061 22880
rect 4997 22820 5001 22876
rect 5001 22820 5057 22876
rect 5057 22820 5061 22876
rect 4997 22816 5061 22820
rect 5077 22876 5141 22880
rect 5077 22820 5081 22876
rect 5081 22820 5137 22876
rect 5137 22820 5141 22876
rect 5077 22816 5141 22820
rect 5157 22876 5221 22880
rect 5157 22820 5161 22876
rect 5161 22820 5217 22876
rect 5217 22820 5221 22876
rect 5157 22816 5221 22820
rect 12848 22876 12912 22880
rect 12848 22820 12852 22876
rect 12852 22820 12908 22876
rect 12908 22820 12912 22876
rect 12848 22816 12912 22820
rect 12928 22876 12992 22880
rect 12928 22820 12932 22876
rect 12932 22820 12988 22876
rect 12988 22820 12992 22876
rect 12928 22816 12992 22820
rect 13008 22876 13072 22880
rect 13008 22820 13012 22876
rect 13012 22820 13068 22876
rect 13068 22820 13072 22876
rect 13008 22816 13072 22820
rect 13088 22876 13152 22880
rect 13088 22820 13092 22876
rect 13092 22820 13148 22876
rect 13148 22820 13152 22876
rect 13088 22816 13152 22820
rect 20778 22876 20842 22880
rect 20778 22820 20782 22876
rect 20782 22820 20838 22876
rect 20838 22820 20842 22876
rect 20778 22816 20842 22820
rect 20858 22876 20922 22880
rect 20858 22820 20862 22876
rect 20862 22820 20918 22876
rect 20918 22820 20922 22876
rect 20858 22816 20922 22820
rect 20938 22876 21002 22880
rect 20938 22820 20942 22876
rect 20942 22820 20998 22876
rect 20998 22820 21002 22876
rect 20938 22816 21002 22820
rect 21018 22876 21082 22880
rect 21018 22820 21022 22876
rect 21022 22820 21078 22876
rect 21078 22820 21082 22876
rect 21018 22816 21082 22820
rect 7972 22808 8036 22812
rect 7972 22752 7986 22808
rect 7986 22752 8036 22808
rect 7972 22748 8036 22752
rect 8524 22672 8588 22676
rect 8524 22616 8538 22672
rect 8538 22616 8588 22672
rect 8524 22612 8588 22616
rect 8340 22476 8404 22540
rect 8882 22332 8946 22336
rect 8882 22276 8886 22332
rect 8886 22276 8942 22332
rect 8942 22276 8946 22332
rect 8882 22272 8946 22276
rect 8962 22332 9026 22336
rect 8962 22276 8966 22332
rect 8966 22276 9022 22332
rect 9022 22276 9026 22332
rect 8962 22272 9026 22276
rect 9042 22332 9106 22336
rect 9042 22276 9046 22332
rect 9046 22276 9102 22332
rect 9102 22276 9106 22332
rect 9042 22272 9106 22276
rect 9122 22332 9186 22336
rect 9122 22276 9126 22332
rect 9126 22276 9182 22332
rect 9182 22276 9186 22332
rect 9122 22272 9186 22276
rect 16813 22332 16877 22336
rect 16813 22276 16817 22332
rect 16817 22276 16873 22332
rect 16873 22276 16877 22332
rect 16813 22272 16877 22276
rect 16893 22332 16957 22336
rect 16893 22276 16897 22332
rect 16897 22276 16953 22332
rect 16953 22276 16957 22332
rect 16893 22272 16957 22276
rect 16973 22332 17037 22336
rect 16973 22276 16977 22332
rect 16977 22276 17033 22332
rect 17033 22276 17037 22332
rect 16973 22272 17037 22276
rect 17053 22332 17117 22336
rect 17053 22276 17057 22332
rect 17057 22276 17113 22332
rect 17113 22276 17117 22332
rect 17053 22272 17117 22276
rect 7052 21932 7116 21996
rect 9444 21992 9508 21996
rect 9444 21936 9494 21992
rect 9494 21936 9508 21992
rect 9444 21932 9508 21936
rect 7972 21796 8036 21860
rect 4917 21788 4981 21792
rect 4917 21732 4921 21788
rect 4921 21732 4977 21788
rect 4977 21732 4981 21788
rect 4917 21728 4981 21732
rect 4997 21788 5061 21792
rect 4997 21732 5001 21788
rect 5001 21732 5057 21788
rect 5057 21732 5061 21788
rect 4997 21728 5061 21732
rect 5077 21788 5141 21792
rect 5077 21732 5081 21788
rect 5081 21732 5137 21788
rect 5137 21732 5141 21788
rect 5077 21728 5141 21732
rect 5157 21788 5221 21792
rect 5157 21732 5161 21788
rect 5161 21732 5217 21788
rect 5217 21732 5221 21788
rect 5157 21728 5221 21732
rect 12848 21788 12912 21792
rect 12848 21732 12852 21788
rect 12852 21732 12908 21788
rect 12908 21732 12912 21788
rect 12848 21728 12912 21732
rect 12928 21788 12992 21792
rect 12928 21732 12932 21788
rect 12932 21732 12988 21788
rect 12988 21732 12992 21788
rect 12928 21728 12992 21732
rect 13008 21788 13072 21792
rect 13008 21732 13012 21788
rect 13012 21732 13068 21788
rect 13068 21732 13072 21788
rect 13008 21728 13072 21732
rect 13088 21788 13152 21792
rect 13088 21732 13092 21788
rect 13092 21732 13148 21788
rect 13148 21732 13152 21788
rect 13088 21728 13152 21732
rect 20778 21788 20842 21792
rect 20778 21732 20782 21788
rect 20782 21732 20838 21788
rect 20838 21732 20842 21788
rect 20778 21728 20842 21732
rect 20858 21788 20922 21792
rect 20858 21732 20862 21788
rect 20862 21732 20918 21788
rect 20918 21732 20922 21788
rect 20858 21728 20922 21732
rect 20938 21788 21002 21792
rect 20938 21732 20942 21788
rect 20942 21732 20998 21788
rect 20998 21732 21002 21788
rect 20938 21728 21002 21732
rect 21018 21788 21082 21792
rect 21018 21732 21022 21788
rect 21022 21732 21078 21788
rect 21078 21732 21082 21788
rect 21018 21728 21082 21732
rect 7420 21660 7484 21724
rect 6868 21524 6932 21588
rect 8882 21244 8946 21248
rect 8882 21188 8886 21244
rect 8886 21188 8942 21244
rect 8942 21188 8946 21244
rect 8882 21184 8946 21188
rect 8962 21244 9026 21248
rect 8962 21188 8966 21244
rect 8966 21188 9022 21244
rect 9022 21188 9026 21244
rect 8962 21184 9026 21188
rect 9042 21244 9106 21248
rect 9042 21188 9046 21244
rect 9046 21188 9102 21244
rect 9102 21188 9106 21244
rect 9042 21184 9106 21188
rect 9122 21244 9186 21248
rect 9122 21188 9126 21244
rect 9126 21188 9182 21244
rect 9182 21188 9186 21244
rect 9122 21184 9186 21188
rect 16813 21244 16877 21248
rect 16813 21188 16817 21244
rect 16817 21188 16873 21244
rect 16873 21188 16877 21244
rect 16813 21184 16877 21188
rect 16893 21244 16957 21248
rect 16893 21188 16897 21244
rect 16897 21188 16953 21244
rect 16953 21188 16957 21244
rect 16893 21184 16957 21188
rect 16973 21244 17037 21248
rect 16973 21188 16977 21244
rect 16977 21188 17033 21244
rect 17033 21188 17037 21244
rect 16973 21184 17037 21188
rect 17053 21244 17117 21248
rect 17053 21188 17057 21244
rect 17057 21188 17113 21244
rect 17113 21188 17117 21244
rect 17053 21184 17117 21188
rect 8708 20980 8772 21044
rect 8340 20768 8404 20772
rect 8340 20712 8390 20768
rect 8390 20712 8404 20768
rect 8340 20708 8404 20712
rect 4917 20700 4981 20704
rect 4917 20644 4921 20700
rect 4921 20644 4977 20700
rect 4977 20644 4981 20700
rect 4917 20640 4981 20644
rect 4997 20700 5061 20704
rect 4997 20644 5001 20700
rect 5001 20644 5057 20700
rect 5057 20644 5061 20700
rect 4997 20640 5061 20644
rect 5077 20700 5141 20704
rect 5077 20644 5081 20700
rect 5081 20644 5137 20700
rect 5137 20644 5141 20700
rect 5077 20640 5141 20644
rect 5157 20700 5221 20704
rect 5157 20644 5161 20700
rect 5161 20644 5217 20700
rect 5217 20644 5221 20700
rect 5157 20640 5221 20644
rect 12848 20700 12912 20704
rect 12848 20644 12852 20700
rect 12852 20644 12908 20700
rect 12908 20644 12912 20700
rect 12848 20640 12912 20644
rect 12928 20700 12992 20704
rect 12928 20644 12932 20700
rect 12932 20644 12988 20700
rect 12988 20644 12992 20700
rect 12928 20640 12992 20644
rect 13008 20700 13072 20704
rect 13008 20644 13012 20700
rect 13012 20644 13068 20700
rect 13068 20644 13072 20700
rect 13008 20640 13072 20644
rect 13088 20700 13152 20704
rect 13088 20644 13092 20700
rect 13092 20644 13148 20700
rect 13148 20644 13152 20700
rect 13088 20640 13152 20644
rect 20778 20700 20842 20704
rect 20778 20644 20782 20700
rect 20782 20644 20838 20700
rect 20838 20644 20842 20700
rect 20778 20640 20842 20644
rect 20858 20700 20922 20704
rect 20858 20644 20862 20700
rect 20862 20644 20918 20700
rect 20918 20644 20922 20700
rect 20858 20640 20922 20644
rect 20938 20700 21002 20704
rect 20938 20644 20942 20700
rect 20942 20644 20998 20700
rect 20998 20644 21002 20700
rect 20938 20640 21002 20644
rect 21018 20700 21082 20704
rect 21018 20644 21022 20700
rect 21022 20644 21078 20700
rect 21078 20644 21082 20700
rect 21018 20640 21082 20644
rect 9260 20436 9324 20500
rect 8882 20156 8946 20160
rect 8882 20100 8886 20156
rect 8886 20100 8942 20156
rect 8942 20100 8946 20156
rect 8882 20096 8946 20100
rect 8962 20156 9026 20160
rect 8962 20100 8966 20156
rect 8966 20100 9022 20156
rect 9022 20100 9026 20156
rect 8962 20096 9026 20100
rect 9042 20156 9106 20160
rect 9042 20100 9046 20156
rect 9046 20100 9102 20156
rect 9102 20100 9106 20156
rect 9042 20096 9106 20100
rect 9122 20156 9186 20160
rect 9122 20100 9126 20156
rect 9126 20100 9182 20156
rect 9182 20100 9186 20156
rect 9122 20096 9186 20100
rect 16813 20156 16877 20160
rect 16813 20100 16817 20156
rect 16817 20100 16873 20156
rect 16873 20100 16877 20156
rect 16813 20096 16877 20100
rect 16893 20156 16957 20160
rect 16893 20100 16897 20156
rect 16897 20100 16953 20156
rect 16953 20100 16957 20156
rect 16893 20096 16957 20100
rect 16973 20156 17037 20160
rect 16973 20100 16977 20156
rect 16977 20100 17033 20156
rect 17033 20100 17037 20156
rect 16973 20096 17037 20100
rect 17053 20156 17117 20160
rect 17053 20100 17057 20156
rect 17057 20100 17113 20156
rect 17113 20100 17117 20156
rect 17053 20096 17117 20100
rect 7052 19892 7116 19956
rect 9628 19756 9692 19820
rect 4917 19612 4981 19616
rect 4917 19556 4921 19612
rect 4921 19556 4977 19612
rect 4977 19556 4981 19612
rect 4917 19552 4981 19556
rect 4997 19612 5061 19616
rect 4997 19556 5001 19612
rect 5001 19556 5057 19612
rect 5057 19556 5061 19612
rect 4997 19552 5061 19556
rect 5077 19612 5141 19616
rect 5077 19556 5081 19612
rect 5081 19556 5137 19612
rect 5137 19556 5141 19612
rect 5077 19552 5141 19556
rect 5157 19612 5221 19616
rect 5157 19556 5161 19612
rect 5161 19556 5217 19612
rect 5217 19556 5221 19612
rect 5157 19552 5221 19556
rect 12848 19612 12912 19616
rect 12848 19556 12852 19612
rect 12852 19556 12908 19612
rect 12908 19556 12912 19612
rect 12848 19552 12912 19556
rect 12928 19612 12992 19616
rect 12928 19556 12932 19612
rect 12932 19556 12988 19612
rect 12988 19556 12992 19612
rect 12928 19552 12992 19556
rect 13008 19612 13072 19616
rect 13008 19556 13012 19612
rect 13012 19556 13068 19612
rect 13068 19556 13072 19612
rect 13008 19552 13072 19556
rect 13088 19612 13152 19616
rect 13088 19556 13092 19612
rect 13092 19556 13148 19612
rect 13148 19556 13152 19612
rect 13088 19552 13152 19556
rect 20778 19612 20842 19616
rect 20778 19556 20782 19612
rect 20782 19556 20838 19612
rect 20838 19556 20842 19612
rect 20778 19552 20842 19556
rect 20858 19612 20922 19616
rect 20858 19556 20862 19612
rect 20862 19556 20918 19612
rect 20918 19556 20922 19612
rect 20858 19552 20922 19556
rect 20938 19612 21002 19616
rect 20938 19556 20942 19612
rect 20942 19556 20998 19612
rect 20998 19556 21002 19612
rect 20938 19552 21002 19556
rect 21018 19612 21082 19616
rect 21018 19556 21022 19612
rect 21022 19556 21078 19612
rect 21078 19556 21082 19612
rect 21018 19552 21082 19556
rect 6868 19348 6932 19412
rect 10180 19076 10244 19140
rect 8882 19068 8946 19072
rect 8882 19012 8886 19068
rect 8886 19012 8942 19068
rect 8942 19012 8946 19068
rect 8882 19008 8946 19012
rect 8962 19068 9026 19072
rect 8962 19012 8966 19068
rect 8966 19012 9022 19068
rect 9022 19012 9026 19068
rect 8962 19008 9026 19012
rect 9042 19068 9106 19072
rect 9042 19012 9046 19068
rect 9046 19012 9102 19068
rect 9102 19012 9106 19068
rect 9042 19008 9106 19012
rect 9122 19068 9186 19072
rect 9122 19012 9126 19068
rect 9126 19012 9182 19068
rect 9182 19012 9186 19068
rect 9122 19008 9186 19012
rect 16813 19068 16877 19072
rect 16813 19012 16817 19068
rect 16817 19012 16873 19068
rect 16873 19012 16877 19068
rect 16813 19008 16877 19012
rect 16893 19068 16957 19072
rect 16893 19012 16897 19068
rect 16897 19012 16953 19068
rect 16953 19012 16957 19068
rect 16893 19008 16957 19012
rect 16973 19068 17037 19072
rect 16973 19012 16977 19068
rect 16977 19012 17033 19068
rect 17033 19012 17037 19068
rect 16973 19008 17037 19012
rect 17053 19068 17117 19072
rect 17053 19012 17057 19068
rect 17057 19012 17113 19068
rect 17113 19012 17117 19068
rect 17053 19008 17117 19012
rect 7420 19000 7484 19004
rect 7420 18944 7434 19000
rect 7434 18944 7484 19000
rect 7420 18940 7484 18944
rect 5396 18668 5460 18732
rect 4917 18524 4981 18528
rect 4917 18468 4921 18524
rect 4921 18468 4977 18524
rect 4977 18468 4981 18524
rect 4917 18464 4981 18468
rect 4997 18524 5061 18528
rect 4997 18468 5001 18524
rect 5001 18468 5057 18524
rect 5057 18468 5061 18524
rect 4997 18464 5061 18468
rect 5077 18524 5141 18528
rect 5077 18468 5081 18524
rect 5081 18468 5137 18524
rect 5137 18468 5141 18524
rect 5077 18464 5141 18468
rect 5157 18524 5221 18528
rect 5157 18468 5161 18524
rect 5161 18468 5217 18524
rect 5217 18468 5221 18524
rect 5157 18464 5221 18468
rect 12848 18524 12912 18528
rect 12848 18468 12852 18524
rect 12852 18468 12908 18524
rect 12908 18468 12912 18524
rect 12848 18464 12912 18468
rect 12928 18524 12992 18528
rect 12928 18468 12932 18524
rect 12932 18468 12988 18524
rect 12988 18468 12992 18524
rect 12928 18464 12992 18468
rect 13008 18524 13072 18528
rect 13008 18468 13012 18524
rect 13012 18468 13068 18524
rect 13068 18468 13072 18524
rect 13008 18464 13072 18468
rect 13088 18524 13152 18528
rect 13088 18468 13092 18524
rect 13092 18468 13148 18524
rect 13148 18468 13152 18524
rect 13088 18464 13152 18468
rect 20778 18524 20842 18528
rect 20778 18468 20782 18524
rect 20782 18468 20838 18524
rect 20838 18468 20842 18524
rect 20778 18464 20842 18468
rect 20858 18524 20922 18528
rect 20858 18468 20862 18524
rect 20862 18468 20918 18524
rect 20918 18468 20922 18524
rect 20858 18464 20922 18468
rect 20938 18524 21002 18528
rect 20938 18468 20942 18524
rect 20942 18468 20998 18524
rect 20998 18468 21002 18524
rect 20938 18464 21002 18468
rect 21018 18524 21082 18528
rect 21018 18468 21022 18524
rect 21022 18468 21078 18524
rect 21078 18468 21082 18524
rect 21018 18464 21082 18468
rect 8882 17980 8946 17984
rect 8882 17924 8886 17980
rect 8886 17924 8942 17980
rect 8942 17924 8946 17980
rect 8882 17920 8946 17924
rect 8962 17980 9026 17984
rect 8962 17924 8966 17980
rect 8966 17924 9022 17980
rect 9022 17924 9026 17980
rect 8962 17920 9026 17924
rect 9042 17980 9106 17984
rect 9042 17924 9046 17980
rect 9046 17924 9102 17980
rect 9102 17924 9106 17980
rect 9042 17920 9106 17924
rect 9122 17980 9186 17984
rect 9122 17924 9126 17980
rect 9126 17924 9182 17980
rect 9182 17924 9186 17980
rect 9122 17920 9186 17924
rect 16813 17980 16877 17984
rect 16813 17924 16817 17980
rect 16817 17924 16873 17980
rect 16873 17924 16877 17980
rect 16813 17920 16877 17924
rect 16893 17980 16957 17984
rect 16893 17924 16897 17980
rect 16897 17924 16953 17980
rect 16953 17924 16957 17980
rect 16893 17920 16957 17924
rect 16973 17980 17037 17984
rect 16973 17924 16977 17980
rect 16977 17924 17033 17980
rect 17033 17924 17037 17980
rect 16973 17920 17037 17924
rect 17053 17980 17117 17984
rect 17053 17924 17057 17980
rect 17057 17924 17113 17980
rect 17113 17924 17117 17980
rect 17053 17920 17117 17924
rect 4917 17436 4981 17440
rect 4917 17380 4921 17436
rect 4921 17380 4977 17436
rect 4977 17380 4981 17436
rect 4917 17376 4981 17380
rect 4997 17436 5061 17440
rect 4997 17380 5001 17436
rect 5001 17380 5057 17436
rect 5057 17380 5061 17436
rect 4997 17376 5061 17380
rect 5077 17436 5141 17440
rect 5077 17380 5081 17436
rect 5081 17380 5137 17436
rect 5137 17380 5141 17436
rect 5077 17376 5141 17380
rect 5157 17436 5221 17440
rect 5157 17380 5161 17436
rect 5161 17380 5217 17436
rect 5217 17380 5221 17436
rect 5157 17376 5221 17380
rect 12848 17436 12912 17440
rect 12848 17380 12852 17436
rect 12852 17380 12908 17436
rect 12908 17380 12912 17436
rect 12848 17376 12912 17380
rect 12928 17436 12992 17440
rect 12928 17380 12932 17436
rect 12932 17380 12988 17436
rect 12988 17380 12992 17436
rect 12928 17376 12992 17380
rect 13008 17436 13072 17440
rect 13008 17380 13012 17436
rect 13012 17380 13068 17436
rect 13068 17380 13072 17436
rect 13008 17376 13072 17380
rect 13088 17436 13152 17440
rect 13088 17380 13092 17436
rect 13092 17380 13148 17436
rect 13148 17380 13152 17436
rect 13088 17376 13152 17380
rect 20778 17436 20842 17440
rect 20778 17380 20782 17436
rect 20782 17380 20838 17436
rect 20838 17380 20842 17436
rect 20778 17376 20842 17380
rect 20858 17436 20922 17440
rect 20858 17380 20862 17436
rect 20862 17380 20918 17436
rect 20918 17380 20922 17436
rect 20858 17376 20922 17380
rect 20938 17436 21002 17440
rect 20938 17380 20942 17436
rect 20942 17380 20998 17436
rect 20998 17380 21002 17436
rect 20938 17376 21002 17380
rect 21018 17436 21082 17440
rect 21018 17380 21022 17436
rect 21022 17380 21078 17436
rect 21078 17380 21082 17436
rect 21018 17376 21082 17380
rect 8882 16892 8946 16896
rect 8882 16836 8886 16892
rect 8886 16836 8942 16892
rect 8942 16836 8946 16892
rect 8882 16832 8946 16836
rect 8962 16892 9026 16896
rect 8962 16836 8966 16892
rect 8966 16836 9022 16892
rect 9022 16836 9026 16892
rect 8962 16832 9026 16836
rect 9042 16892 9106 16896
rect 9042 16836 9046 16892
rect 9046 16836 9102 16892
rect 9102 16836 9106 16892
rect 9042 16832 9106 16836
rect 9122 16892 9186 16896
rect 9122 16836 9126 16892
rect 9126 16836 9182 16892
rect 9182 16836 9186 16892
rect 9122 16832 9186 16836
rect 16813 16892 16877 16896
rect 16813 16836 16817 16892
rect 16817 16836 16873 16892
rect 16873 16836 16877 16892
rect 16813 16832 16877 16836
rect 16893 16892 16957 16896
rect 16893 16836 16897 16892
rect 16897 16836 16953 16892
rect 16953 16836 16957 16892
rect 16893 16832 16957 16836
rect 16973 16892 17037 16896
rect 16973 16836 16977 16892
rect 16977 16836 17033 16892
rect 17033 16836 17037 16892
rect 16973 16832 17037 16836
rect 17053 16892 17117 16896
rect 17053 16836 17057 16892
rect 17057 16836 17113 16892
rect 17113 16836 17117 16892
rect 17053 16832 17117 16836
rect 4917 16348 4981 16352
rect 4917 16292 4921 16348
rect 4921 16292 4977 16348
rect 4977 16292 4981 16348
rect 4917 16288 4981 16292
rect 4997 16348 5061 16352
rect 4997 16292 5001 16348
rect 5001 16292 5057 16348
rect 5057 16292 5061 16348
rect 4997 16288 5061 16292
rect 5077 16348 5141 16352
rect 5077 16292 5081 16348
rect 5081 16292 5137 16348
rect 5137 16292 5141 16348
rect 5077 16288 5141 16292
rect 5157 16348 5221 16352
rect 5157 16292 5161 16348
rect 5161 16292 5217 16348
rect 5217 16292 5221 16348
rect 5157 16288 5221 16292
rect 12848 16348 12912 16352
rect 12848 16292 12852 16348
rect 12852 16292 12908 16348
rect 12908 16292 12912 16348
rect 12848 16288 12912 16292
rect 12928 16348 12992 16352
rect 12928 16292 12932 16348
rect 12932 16292 12988 16348
rect 12988 16292 12992 16348
rect 12928 16288 12992 16292
rect 13008 16348 13072 16352
rect 13008 16292 13012 16348
rect 13012 16292 13068 16348
rect 13068 16292 13072 16348
rect 13008 16288 13072 16292
rect 13088 16348 13152 16352
rect 13088 16292 13092 16348
rect 13092 16292 13148 16348
rect 13148 16292 13152 16348
rect 13088 16288 13152 16292
rect 20778 16348 20842 16352
rect 20778 16292 20782 16348
rect 20782 16292 20838 16348
rect 20838 16292 20842 16348
rect 20778 16288 20842 16292
rect 20858 16348 20922 16352
rect 20858 16292 20862 16348
rect 20862 16292 20918 16348
rect 20918 16292 20922 16348
rect 20858 16288 20922 16292
rect 20938 16348 21002 16352
rect 20938 16292 20942 16348
rect 20942 16292 20998 16348
rect 20998 16292 21002 16348
rect 20938 16288 21002 16292
rect 21018 16348 21082 16352
rect 21018 16292 21022 16348
rect 21022 16292 21078 16348
rect 21078 16292 21082 16348
rect 21018 16288 21082 16292
rect 8882 15804 8946 15808
rect 8882 15748 8886 15804
rect 8886 15748 8942 15804
rect 8942 15748 8946 15804
rect 8882 15744 8946 15748
rect 8962 15804 9026 15808
rect 8962 15748 8966 15804
rect 8966 15748 9022 15804
rect 9022 15748 9026 15804
rect 8962 15744 9026 15748
rect 9042 15804 9106 15808
rect 9042 15748 9046 15804
rect 9046 15748 9102 15804
rect 9102 15748 9106 15804
rect 9042 15744 9106 15748
rect 9122 15804 9186 15808
rect 9122 15748 9126 15804
rect 9126 15748 9182 15804
rect 9182 15748 9186 15804
rect 9122 15744 9186 15748
rect 16813 15804 16877 15808
rect 16813 15748 16817 15804
rect 16817 15748 16873 15804
rect 16873 15748 16877 15804
rect 16813 15744 16877 15748
rect 16893 15804 16957 15808
rect 16893 15748 16897 15804
rect 16897 15748 16953 15804
rect 16953 15748 16957 15804
rect 16893 15744 16957 15748
rect 16973 15804 17037 15808
rect 16973 15748 16977 15804
rect 16977 15748 17033 15804
rect 17033 15748 17037 15804
rect 16973 15744 17037 15748
rect 17053 15804 17117 15808
rect 17053 15748 17057 15804
rect 17057 15748 17113 15804
rect 17113 15748 17117 15804
rect 17053 15744 17117 15748
rect 4917 15260 4981 15264
rect 4917 15204 4921 15260
rect 4921 15204 4977 15260
rect 4977 15204 4981 15260
rect 4917 15200 4981 15204
rect 4997 15260 5061 15264
rect 4997 15204 5001 15260
rect 5001 15204 5057 15260
rect 5057 15204 5061 15260
rect 4997 15200 5061 15204
rect 5077 15260 5141 15264
rect 5077 15204 5081 15260
rect 5081 15204 5137 15260
rect 5137 15204 5141 15260
rect 5077 15200 5141 15204
rect 5157 15260 5221 15264
rect 5157 15204 5161 15260
rect 5161 15204 5217 15260
rect 5217 15204 5221 15260
rect 5157 15200 5221 15204
rect 12848 15260 12912 15264
rect 12848 15204 12852 15260
rect 12852 15204 12908 15260
rect 12908 15204 12912 15260
rect 12848 15200 12912 15204
rect 12928 15260 12992 15264
rect 12928 15204 12932 15260
rect 12932 15204 12988 15260
rect 12988 15204 12992 15260
rect 12928 15200 12992 15204
rect 13008 15260 13072 15264
rect 13008 15204 13012 15260
rect 13012 15204 13068 15260
rect 13068 15204 13072 15260
rect 13008 15200 13072 15204
rect 13088 15260 13152 15264
rect 13088 15204 13092 15260
rect 13092 15204 13148 15260
rect 13148 15204 13152 15260
rect 13088 15200 13152 15204
rect 20778 15260 20842 15264
rect 20778 15204 20782 15260
rect 20782 15204 20838 15260
rect 20838 15204 20842 15260
rect 20778 15200 20842 15204
rect 20858 15260 20922 15264
rect 20858 15204 20862 15260
rect 20862 15204 20918 15260
rect 20918 15204 20922 15260
rect 20858 15200 20922 15204
rect 20938 15260 21002 15264
rect 20938 15204 20942 15260
rect 20942 15204 20998 15260
rect 20998 15204 21002 15260
rect 20938 15200 21002 15204
rect 21018 15260 21082 15264
rect 21018 15204 21022 15260
rect 21022 15204 21078 15260
rect 21078 15204 21082 15260
rect 21018 15200 21082 15204
rect 8882 14716 8946 14720
rect 8882 14660 8886 14716
rect 8886 14660 8942 14716
rect 8942 14660 8946 14716
rect 8882 14656 8946 14660
rect 8962 14716 9026 14720
rect 8962 14660 8966 14716
rect 8966 14660 9022 14716
rect 9022 14660 9026 14716
rect 8962 14656 9026 14660
rect 9042 14716 9106 14720
rect 9042 14660 9046 14716
rect 9046 14660 9102 14716
rect 9102 14660 9106 14716
rect 9042 14656 9106 14660
rect 9122 14716 9186 14720
rect 9122 14660 9126 14716
rect 9126 14660 9182 14716
rect 9182 14660 9186 14716
rect 9122 14656 9186 14660
rect 16813 14716 16877 14720
rect 16813 14660 16817 14716
rect 16817 14660 16873 14716
rect 16873 14660 16877 14716
rect 16813 14656 16877 14660
rect 16893 14716 16957 14720
rect 16893 14660 16897 14716
rect 16897 14660 16953 14716
rect 16953 14660 16957 14716
rect 16893 14656 16957 14660
rect 16973 14716 17037 14720
rect 16973 14660 16977 14716
rect 16977 14660 17033 14716
rect 17033 14660 17037 14716
rect 16973 14656 17037 14660
rect 17053 14716 17117 14720
rect 17053 14660 17057 14716
rect 17057 14660 17113 14716
rect 17113 14660 17117 14716
rect 17053 14656 17117 14660
rect 4917 14172 4981 14176
rect 4917 14116 4921 14172
rect 4921 14116 4977 14172
rect 4977 14116 4981 14172
rect 4917 14112 4981 14116
rect 4997 14172 5061 14176
rect 4997 14116 5001 14172
rect 5001 14116 5057 14172
rect 5057 14116 5061 14172
rect 4997 14112 5061 14116
rect 5077 14172 5141 14176
rect 5077 14116 5081 14172
rect 5081 14116 5137 14172
rect 5137 14116 5141 14172
rect 5077 14112 5141 14116
rect 5157 14172 5221 14176
rect 5157 14116 5161 14172
rect 5161 14116 5217 14172
rect 5217 14116 5221 14172
rect 5157 14112 5221 14116
rect 12848 14172 12912 14176
rect 12848 14116 12852 14172
rect 12852 14116 12908 14172
rect 12908 14116 12912 14172
rect 12848 14112 12912 14116
rect 12928 14172 12992 14176
rect 12928 14116 12932 14172
rect 12932 14116 12988 14172
rect 12988 14116 12992 14172
rect 12928 14112 12992 14116
rect 13008 14172 13072 14176
rect 13008 14116 13012 14172
rect 13012 14116 13068 14172
rect 13068 14116 13072 14172
rect 13008 14112 13072 14116
rect 13088 14172 13152 14176
rect 13088 14116 13092 14172
rect 13092 14116 13148 14172
rect 13148 14116 13152 14172
rect 13088 14112 13152 14116
rect 20778 14172 20842 14176
rect 20778 14116 20782 14172
rect 20782 14116 20838 14172
rect 20838 14116 20842 14172
rect 20778 14112 20842 14116
rect 20858 14172 20922 14176
rect 20858 14116 20862 14172
rect 20862 14116 20918 14172
rect 20918 14116 20922 14172
rect 20858 14112 20922 14116
rect 20938 14172 21002 14176
rect 20938 14116 20942 14172
rect 20942 14116 20998 14172
rect 20998 14116 21002 14172
rect 20938 14112 21002 14116
rect 21018 14172 21082 14176
rect 21018 14116 21022 14172
rect 21022 14116 21078 14172
rect 21078 14116 21082 14172
rect 21018 14112 21082 14116
rect 8882 13628 8946 13632
rect 8882 13572 8886 13628
rect 8886 13572 8942 13628
rect 8942 13572 8946 13628
rect 8882 13568 8946 13572
rect 8962 13628 9026 13632
rect 8962 13572 8966 13628
rect 8966 13572 9022 13628
rect 9022 13572 9026 13628
rect 8962 13568 9026 13572
rect 9042 13628 9106 13632
rect 9042 13572 9046 13628
rect 9046 13572 9102 13628
rect 9102 13572 9106 13628
rect 9042 13568 9106 13572
rect 9122 13628 9186 13632
rect 9122 13572 9126 13628
rect 9126 13572 9182 13628
rect 9182 13572 9186 13628
rect 9122 13568 9186 13572
rect 16813 13628 16877 13632
rect 16813 13572 16817 13628
rect 16817 13572 16873 13628
rect 16873 13572 16877 13628
rect 16813 13568 16877 13572
rect 16893 13628 16957 13632
rect 16893 13572 16897 13628
rect 16897 13572 16953 13628
rect 16953 13572 16957 13628
rect 16893 13568 16957 13572
rect 16973 13628 17037 13632
rect 16973 13572 16977 13628
rect 16977 13572 17033 13628
rect 17033 13572 17037 13628
rect 16973 13568 17037 13572
rect 17053 13628 17117 13632
rect 17053 13572 17057 13628
rect 17057 13572 17113 13628
rect 17113 13572 17117 13628
rect 17053 13568 17117 13572
rect 9444 13152 9508 13156
rect 9444 13096 9458 13152
rect 9458 13096 9508 13152
rect 9444 13092 9508 13096
rect 4917 13084 4981 13088
rect 4917 13028 4921 13084
rect 4921 13028 4977 13084
rect 4977 13028 4981 13084
rect 4917 13024 4981 13028
rect 4997 13084 5061 13088
rect 4997 13028 5001 13084
rect 5001 13028 5057 13084
rect 5057 13028 5061 13084
rect 4997 13024 5061 13028
rect 5077 13084 5141 13088
rect 5077 13028 5081 13084
rect 5081 13028 5137 13084
rect 5137 13028 5141 13084
rect 5077 13024 5141 13028
rect 5157 13084 5221 13088
rect 5157 13028 5161 13084
rect 5161 13028 5217 13084
rect 5217 13028 5221 13084
rect 5157 13024 5221 13028
rect 12848 13084 12912 13088
rect 12848 13028 12852 13084
rect 12852 13028 12908 13084
rect 12908 13028 12912 13084
rect 12848 13024 12912 13028
rect 12928 13084 12992 13088
rect 12928 13028 12932 13084
rect 12932 13028 12988 13084
rect 12988 13028 12992 13084
rect 12928 13024 12992 13028
rect 13008 13084 13072 13088
rect 13008 13028 13012 13084
rect 13012 13028 13068 13084
rect 13068 13028 13072 13084
rect 13008 13024 13072 13028
rect 13088 13084 13152 13088
rect 13088 13028 13092 13084
rect 13092 13028 13148 13084
rect 13148 13028 13152 13084
rect 13088 13024 13152 13028
rect 20778 13084 20842 13088
rect 20778 13028 20782 13084
rect 20782 13028 20838 13084
rect 20838 13028 20842 13084
rect 20778 13024 20842 13028
rect 20858 13084 20922 13088
rect 20858 13028 20862 13084
rect 20862 13028 20918 13084
rect 20918 13028 20922 13084
rect 20858 13024 20922 13028
rect 20938 13084 21002 13088
rect 20938 13028 20942 13084
rect 20942 13028 20998 13084
rect 20998 13028 21002 13084
rect 20938 13024 21002 13028
rect 21018 13084 21082 13088
rect 21018 13028 21022 13084
rect 21022 13028 21078 13084
rect 21078 13028 21082 13084
rect 21018 13024 21082 13028
rect 5396 12820 5460 12884
rect 8882 12540 8946 12544
rect 8882 12484 8886 12540
rect 8886 12484 8942 12540
rect 8942 12484 8946 12540
rect 8882 12480 8946 12484
rect 8962 12540 9026 12544
rect 8962 12484 8966 12540
rect 8966 12484 9022 12540
rect 9022 12484 9026 12540
rect 8962 12480 9026 12484
rect 9042 12540 9106 12544
rect 9042 12484 9046 12540
rect 9046 12484 9102 12540
rect 9102 12484 9106 12540
rect 9042 12480 9106 12484
rect 9122 12540 9186 12544
rect 9122 12484 9126 12540
rect 9126 12484 9182 12540
rect 9182 12484 9186 12540
rect 9122 12480 9186 12484
rect 16813 12540 16877 12544
rect 16813 12484 16817 12540
rect 16817 12484 16873 12540
rect 16873 12484 16877 12540
rect 16813 12480 16877 12484
rect 16893 12540 16957 12544
rect 16893 12484 16897 12540
rect 16897 12484 16953 12540
rect 16953 12484 16957 12540
rect 16893 12480 16957 12484
rect 16973 12540 17037 12544
rect 16973 12484 16977 12540
rect 16977 12484 17033 12540
rect 17033 12484 17037 12540
rect 16973 12480 17037 12484
rect 17053 12540 17117 12544
rect 17053 12484 17057 12540
rect 17057 12484 17113 12540
rect 17113 12484 17117 12540
rect 17053 12480 17117 12484
rect 4917 11996 4981 12000
rect 4917 11940 4921 11996
rect 4921 11940 4977 11996
rect 4977 11940 4981 11996
rect 4917 11936 4981 11940
rect 4997 11996 5061 12000
rect 4997 11940 5001 11996
rect 5001 11940 5057 11996
rect 5057 11940 5061 11996
rect 4997 11936 5061 11940
rect 5077 11996 5141 12000
rect 5077 11940 5081 11996
rect 5081 11940 5137 11996
rect 5137 11940 5141 11996
rect 5077 11936 5141 11940
rect 5157 11996 5221 12000
rect 5157 11940 5161 11996
rect 5161 11940 5217 11996
rect 5217 11940 5221 11996
rect 5157 11936 5221 11940
rect 12848 11996 12912 12000
rect 12848 11940 12852 11996
rect 12852 11940 12908 11996
rect 12908 11940 12912 11996
rect 12848 11936 12912 11940
rect 12928 11996 12992 12000
rect 12928 11940 12932 11996
rect 12932 11940 12988 11996
rect 12988 11940 12992 11996
rect 12928 11936 12992 11940
rect 13008 11996 13072 12000
rect 13008 11940 13012 11996
rect 13012 11940 13068 11996
rect 13068 11940 13072 11996
rect 13008 11936 13072 11940
rect 13088 11996 13152 12000
rect 13088 11940 13092 11996
rect 13092 11940 13148 11996
rect 13148 11940 13152 11996
rect 13088 11936 13152 11940
rect 20778 11996 20842 12000
rect 20778 11940 20782 11996
rect 20782 11940 20838 11996
rect 20838 11940 20842 11996
rect 20778 11936 20842 11940
rect 20858 11996 20922 12000
rect 20858 11940 20862 11996
rect 20862 11940 20918 11996
rect 20918 11940 20922 11996
rect 20858 11936 20922 11940
rect 20938 11996 21002 12000
rect 20938 11940 20942 11996
rect 20942 11940 20998 11996
rect 20998 11940 21002 11996
rect 20938 11936 21002 11940
rect 21018 11996 21082 12000
rect 21018 11940 21022 11996
rect 21022 11940 21078 11996
rect 21078 11940 21082 11996
rect 21018 11936 21082 11940
rect 8882 11452 8946 11456
rect 8882 11396 8886 11452
rect 8886 11396 8942 11452
rect 8942 11396 8946 11452
rect 8882 11392 8946 11396
rect 8962 11452 9026 11456
rect 8962 11396 8966 11452
rect 8966 11396 9022 11452
rect 9022 11396 9026 11452
rect 8962 11392 9026 11396
rect 9042 11452 9106 11456
rect 9042 11396 9046 11452
rect 9046 11396 9102 11452
rect 9102 11396 9106 11452
rect 9042 11392 9106 11396
rect 9122 11452 9186 11456
rect 9122 11396 9126 11452
rect 9126 11396 9182 11452
rect 9182 11396 9186 11452
rect 9122 11392 9186 11396
rect 16813 11452 16877 11456
rect 16813 11396 16817 11452
rect 16817 11396 16873 11452
rect 16873 11396 16877 11452
rect 16813 11392 16877 11396
rect 16893 11452 16957 11456
rect 16893 11396 16897 11452
rect 16897 11396 16953 11452
rect 16953 11396 16957 11452
rect 16893 11392 16957 11396
rect 16973 11452 17037 11456
rect 16973 11396 16977 11452
rect 16977 11396 17033 11452
rect 17033 11396 17037 11452
rect 16973 11392 17037 11396
rect 17053 11452 17117 11456
rect 17053 11396 17057 11452
rect 17057 11396 17113 11452
rect 17113 11396 17117 11452
rect 17053 11392 17117 11396
rect 4917 10908 4981 10912
rect 4917 10852 4921 10908
rect 4921 10852 4977 10908
rect 4977 10852 4981 10908
rect 4917 10848 4981 10852
rect 4997 10908 5061 10912
rect 4997 10852 5001 10908
rect 5001 10852 5057 10908
rect 5057 10852 5061 10908
rect 4997 10848 5061 10852
rect 5077 10908 5141 10912
rect 5077 10852 5081 10908
rect 5081 10852 5137 10908
rect 5137 10852 5141 10908
rect 5077 10848 5141 10852
rect 5157 10908 5221 10912
rect 5157 10852 5161 10908
rect 5161 10852 5217 10908
rect 5217 10852 5221 10908
rect 5157 10848 5221 10852
rect 12848 10908 12912 10912
rect 12848 10852 12852 10908
rect 12852 10852 12908 10908
rect 12908 10852 12912 10908
rect 12848 10848 12912 10852
rect 12928 10908 12992 10912
rect 12928 10852 12932 10908
rect 12932 10852 12988 10908
rect 12988 10852 12992 10908
rect 12928 10848 12992 10852
rect 13008 10908 13072 10912
rect 13008 10852 13012 10908
rect 13012 10852 13068 10908
rect 13068 10852 13072 10908
rect 13008 10848 13072 10852
rect 13088 10908 13152 10912
rect 13088 10852 13092 10908
rect 13092 10852 13148 10908
rect 13148 10852 13152 10908
rect 13088 10848 13152 10852
rect 20778 10908 20842 10912
rect 20778 10852 20782 10908
rect 20782 10852 20838 10908
rect 20838 10852 20842 10908
rect 20778 10848 20842 10852
rect 20858 10908 20922 10912
rect 20858 10852 20862 10908
rect 20862 10852 20918 10908
rect 20918 10852 20922 10908
rect 20858 10848 20922 10852
rect 20938 10908 21002 10912
rect 20938 10852 20942 10908
rect 20942 10852 20998 10908
rect 20998 10852 21002 10908
rect 20938 10848 21002 10852
rect 21018 10908 21082 10912
rect 21018 10852 21022 10908
rect 21022 10852 21078 10908
rect 21078 10852 21082 10908
rect 21018 10848 21082 10852
rect 8882 10364 8946 10368
rect 8882 10308 8886 10364
rect 8886 10308 8942 10364
rect 8942 10308 8946 10364
rect 8882 10304 8946 10308
rect 8962 10364 9026 10368
rect 8962 10308 8966 10364
rect 8966 10308 9022 10364
rect 9022 10308 9026 10364
rect 8962 10304 9026 10308
rect 9042 10364 9106 10368
rect 9042 10308 9046 10364
rect 9046 10308 9102 10364
rect 9102 10308 9106 10364
rect 9042 10304 9106 10308
rect 9122 10364 9186 10368
rect 9122 10308 9126 10364
rect 9126 10308 9182 10364
rect 9182 10308 9186 10364
rect 9122 10304 9186 10308
rect 16813 10364 16877 10368
rect 16813 10308 16817 10364
rect 16817 10308 16873 10364
rect 16873 10308 16877 10364
rect 16813 10304 16877 10308
rect 16893 10364 16957 10368
rect 16893 10308 16897 10364
rect 16897 10308 16953 10364
rect 16953 10308 16957 10364
rect 16893 10304 16957 10308
rect 16973 10364 17037 10368
rect 16973 10308 16977 10364
rect 16977 10308 17033 10364
rect 17033 10308 17037 10364
rect 16973 10304 17037 10308
rect 17053 10364 17117 10368
rect 17053 10308 17057 10364
rect 17057 10308 17113 10364
rect 17113 10308 17117 10364
rect 17053 10304 17117 10308
rect 7236 10236 7300 10300
rect 12204 9828 12268 9892
rect 4917 9820 4981 9824
rect 4917 9764 4921 9820
rect 4921 9764 4977 9820
rect 4977 9764 4981 9820
rect 4917 9760 4981 9764
rect 4997 9820 5061 9824
rect 4997 9764 5001 9820
rect 5001 9764 5057 9820
rect 5057 9764 5061 9820
rect 4997 9760 5061 9764
rect 5077 9820 5141 9824
rect 5077 9764 5081 9820
rect 5081 9764 5137 9820
rect 5137 9764 5141 9820
rect 5077 9760 5141 9764
rect 5157 9820 5221 9824
rect 5157 9764 5161 9820
rect 5161 9764 5217 9820
rect 5217 9764 5221 9820
rect 5157 9760 5221 9764
rect 12848 9820 12912 9824
rect 12848 9764 12852 9820
rect 12852 9764 12908 9820
rect 12908 9764 12912 9820
rect 12848 9760 12912 9764
rect 12928 9820 12992 9824
rect 12928 9764 12932 9820
rect 12932 9764 12988 9820
rect 12988 9764 12992 9820
rect 12928 9760 12992 9764
rect 13008 9820 13072 9824
rect 13008 9764 13012 9820
rect 13012 9764 13068 9820
rect 13068 9764 13072 9820
rect 13008 9760 13072 9764
rect 13088 9820 13152 9824
rect 13088 9764 13092 9820
rect 13092 9764 13148 9820
rect 13148 9764 13152 9820
rect 13088 9760 13152 9764
rect 20778 9820 20842 9824
rect 20778 9764 20782 9820
rect 20782 9764 20838 9820
rect 20838 9764 20842 9820
rect 20778 9760 20842 9764
rect 20858 9820 20922 9824
rect 20858 9764 20862 9820
rect 20862 9764 20918 9820
rect 20918 9764 20922 9820
rect 20858 9760 20922 9764
rect 20938 9820 21002 9824
rect 20938 9764 20942 9820
rect 20942 9764 20998 9820
rect 20998 9764 21002 9820
rect 20938 9760 21002 9764
rect 21018 9820 21082 9824
rect 21018 9764 21022 9820
rect 21022 9764 21078 9820
rect 21078 9764 21082 9820
rect 21018 9760 21082 9764
rect 13308 9284 13372 9348
rect 8882 9276 8946 9280
rect 8882 9220 8886 9276
rect 8886 9220 8942 9276
rect 8942 9220 8946 9276
rect 8882 9216 8946 9220
rect 8962 9276 9026 9280
rect 8962 9220 8966 9276
rect 8966 9220 9022 9276
rect 9022 9220 9026 9276
rect 8962 9216 9026 9220
rect 9042 9276 9106 9280
rect 9042 9220 9046 9276
rect 9046 9220 9102 9276
rect 9102 9220 9106 9276
rect 9042 9216 9106 9220
rect 9122 9276 9186 9280
rect 9122 9220 9126 9276
rect 9126 9220 9182 9276
rect 9182 9220 9186 9276
rect 9122 9216 9186 9220
rect 16813 9276 16877 9280
rect 16813 9220 16817 9276
rect 16817 9220 16873 9276
rect 16873 9220 16877 9276
rect 16813 9216 16877 9220
rect 16893 9276 16957 9280
rect 16893 9220 16897 9276
rect 16897 9220 16953 9276
rect 16953 9220 16957 9276
rect 16893 9216 16957 9220
rect 16973 9276 17037 9280
rect 16973 9220 16977 9276
rect 16977 9220 17033 9276
rect 17033 9220 17037 9276
rect 16973 9216 17037 9220
rect 17053 9276 17117 9280
rect 17053 9220 17057 9276
rect 17057 9220 17113 9276
rect 17113 9220 17117 9276
rect 17053 9216 17117 9220
rect 5396 9012 5460 9076
rect 12572 9012 12636 9076
rect 4917 8732 4981 8736
rect 4917 8676 4921 8732
rect 4921 8676 4977 8732
rect 4977 8676 4981 8732
rect 4917 8672 4981 8676
rect 4997 8732 5061 8736
rect 4997 8676 5001 8732
rect 5001 8676 5057 8732
rect 5057 8676 5061 8732
rect 4997 8672 5061 8676
rect 5077 8732 5141 8736
rect 5077 8676 5081 8732
rect 5081 8676 5137 8732
rect 5137 8676 5141 8732
rect 5077 8672 5141 8676
rect 5157 8732 5221 8736
rect 5157 8676 5161 8732
rect 5161 8676 5217 8732
rect 5217 8676 5221 8732
rect 5157 8672 5221 8676
rect 12848 8732 12912 8736
rect 12848 8676 12852 8732
rect 12852 8676 12908 8732
rect 12908 8676 12912 8732
rect 12848 8672 12912 8676
rect 12928 8732 12992 8736
rect 12928 8676 12932 8732
rect 12932 8676 12988 8732
rect 12988 8676 12992 8732
rect 12928 8672 12992 8676
rect 13008 8732 13072 8736
rect 13008 8676 13012 8732
rect 13012 8676 13068 8732
rect 13068 8676 13072 8732
rect 13008 8672 13072 8676
rect 13088 8732 13152 8736
rect 13088 8676 13092 8732
rect 13092 8676 13148 8732
rect 13148 8676 13152 8732
rect 13088 8672 13152 8676
rect 20778 8732 20842 8736
rect 20778 8676 20782 8732
rect 20782 8676 20838 8732
rect 20838 8676 20842 8732
rect 20778 8672 20842 8676
rect 20858 8732 20922 8736
rect 20858 8676 20862 8732
rect 20862 8676 20918 8732
rect 20918 8676 20922 8732
rect 20858 8672 20922 8676
rect 20938 8732 21002 8736
rect 20938 8676 20942 8732
rect 20942 8676 20998 8732
rect 20998 8676 21002 8732
rect 20938 8672 21002 8676
rect 21018 8732 21082 8736
rect 21018 8676 21022 8732
rect 21022 8676 21078 8732
rect 21078 8676 21082 8732
rect 21018 8672 21082 8676
rect 12572 8468 12636 8532
rect 13308 8332 13372 8396
rect 13492 8196 13556 8260
rect 8882 8188 8946 8192
rect 8882 8132 8886 8188
rect 8886 8132 8942 8188
rect 8942 8132 8946 8188
rect 8882 8128 8946 8132
rect 8962 8188 9026 8192
rect 8962 8132 8966 8188
rect 8966 8132 9022 8188
rect 9022 8132 9026 8188
rect 8962 8128 9026 8132
rect 9042 8188 9106 8192
rect 9042 8132 9046 8188
rect 9046 8132 9102 8188
rect 9102 8132 9106 8188
rect 9042 8128 9106 8132
rect 9122 8188 9186 8192
rect 9122 8132 9126 8188
rect 9126 8132 9182 8188
rect 9182 8132 9186 8188
rect 9122 8128 9186 8132
rect 16813 8188 16877 8192
rect 16813 8132 16817 8188
rect 16817 8132 16873 8188
rect 16873 8132 16877 8188
rect 16813 8128 16877 8132
rect 16893 8188 16957 8192
rect 16893 8132 16897 8188
rect 16897 8132 16953 8188
rect 16953 8132 16957 8188
rect 16893 8128 16957 8132
rect 16973 8188 17037 8192
rect 16973 8132 16977 8188
rect 16977 8132 17033 8188
rect 17033 8132 17037 8188
rect 16973 8128 17037 8132
rect 17053 8188 17117 8192
rect 17053 8132 17057 8188
rect 17057 8132 17113 8188
rect 17113 8132 17117 8188
rect 17053 8128 17117 8132
rect 7236 7848 7300 7852
rect 7236 7792 7286 7848
rect 7286 7792 7300 7848
rect 7236 7788 7300 7792
rect 4917 7644 4981 7648
rect 4917 7588 4921 7644
rect 4921 7588 4977 7644
rect 4977 7588 4981 7644
rect 4917 7584 4981 7588
rect 4997 7644 5061 7648
rect 4997 7588 5001 7644
rect 5001 7588 5057 7644
rect 5057 7588 5061 7644
rect 4997 7584 5061 7588
rect 5077 7644 5141 7648
rect 5077 7588 5081 7644
rect 5081 7588 5137 7644
rect 5137 7588 5141 7644
rect 5077 7584 5141 7588
rect 5157 7644 5221 7648
rect 5157 7588 5161 7644
rect 5161 7588 5217 7644
rect 5217 7588 5221 7644
rect 5157 7584 5221 7588
rect 12848 7644 12912 7648
rect 12848 7588 12852 7644
rect 12852 7588 12908 7644
rect 12908 7588 12912 7644
rect 12848 7584 12912 7588
rect 12928 7644 12992 7648
rect 12928 7588 12932 7644
rect 12932 7588 12988 7644
rect 12988 7588 12992 7644
rect 12928 7584 12992 7588
rect 13008 7644 13072 7648
rect 13008 7588 13012 7644
rect 13012 7588 13068 7644
rect 13068 7588 13072 7644
rect 13008 7584 13072 7588
rect 13088 7644 13152 7648
rect 13088 7588 13092 7644
rect 13092 7588 13148 7644
rect 13148 7588 13152 7644
rect 13088 7584 13152 7588
rect 20778 7644 20842 7648
rect 20778 7588 20782 7644
rect 20782 7588 20838 7644
rect 20838 7588 20842 7644
rect 20778 7584 20842 7588
rect 20858 7644 20922 7648
rect 20858 7588 20862 7644
rect 20862 7588 20918 7644
rect 20918 7588 20922 7644
rect 20858 7584 20922 7588
rect 20938 7644 21002 7648
rect 20938 7588 20942 7644
rect 20942 7588 20998 7644
rect 20998 7588 21002 7644
rect 20938 7584 21002 7588
rect 21018 7644 21082 7648
rect 21018 7588 21022 7644
rect 21022 7588 21078 7644
rect 21078 7588 21082 7644
rect 21018 7584 21082 7588
rect 8882 7100 8946 7104
rect 8882 7044 8886 7100
rect 8886 7044 8942 7100
rect 8942 7044 8946 7100
rect 8882 7040 8946 7044
rect 8962 7100 9026 7104
rect 8962 7044 8966 7100
rect 8966 7044 9022 7100
rect 9022 7044 9026 7100
rect 8962 7040 9026 7044
rect 9042 7100 9106 7104
rect 9042 7044 9046 7100
rect 9046 7044 9102 7100
rect 9102 7044 9106 7100
rect 9042 7040 9106 7044
rect 9122 7100 9186 7104
rect 9122 7044 9126 7100
rect 9126 7044 9182 7100
rect 9182 7044 9186 7100
rect 9122 7040 9186 7044
rect 16813 7100 16877 7104
rect 16813 7044 16817 7100
rect 16817 7044 16873 7100
rect 16873 7044 16877 7100
rect 16813 7040 16877 7044
rect 16893 7100 16957 7104
rect 16893 7044 16897 7100
rect 16897 7044 16953 7100
rect 16953 7044 16957 7100
rect 16893 7040 16957 7044
rect 16973 7100 17037 7104
rect 16973 7044 16977 7100
rect 16977 7044 17033 7100
rect 17033 7044 17037 7100
rect 16973 7040 17037 7044
rect 17053 7100 17117 7104
rect 17053 7044 17057 7100
rect 17057 7044 17113 7100
rect 17113 7044 17117 7100
rect 17053 7040 17117 7044
rect 4917 6556 4981 6560
rect 4917 6500 4921 6556
rect 4921 6500 4977 6556
rect 4977 6500 4981 6556
rect 4917 6496 4981 6500
rect 4997 6556 5061 6560
rect 4997 6500 5001 6556
rect 5001 6500 5057 6556
rect 5057 6500 5061 6556
rect 4997 6496 5061 6500
rect 5077 6556 5141 6560
rect 5077 6500 5081 6556
rect 5081 6500 5137 6556
rect 5137 6500 5141 6556
rect 5077 6496 5141 6500
rect 5157 6556 5221 6560
rect 5157 6500 5161 6556
rect 5161 6500 5217 6556
rect 5217 6500 5221 6556
rect 5157 6496 5221 6500
rect 12848 6556 12912 6560
rect 12848 6500 12852 6556
rect 12852 6500 12908 6556
rect 12908 6500 12912 6556
rect 12848 6496 12912 6500
rect 12928 6556 12992 6560
rect 12928 6500 12932 6556
rect 12932 6500 12988 6556
rect 12988 6500 12992 6556
rect 12928 6496 12992 6500
rect 13008 6556 13072 6560
rect 13008 6500 13012 6556
rect 13012 6500 13068 6556
rect 13068 6500 13072 6556
rect 13008 6496 13072 6500
rect 13088 6556 13152 6560
rect 13088 6500 13092 6556
rect 13092 6500 13148 6556
rect 13148 6500 13152 6556
rect 13088 6496 13152 6500
rect 20778 6556 20842 6560
rect 20778 6500 20782 6556
rect 20782 6500 20838 6556
rect 20838 6500 20842 6556
rect 20778 6496 20842 6500
rect 20858 6556 20922 6560
rect 20858 6500 20862 6556
rect 20862 6500 20918 6556
rect 20918 6500 20922 6556
rect 20858 6496 20922 6500
rect 20938 6556 21002 6560
rect 20938 6500 20942 6556
rect 20942 6500 20998 6556
rect 20998 6500 21002 6556
rect 20938 6496 21002 6500
rect 21018 6556 21082 6560
rect 21018 6500 21022 6556
rect 21022 6500 21078 6556
rect 21078 6500 21082 6556
rect 21018 6496 21082 6500
rect 8882 6012 8946 6016
rect 8882 5956 8886 6012
rect 8886 5956 8942 6012
rect 8942 5956 8946 6012
rect 8882 5952 8946 5956
rect 8962 6012 9026 6016
rect 8962 5956 8966 6012
rect 8966 5956 9022 6012
rect 9022 5956 9026 6012
rect 8962 5952 9026 5956
rect 9042 6012 9106 6016
rect 9042 5956 9046 6012
rect 9046 5956 9102 6012
rect 9102 5956 9106 6012
rect 9042 5952 9106 5956
rect 9122 6012 9186 6016
rect 9122 5956 9126 6012
rect 9126 5956 9182 6012
rect 9182 5956 9186 6012
rect 9122 5952 9186 5956
rect 16813 6012 16877 6016
rect 16813 5956 16817 6012
rect 16817 5956 16873 6012
rect 16873 5956 16877 6012
rect 16813 5952 16877 5956
rect 16893 6012 16957 6016
rect 16893 5956 16897 6012
rect 16897 5956 16953 6012
rect 16953 5956 16957 6012
rect 16893 5952 16957 5956
rect 16973 6012 17037 6016
rect 16973 5956 16977 6012
rect 16977 5956 17033 6012
rect 17033 5956 17037 6012
rect 16973 5952 17037 5956
rect 17053 6012 17117 6016
rect 17053 5956 17057 6012
rect 17057 5956 17113 6012
rect 17113 5956 17117 6012
rect 17053 5952 17117 5956
rect 4917 5468 4981 5472
rect 4917 5412 4921 5468
rect 4921 5412 4977 5468
rect 4977 5412 4981 5468
rect 4917 5408 4981 5412
rect 4997 5468 5061 5472
rect 4997 5412 5001 5468
rect 5001 5412 5057 5468
rect 5057 5412 5061 5468
rect 4997 5408 5061 5412
rect 5077 5468 5141 5472
rect 5077 5412 5081 5468
rect 5081 5412 5137 5468
rect 5137 5412 5141 5468
rect 5077 5408 5141 5412
rect 5157 5468 5221 5472
rect 5157 5412 5161 5468
rect 5161 5412 5217 5468
rect 5217 5412 5221 5468
rect 5157 5408 5221 5412
rect 12848 5468 12912 5472
rect 12848 5412 12852 5468
rect 12852 5412 12908 5468
rect 12908 5412 12912 5468
rect 12848 5408 12912 5412
rect 12928 5468 12992 5472
rect 12928 5412 12932 5468
rect 12932 5412 12988 5468
rect 12988 5412 12992 5468
rect 12928 5408 12992 5412
rect 13008 5468 13072 5472
rect 13008 5412 13012 5468
rect 13012 5412 13068 5468
rect 13068 5412 13072 5468
rect 13008 5408 13072 5412
rect 13088 5468 13152 5472
rect 13088 5412 13092 5468
rect 13092 5412 13148 5468
rect 13148 5412 13152 5468
rect 13088 5408 13152 5412
rect 20778 5468 20842 5472
rect 20778 5412 20782 5468
rect 20782 5412 20838 5468
rect 20838 5412 20842 5468
rect 20778 5408 20842 5412
rect 20858 5468 20922 5472
rect 20858 5412 20862 5468
rect 20862 5412 20918 5468
rect 20918 5412 20922 5468
rect 20858 5408 20922 5412
rect 20938 5468 21002 5472
rect 20938 5412 20942 5468
rect 20942 5412 20998 5468
rect 20998 5412 21002 5468
rect 20938 5408 21002 5412
rect 21018 5468 21082 5472
rect 21018 5412 21022 5468
rect 21022 5412 21078 5468
rect 21078 5412 21082 5468
rect 21018 5408 21082 5412
rect 8882 4924 8946 4928
rect 8882 4868 8886 4924
rect 8886 4868 8942 4924
rect 8942 4868 8946 4924
rect 8882 4864 8946 4868
rect 8962 4924 9026 4928
rect 8962 4868 8966 4924
rect 8966 4868 9022 4924
rect 9022 4868 9026 4924
rect 8962 4864 9026 4868
rect 9042 4924 9106 4928
rect 9042 4868 9046 4924
rect 9046 4868 9102 4924
rect 9102 4868 9106 4924
rect 9042 4864 9106 4868
rect 9122 4924 9186 4928
rect 9122 4868 9126 4924
rect 9126 4868 9182 4924
rect 9182 4868 9186 4924
rect 9122 4864 9186 4868
rect 16813 4924 16877 4928
rect 16813 4868 16817 4924
rect 16817 4868 16873 4924
rect 16873 4868 16877 4924
rect 16813 4864 16877 4868
rect 16893 4924 16957 4928
rect 16893 4868 16897 4924
rect 16897 4868 16953 4924
rect 16953 4868 16957 4924
rect 16893 4864 16957 4868
rect 16973 4924 17037 4928
rect 16973 4868 16977 4924
rect 16977 4868 17033 4924
rect 17033 4868 17037 4924
rect 16973 4864 17037 4868
rect 17053 4924 17117 4928
rect 17053 4868 17057 4924
rect 17057 4868 17113 4924
rect 17113 4868 17117 4924
rect 17053 4864 17117 4868
rect 12204 4448 12268 4452
rect 12204 4392 12218 4448
rect 12218 4392 12268 4448
rect 12204 4388 12268 4392
rect 4917 4380 4981 4384
rect 4917 4324 4921 4380
rect 4921 4324 4977 4380
rect 4977 4324 4981 4380
rect 4917 4320 4981 4324
rect 4997 4380 5061 4384
rect 4997 4324 5001 4380
rect 5001 4324 5057 4380
rect 5057 4324 5061 4380
rect 4997 4320 5061 4324
rect 5077 4380 5141 4384
rect 5077 4324 5081 4380
rect 5081 4324 5137 4380
rect 5137 4324 5141 4380
rect 5077 4320 5141 4324
rect 5157 4380 5221 4384
rect 5157 4324 5161 4380
rect 5161 4324 5217 4380
rect 5217 4324 5221 4380
rect 5157 4320 5221 4324
rect 12848 4380 12912 4384
rect 12848 4324 12852 4380
rect 12852 4324 12908 4380
rect 12908 4324 12912 4380
rect 12848 4320 12912 4324
rect 12928 4380 12992 4384
rect 12928 4324 12932 4380
rect 12932 4324 12988 4380
rect 12988 4324 12992 4380
rect 12928 4320 12992 4324
rect 13008 4380 13072 4384
rect 13008 4324 13012 4380
rect 13012 4324 13068 4380
rect 13068 4324 13072 4380
rect 13008 4320 13072 4324
rect 13088 4380 13152 4384
rect 13088 4324 13092 4380
rect 13092 4324 13148 4380
rect 13148 4324 13152 4380
rect 13088 4320 13152 4324
rect 20778 4380 20842 4384
rect 20778 4324 20782 4380
rect 20782 4324 20838 4380
rect 20838 4324 20842 4380
rect 20778 4320 20842 4324
rect 20858 4380 20922 4384
rect 20858 4324 20862 4380
rect 20862 4324 20918 4380
rect 20918 4324 20922 4380
rect 20858 4320 20922 4324
rect 20938 4380 21002 4384
rect 20938 4324 20942 4380
rect 20942 4324 20998 4380
rect 20998 4324 21002 4380
rect 20938 4320 21002 4324
rect 21018 4380 21082 4384
rect 21018 4324 21022 4380
rect 21022 4324 21078 4380
rect 21078 4324 21082 4380
rect 21018 4320 21082 4324
rect 13492 4116 13556 4180
rect 8882 3836 8946 3840
rect 8882 3780 8886 3836
rect 8886 3780 8942 3836
rect 8942 3780 8946 3836
rect 8882 3776 8946 3780
rect 8962 3836 9026 3840
rect 8962 3780 8966 3836
rect 8966 3780 9022 3836
rect 9022 3780 9026 3836
rect 8962 3776 9026 3780
rect 9042 3836 9106 3840
rect 9042 3780 9046 3836
rect 9046 3780 9102 3836
rect 9102 3780 9106 3836
rect 9042 3776 9106 3780
rect 9122 3836 9186 3840
rect 9122 3780 9126 3836
rect 9126 3780 9182 3836
rect 9182 3780 9186 3836
rect 9122 3776 9186 3780
rect 16813 3836 16877 3840
rect 16813 3780 16817 3836
rect 16817 3780 16873 3836
rect 16873 3780 16877 3836
rect 16813 3776 16877 3780
rect 16893 3836 16957 3840
rect 16893 3780 16897 3836
rect 16897 3780 16953 3836
rect 16953 3780 16957 3836
rect 16893 3776 16957 3780
rect 16973 3836 17037 3840
rect 16973 3780 16977 3836
rect 16977 3780 17033 3836
rect 17033 3780 17037 3836
rect 16973 3776 17037 3780
rect 17053 3836 17117 3840
rect 17053 3780 17057 3836
rect 17057 3780 17113 3836
rect 17113 3780 17117 3836
rect 17053 3776 17117 3780
rect 4917 3292 4981 3296
rect 4917 3236 4921 3292
rect 4921 3236 4977 3292
rect 4977 3236 4981 3292
rect 4917 3232 4981 3236
rect 4997 3292 5061 3296
rect 4997 3236 5001 3292
rect 5001 3236 5057 3292
rect 5057 3236 5061 3292
rect 4997 3232 5061 3236
rect 5077 3292 5141 3296
rect 5077 3236 5081 3292
rect 5081 3236 5137 3292
rect 5137 3236 5141 3292
rect 5077 3232 5141 3236
rect 5157 3292 5221 3296
rect 5157 3236 5161 3292
rect 5161 3236 5217 3292
rect 5217 3236 5221 3292
rect 5157 3232 5221 3236
rect 12848 3292 12912 3296
rect 12848 3236 12852 3292
rect 12852 3236 12908 3292
rect 12908 3236 12912 3292
rect 12848 3232 12912 3236
rect 12928 3292 12992 3296
rect 12928 3236 12932 3292
rect 12932 3236 12988 3292
rect 12988 3236 12992 3292
rect 12928 3232 12992 3236
rect 13008 3292 13072 3296
rect 13008 3236 13012 3292
rect 13012 3236 13068 3292
rect 13068 3236 13072 3292
rect 13008 3232 13072 3236
rect 13088 3292 13152 3296
rect 13088 3236 13092 3292
rect 13092 3236 13148 3292
rect 13148 3236 13152 3292
rect 13088 3232 13152 3236
rect 20778 3292 20842 3296
rect 20778 3236 20782 3292
rect 20782 3236 20838 3292
rect 20838 3236 20842 3292
rect 20778 3232 20842 3236
rect 20858 3292 20922 3296
rect 20858 3236 20862 3292
rect 20862 3236 20918 3292
rect 20918 3236 20922 3292
rect 20858 3232 20922 3236
rect 20938 3292 21002 3296
rect 20938 3236 20942 3292
rect 20942 3236 20998 3292
rect 20998 3236 21002 3292
rect 20938 3232 21002 3236
rect 21018 3292 21082 3296
rect 21018 3236 21022 3292
rect 21022 3236 21078 3292
rect 21078 3236 21082 3292
rect 21018 3232 21082 3236
rect 9444 3164 9508 3228
rect 8882 2748 8946 2752
rect 8882 2692 8886 2748
rect 8886 2692 8942 2748
rect 8942 2692 8946 2748
rect 8882 2688 8946 2692
rect 8962 2748 9026 2752
rect 8962 2692 8966 2748
rect 8966 2692 9022 2748
rect 9022 2692 9026 2748
rect 8962 2688 9026 2692
rect 9042 2748 9106 2752
rect 9042 2692 9046 2748
rect 9046 2692 9102 2748
rect 9102 2692 9106 2748
rect 9042 2688 9106 2692
rect 9122 2748 9186 2752
rect 9122 2692 9126 2748
rect 9126 2692 9182 2748
rect 9182 2692 9186 2748
rect 9122 2688 9186 2692
rect 16813 2748 16877 2752
rect 16813 2692 16817 2748
rect 16817 2692 16873 2748
rect 16873 2692 16877 2748
rect 16813 2688 16877 2692
rect 16893 2748 16957 2752
rect 16893 2692 16897 2748
rect 16897 2692 16953 2748
rect 16953 2692 16957 2748
rect 16893 2688 16957 2692
rect 16973 2748 17037 2752
rect 16973 2692 16977 2748
rect 16977 2692 17033 2748
rect 17033 2692 17037 2748
rect 16973 2688 17037 2692
rect 17053 2748 17117 2752
rect 17053 2692 17057 2748
rect 17057 2692 17113 2748
rect 17113 2692 17117 2748
rect 17053 2688 17117 2692
rect 4917 2204 4981 2208
rect 4917 2148 4921 2204
rect 4921 2148 4977 2204
rect 4977 2148 4981 2204
rect 4917 2144 4981 2148
rect 4997 2204 5061 2208
rect 4997 2148 5001 2204
rect 5001 2148 5057 2204
rect 5057 2148 5061 2204
rect 4997 2144 5061 2148
rect 5077 2204 5141 2208
rect 5077 2148 5081 2204
rect 5081 2148 5137 2204
rect 5137 2148 5141 2204
rect 5077 2144 5141 2148
rect 5157 2204 5221 2208
rect 5157 2148 5161 2204
rect 5161 2148 5217 2204
rect 5217 2148 5221 2204
rect 5157 2144 5221 2148
rect 12848 2204 12912 2208
rect 12848 2148 12852 2204
rect 12852 2148 12908 2204
rect 12908 2148 12912 2204
rect 12848 2144 12912 2148
rect 12928 2204 12992 2208
rect 12928 2148 12932 2204
rect 12932 2148 12988 2204
rect 12988 2148 12992 2204
rect 12928 2144 12992 2148
rect 13008 2204 13072 2208
rect 13008 2148 13012 2204
rect 13012 2148 13068 2204
rect 13068 2148 13072 2204
rect 13008 2144 13072 2148
rect 13088 2204 13152 2208
rect 13088 2148 13092 2204
rect 13092 2148 13148 2204
rect 13148 2148 13152 2204
rect 13088 2144 13152 2148
rect 20778 2204 20842 2208
rect 20778 2148 20782 2204
rect 20782 2148 20838 2204
rect 20838 2148 20842 2204
rect 20778 2144 20842 2148
rect 20858 2204 20922 2208
rect 20858 2148 20862 2204
rect 20862 2148 20918 2204
rect 20918 2148 20922 2204
rect 20858 2144 20922 2148
rect 20938 2204 21002 2208
rect 20938 2148 20942 2204
rect 20942 2148 20998 2204
rect 20998 2148 21002 2204
rect 20938 2144 21002 2148
rect 21018 2204 21082 2208
rect 21018 2148 21022 2204
rect 21022 2148 21078 2204
rect 21078 2148 21082 2204
rect 21018 2144 21082 2148
rect 5396 1864 5460 1868
rect 5396 1808 5446 1864
rect 5446 1808 5460 1864
rect 5396 1804 5460 1808
<< metal4 >>
rect 4909 46816 5229 47376
rect 4909 46752 4917 46816
rect 4981 46752 4997 46816
rect 5061 46752 5077 46816
rect 5141 46752 5157 46816
rect 5221 46752 5229 46816
rect 4909 45728 5229 46752
rect 4909 45664 4917 45728
rect 4981 45664 4997 45728
rect 5061 45664 5077 45728
rect 5141 45664 5157 45728
rect 5221 45664 5229 45728
rect 4909 44640 5229 45664
rect 4909 44576 4917 44640
rect 4981 44576 4997 44640
rect 5061 44576 5077 44640
rect 5141 44576 5157 44640
rect 5221 44576 5229 44640
rect 4909 43552 5229 44576
rect 4909 43488 4917 43552
rect 4981 43488 4997 43552
rect 5061 43488 5077 43552
rect 5141 43488 5157 43552
rect 5221 43488 5229 43552
rect 4909 42464 5229 43488
rect 4909 42400 4917 42464
rect 4981 42400 4997 42464
rect 5061 42400 5077 42464
rect 5141 42400 5157 42464
rect 5221 42400 5229 42464
rect 4909 41376 5229 42400
rect 4909 41312 4917 41376
rect 4981 41312 4997 41376
rect 5061 41312 5077 41376
rect 5141 41312 5157 41376
rect 5221 41312 5229 41376
rect 4909 40288 5229 41312
rect 4909 40224 4917 40288
rect 4981 40286 4997 40288
rect 5061 40286 5077 40288
rect 5141 40286 5157 40288
rect 5221 40224 5229 40288
rect 4909 40050 4951 40224
rect 5187 40050 5229 40224
rect 4909 39200 5229 40050
rect 4909 39136 4917 39200
rect 4981 39136 4997 39200
rect 5061 39136 5077 39200
rect 5141 39136 5157 39200
rect 5221 39136 5229 39200
rect 4909 38112 5229 39136
rect 4909 38048 4917 38112
rect 4981 38048 4997 38112
rect 5061 38048 5077 38112
rect 5141 38048 5157 38112
rect 5221 38048 5229 38112
rect 4909 37024 5229 38048
rect 4909 36960 4917 37024
rect 4981 36960 4997 37024
rect 5061 36960 5077 37024
rect 5141 36960 5157 37024
rect 5221 36960 5229 37024
rect 4909 35936 5229 36960
rect 4909 35872 4917 35936
rect 4981 35872 4997 35936
rect 5061 35872 5077 35936
rect 5141 35872 5157 35936
rect 5221 35872 5229 35936
rect 4909 34848 5229 35872
rect 4909 34784 4917 34848
rect 4981 34784 4997 34848
rect 5061 34784 5077 34848
rect 5141 34784 5157 34848
rect 5221 34784 5229 34848
rect 4909 33760 5229 34784
rect 8874 47360 9194 47376
rect 8874 47296 8882 47360
rect 8946 47296 8962 47360
rect 9026 47296 9042 47360
rect 9106 47296 9122 47360
rect 9186 47296 9194 47360
rect 8874 46272 9194 47296
rect 8874 46208 8882 46272
rect 8946 46208 8962 46272
rect 9026 46208 9042 46272
rect 9106 46208 9122 46272
rect 9186 46208 9194 46272
rect 8874 45184 9194 46208
rect 8874 45120 8882 45184
rect 8946 45120 8962 45184
rect 9026 45120 9042 45184
rect 9106 45120 9122 45184
rect 9186 45120 9194 45184
rect 8874 44096 9194 45120
rect 8874 44032 8882 44096
rect 8946 44032 8962 44096
rect 9026 44032 9042 44096
rect 9106 44032 9122 44096
rect 9186 44032 9194 44096
rect 8874 43008 9194 44032
rect 8874 42944 8882 43008
rect 8946 42944 8962 43008
rect 9026 42944 9042 43008
rect 9106 42944 9122 43008
rect 9186 42944 9194 43008
rect 8874 41920 9194 42944
rect 8874 41856 8882 41920
rect 8946 41856 8962 41920
rect 9026 41856 9042 41920
rect 9106 41856 9122 41920
rect 9186 41856 9194 41920
rect 8874 40832 9194 41856
rect 8874 40768 8882 40832
rect 8946 40768 8962 40832
rect 9026 40768 9042 40832
rect 9106 40768 9122 40832
rect 9186 40768 9194 40832
rect 8874 39744 9194 40768
rect 8874 39680 8882 39744
rect 8946 39680 8962 39744
rect 9026 39680 9042 39744
rect 9106 39680 9122 39744
rect 9186 39680 9194 39744
rect 8874 38656 9194 39680
rect 8874 38592 8882 38656
rect 8946 38592 8962 38656
rect 9026 38592 9042 38656
rect 9106 38592 9122 38656
rect 9186 38592 9194 38656
rect 8874 37568 9194 38592
rect 8874 37504 8882 37568
rect 8946 37504 8962 37568
rect 9026 37504 9042 37568
rect 9106 37504 9122 37568
rect 9186 37504 9194 37568
rect 8874 36480 9194 37504
rect 8874 36416 8882 36480
rect 8946 36416 8962 36480
rect 9026 36416 9042 36480
rect 9106 36416 9122 36480
rect 9186 36416 9194 36480
rect 8874 35392 9194 36416
rect 8874 35328 8882 35392
rect 8946 35328 8962 35392
rect 9026 35328 9042 35392
rect 9106 35328 9122 35392
rect 9186 35328 9194 35392
rect 8874 34304 9194 35328
rect 8874 34240 8882 34304
rect 8946 34240 8962 34304
rect 9026 34240 9042 34304
rect 9106 34240 9122 34304
rect 9186 34240 9194 34304
rect 5395 34236 5461 34237
rect 5395 34172 5396 34236
rect 5460 34172 5461 34236
rect 5395 34171 5461 34172
rect 4909 33696 4917 33760
rect 4981 33696 4997 33760
rect 5061 33696 5077 33760
rect 5141 33696 5157 33760
rect 5221 33696 5229 33760
rect 4909 32672 5229 33696
rect 4909 32608 4917 32672
rect 4981 32608 4997 32672
rect 5061 32608 5077 32672
rect 5141 32608 5157 32672
rect 5221 32608 5229 32672
rect 4909 31584 5229 32608
rect 5398 31653 5458 34171
rect 8874 33216 9194 34240
rect 8874 33152 8882 33216
rect 8946 33152 8962 33216
rect 9026 33152 9042 33216
rect 9106 33152 9122 33216
rect 9186 33152 9194 33216
rect 8874 32678 9194 33152
rect 8874 32442 8916 32678
rect 9152 32442 9194 32678
rect 8874 32128 9194 32442
rect 8874 32064 8882 32128
rect 8946 32064 8962 32128
rect 9026 32064 9042 32128
rect 9106 32064 9122 32128
rect 9186 32064 9194 32128
rect 5395 31652 5461 31653
rect 5395 31588 5396 31652
rect 5460 31588 5461 31652
rect 5395 31587 5461 31588
rect 4909 31520 4917 31584
rect 4981 31520 4997 31584
rect 5061 31520 5077 31584
rect 5141 31520 5157 31584
rect 5221 31520 5229 31584
rect 4909 30496 5229 31520
rect 4909 30432 4917 30496
rect 4981 30432 4997 30496
rect 5061 30432 5077 30496
rect 5141 30432 5157 30496
rect 5221 30432 5229 30496
rect 4909 29408 5229 30432
rect 4909 29344 4917 29408
rect 4981 29344 4997 29408
rect 5061 29344 5077 29408
rect 5141 29344 5157 29408
rect 5221 29344 5229 29408
rect 4909 28320 5229 29344
rect 8874 31040 9194 32064
rect 8874 30976 8882 31040
rect 8946 30976 8962 31040
rect 9026 30976 9042 31040
rect 9106 30976 9122 31040
rect 9186 30976 9194 31040
rect 8874 29952 9194 30976
rect 8874 29888 8882 29952
rect 8946 29888 8962 29952
rect 9026 29888 9042 29952
rect 9106 29888 9122 29952
rect 9186 29888 9194 29952
rect 8874 28864 9194 29888
rect 8874 28800 8882 28864
rect 8946 28800 8962 28864
rect 9026 28800 9042 28864
rect 9106 28800 9122 28864
rect 9186 28800 9194 28864
rect 5395 28524 5461 28525
rect 5395 28460 5396 28524
rect 5460 28460 5461 28524
rect 5395 28459 5461 28460
rect 8339 28524 8405 28525
rect 8339 28460 8340 28524
rect 8404 28460 8405 28524
rect 8339 28459 8405 28460
rect 4909 28256 4917 28320
rect 4981 28256 4997 28320
rect 5061 28256 5077 28320
rect 5141 28256 5157 28320
rect 5221 28256 5229 28320
rect 4909 27232 5229 28256
rect 4909 27168 4917 27232
rect 4981 27168 4997 27232
rect 5061 27168 5077 27232
rect 5141 27168 5157 27232
rect 5221 27168 5229 27232
rect 4909 26144 5229 27168
rect 4909 26080 4917 26144
rect 4981 26080 4997 26144
rect 5061 26080 5077 26144
rect 5141 26080 5157 26144
rect 5221 26080 5229 26144
rect 4909 25070 5229 26080
rect 4909 25056 4951 25070
rect 5187 25056 5229 25070
rect 4909 24992 4917 25056
rect 5221 24992 5229 25056
rect 4909 24834 4951 24992
rect 5187 24834 5229 24992
rect 4909 23968 5229 24834
rect 4909 23904 4917 23968
rect 4981 23904 4997 23968
rect 5061 23904 5077 23968
rect 5141 23904 5157 23968
rect 5221 23904 5229 23968
rect 4909 22880 5229 23904
rect 5398 23085 5458 28459
rect 5395 23084 5461 23085
rect 5395 23020 5396 23084
rect 5460 23020 5461 23084
rect 5395 23019 5461 23020
rect 4909 22816 4917 22880
rect 4981 22816 4997 22880
rect 5061 22816 5077 22880
rect 5141 22816 5157 22880
rect 5221 22816 5229 22880
rect 4909 21792 5229 22816
rect 7971 22812 8037 22813
rect 7971 22748 7972 22812
rect 8036 22748 8037 22812
rect 7971 22747 8037 22748
rect 7051 21996 7117 21997
rect 7051 21932 7052 21996
rect 7116 21932 7117 21996
rect 7051 21931 7117 21932
rect 4909 21728 4917 21792
rect 4981 21728 4997 21792
rect 5061 21728 5077 21792
rect 5141 21728 5157 21792
rect 5221 21728 5229 21792
rect 4909 20704 5229 21728
rect 6867 21588 6933 21589
rect 6867 21524 6868 21588
rect 6932 21524 6933 21588
rect 6867 21523 6933 21524
rect 4909 20640 4917 20704
rect 4981 20640 4997 20704
rect 5061 20640 5077 20704
rect 5141 20640 5157 20704
rect 5221 20640 5229 20704
rect 4909 19616 5229 20640
rect 4909 19552 4917 19616
rect 4981 19552 4997 19616
rect 5061 19552 5077 19616
rect 5141 19552 5157 19616
rect 5221 19552 5229 19616
rect 4909 18528 5229 19552
rect 6870 19413 6930 21523
rect 7054 19957 7114 21931
rect 7974 21861 8034 22747
rect 8342 22541 8402 28459
rect 8874 27776 9194 28800
rect 8874 27712 8882 27776
rect 8946 27712 8962 27776
rect 9026 27712 9042 27776
rect 9106 27712 9122 27776
rect 9186 27712 9194 27776
rect 8523 27028 8589 27029
rect 8523 26964 8524 27028
rect 8588 26964 8589 27028
rect 8523 26963 8589 26964
rect 8526 24309 8586 26963
rect 8707 26756 8773 26757
rect 8707 26692 8708 26756
rect 8772 26692 8773 26756
rect 8707 26691 8773 26692
rect 8523 24308 8589 24309
rect 8523 24244 8524 24308
rect 8588 24244 8589 24308
rect 8523 24243 8589 24244
rect 8526 22677 8586 24243
rect 8523 22676 8589 22677
rect 8523 22612 8524 22676
rect 8588 22612 8589 22676
rect 8523 22611 8589 22612
rect 8339 22540 8405 22541
rect 8339 22476 8340 22540
rect 8404 22476 8405 22540
rect 8339 22475 8405 22476
rect 7971 21860 8037 21861
rect 7971 21796 7972 21860
rect 8036 21796 8037 21860
rect 7971 21795 8037 21796
rect 7419 21724 7485 21725
rect 7419 21660 7420 21724
rect 7484 21660 7485 21724
rect 7419 21659 7485 21660
rect 7051 19956 7117 19957
rect 7051 19892 7052 19956
rect 7116 19892 7117 19956
rect 7051 19891 7117 19892
rect 6867 19412 6933 19413
rect 6867 19348 6868 19412
rect 6932 19348 6933 19412
rect 6867 19347 6933 19348
rect 7422 19005 7482 21659
rect 8342 20773 8402 22475
rect 8710 21045 8770 26691
rect 8874 26688 9194 27712
rect 12840 46816 13160 47376
rect 12840 46752 12848 46816
rect 12912 46752 12928 46816
rect 12992 46752 13008 46816
rect 13072 46752 13088 46816
rect 13152 46752 13160 46816
rect 12840 45728 13160 46752
rect 12840 45664 12848 45728
rect 12912 45664 12928 45728
rect 12992 45664 13008 45728
rect 13072 45664 13088 45728
rect 13152 45664 13160 45728
rect 12840 44640 13160 45664
rect 12840 44576 12848 44640
rect 12912 44576 12928 44640
rect 12992 44576 13008 44640
rect 13072 44576 13088 44640
rect 13152 44576 13160 44640
rect 12840 43552 13160 44576
rect 12840 43488 12848 43552
rect 12912 43488 12928 43552
rect 12992 43488 13008 43552
rect 13072 43488 13088 43552
rect 13152 43488 13160 43552
rect 12840 42464 13160 43488
rect 12840 42400 12848 42464
rect 12912 42400 12928 42464
rect 12992 42400 13008 42464
rect 13072 42400 13088 42464
rect 13152 42400 13160 42464
rect 12840 41376 13160 42400
rect 12840 41312 12848 41376
rect 12912 41312 12928 41376
rect 12992 41312 13008 41376
rect 13072 41312 13088 41376
rect 13152 41312 13160 41376
rect 12840 40288 13160 41312
rect 12840 40224 12848 40288
rect 12912 40286 12928 40288
rect 12992 40286 13008 40288
rect 13072 40286 13088 40288
rect 13152 40224 13160 40288
rect 12840 40050 12882 40224
rect 13118 40050 13160 40224
rect 12840 39200 13160 40050
rect 12840 39136 12848 39200
rect 12912 39136 12928 39200
rect 12992 39136 13008 39200
rect 13072 39136 13088 39200
rect 13152 39136 13160 39200
rect 12840 38112 13160 39136
rect 12840 38048 12848 38112
rect 12912 38048 12928 38112
rect 12992 38048 13008 38112
rect 13072 38048 13088 38112
rect 13152 38048 13160 38112
rect 12840 37024 13160 38048
rect 12840 36960 12848 37024
rect 12912 36960 12928 37024
rect 12992 36960 13008 37024
rect 13072 36960 13088 37024
rect 13152 36960 13160 37024
rect 12840 35936 13160 36960
rect 12840 35872 12848 35936
rect 12912 35872 12928 35936
rect 12992 35872 13008 35936
rect 13072 35872 13088 35936
rect 13152 35872 13160 35936
rect 12840 34848 13160 35872
rect 12840 34784 12848 34848
rect 12912 34784 12928 34848
rect 12992 34784 13008 34848
rect 13072 34784 13088 34848
rect 13152 34784 13160 34848
rect 12840 33760 13160 34784
rect 12840 33696 12848 33760
rect 12912 33696 12928 33760
rect 12992 33696 13008 33760
rect 13072 33696 13088 33760
rect 13152 33696 13160 33760
rect 12840 32672 13160 33696
rect 12840 32608 12848 32672
rect 12912 32608 12928 32672
rect 12992 32608 13008 32672
rect 13072 32608 13088 32672
rect 13152 32608 13160 32672
rect 12840 31584 13160 32608
rect 12840 31520 12848 31584
rect 12912 31520 12928 31584
rect 12992 31520 13008 31584
rect 13072 31520 13088 31584
rect 13152 31520 13160 31584
rect 12840 30496 13160 31520
rect 12840 30432 12848 30496
rect 12912 30432 12928 30496
rect 12992 30432 13008 30496
rect 13072 30432 13088 30496
rect 13152 30432 13160 30496
rect 12840 29408 13160 30432
rect 12840 29344 12848 29408
rect 12912 29344 12928 29408
rect 12992 29344 13008 29408
rect 13072 29344 13088 29408
rect 13152 29344 13160 29408
rect 12840 28320 13160 29344
rect 12840 28256 12848 28320
rect 12912 28256 12928 28320
rect 12992 28256 13008 28320
rect 13072 28256 13088 28320
rect 13152 28256 13160 28320
rect 9627 27300 9693 27301
rect 9627 27236 9628 27300
rect 9692 27236 9693 27300
rect 9627 27235 9693 27236
rect 8874 26624 8882 26688
rect 8946 26624 8962 26688
rect 9026 26624 9042 26688
rect 9106 26624 9122 26688
rect 9186 26624 9194 26688
rect 8874 25600 9194 26624
rect 9443 26076 9509 26077
rect 9443 26012 9444 26076
rect 9508 26012 9509 26076
rect 9443 26011 9509 26012
rect 8874 25536 8882 25600
rect 8946 25536 8962 25600
rect 9026 25536 9042 25600
rect 9106 25536 9122 25600
rect 9186 25536 9194 25600
rect 8874 24512 9194 25536
rect 9259 24852 9325 24853
rect 9259 24788 9260 24852
rect 9324 24788 9325 24852
rect 9259 24787 9325 24788
rect 8874 24448 8882 24512
rect 8946 24448 8962 24512
rect 9026 24448 9042 24512
rect 9106 24448 9122 24512
rect 9186 24448 9194 24512
rect 8874 23424 9194 24448
rect 8874 23360 8882 23424
rect 8946 23360 8962 23424
rect 9026 23360 9042 23424
rect 9106 23360 9122 23424
rect 9186 23360 9194 23424
rect 8874 22336 9194 23360
rect 8874 22272 8882 22336
rect 8946 22272 8962 22336
rect 9026 22272 9042 22336
rect 9106 22272 9122 22336
rect 9186 22272 9194 22336
rect 8874 21248 9194 22272
rect 8874 21184 8882 21248
rect 8946 21184 8962 21248
rect 9026 21184 9042 21248
rect 9106 21184 9122 21248
rect 9186 21184 9194 21248
rect 8707 21044 8773 21045
rect 8707 20980 8708 21044
rect 8772 20980 8773 21044
rect 8707 20979 8773 20980
rect 8339 20772 8405 20773
rect 8339 20708 8340 20772
rect 8404 20708 8405 20772
rect 8339 20707 8405 20708
rect 8874 20160 9194 21184
rect 9262 20501 9322 24787
rect 9446 21997 9506 26011
rect 9443 21996 9509 21997
rect 9443 21932 9444 21996
rect 9508 21932 9509 21996
rect 9443 21931 9509 21932
rect 9259 20500 9325 20501
rect 9259 20436 9260 20500
rect 9324 20436 9325 20500
rect 9259 20435 9325 20436
rect 8874 20096 8882 20160
rect 8946 20096 8962 20160
rect 9026 20096 9042 20160
rect 9106 20096 9122 20160
rect 9186 20096 9194 20160
rect 8874 19072 9194 20096
rect 9630 19821 9690 27235
rect 12840 27232 13160 28256
rect 12840 27168 12848 27232
rect 12912 27168 12928 27232
rect 12992 27168 13008 27232
rect 13072 27168 13088 27232
rect 13152 27168 13160 27232
rect 10179 27028 10245 27029
rect 10179 26964 10180 27028
rect 10244 26964 10245 27028
rect 10179 26963 10245 26964
rect 9627 19820 9693 19821
rect 9627 19756 9628 19820
rect 9692 19756 9693 19820
rect 9627 19755 9693 19756
rect 10182 19141 10242 26963
rect 12840 26144 13160 27168
rect 12840 26080 12848 26144
rect 12912 26080 12928 26144
rect 12992 26080 13008 26144
rect 13072 26080 13088 26144
rect 13152 26080 13160 26144
rect 12840 25070 13160 26080
rect 12840 25056 12882 25070
rect 13118 25056 13160 25070
rect 12840 24992 12848 25056
rect 13152 24992 13160 25056
rect 12840 24834 12882 24992
rect 13118 24834 13160 24992
rect 12840 23968 13160 24834
rect 12840 23904 12848 23968
rect 12912 23904 12928 23968
rect 12992 23904 13008 23968
rect 13072 23904 13088 23968
rect 13152 23904 13160 23968
rect 12840 22880 13160 23904
rect 12840 22816 12848 22880
rect 12912 22816 12928 22880
rect 12992 22816 13008 22880
rect 13072 22816 13088 22880
rect 13152 22816 13160 22880
rect 12840 21792 13160 22816
rect 12840 21728 12848 21792
rect 12912 21728 12928 21792
rect 12992 21728 13008 21792
rect 13072 21728 13088 21792
rect 13152 21728 13160 21792
rect 12840 20704 13160 21728
rect 12840 20640 12848 20704
rect 12912 20640 12928 20704
rect 12992 20640 13008 20704
rect 13072 20640 13088 20704
rect 13152 20640 13160 20704
rect 12840 19616 13160 20640
rect 12840 19552 12848 19616
rect 12912 19552 12928 19616
rect 12992 19552 13008 19616
rect 13072 19552 13088 19616
rect 13152 19552 13160 19616
rect 10179 19140 10245 19141
rect 10179 19076 10180 19140
rect 10244 19076 10245 19140
rect 10179 19075 10245 19076
rect 8874 19008 8882 19072
rect 8946 19008 8962 19072
rect 9026 19008 9042 19072
rect 9106 19008 9122 19072
rect 9186 19008 9194 19072
rect 7419 19004 7485 19005
rect 7419 18940 7420 19004
rect 7484 18940 7485 19004
rect 7419 18939 7485 18940
rect 5395 18732 5461 18733
rect 5395 18668 5396 18732
rect 5460 18668 5461 18732
rect 5395 18667 5461 18668
rect 4909 18464 4917 18528
rect 4981 18464 4997 18528
rect 5061 18464 5077 18528
rect 5141 18464 5157 18528
rect 5221 18464 5229 18528
rect 4909 17440 5229 18464
rect 4909 17376 4917 17440
rect 4981 17376 4997 17440
rect 5061 17376 5077 17440
rect 5141 17376 5157 17440
rect 5221 17376 5229 17440
rect 4909 16352 5229 17376
rect 4909 16288 4917 16352
rect 4981 16288 4997 16352
rect 5061 16288 5077 16352
rect 5141 16288 5157 16352
rect 5221 16288 5229 16352
rect 4909 15264 5229 16288
rect 4909 15200 4917 15264
rect 4981 15200 4997 15264
rect 5061 15200 5077 15264
rect 5141 15200 5157 15264
rect 5221 15200 5229 15264
rect 4909 14176 5229 15200
rect 4909 14112 4917 14176
rect 4981 14112 4997 14176
rect 5061 14112 5077 14176
rect 5141 14112 5157 14176
rect 5221 14112 5229 14176
rect 4909 13088 5229 14112
rect 4909 13024 4917 13088
rect 4981 13024 4997 13088
rect 5061 13024 5077 13088
rect 5141 13024 5157 13088
rect 5221 13024 5229 13088
rect 4909 12000 5229 13024
rect 5398 12885 5458 18667
rect 8874 17984 9194 19008
rect 8874 17920 8882 17984
rect 8946 17920 8962 17984
rect 9026 17920 9042 17984
rect 9106 17920 9122 17984
rect 9186 17920 9194 17984
rect 8874 17462 9194 17920
rect 8874 17226 8916 17462
rect 9152 17226 9194 17462
rect 8874 16896 9194 17226
rect 8874 16832 8882 16896
rect 8946 16832 8962 16896
rect 9026 16832 9042 16896
rect 9106 16832 9122 16896
rect 9186 16832 9194 16896
rect 8874 15808 9194 16832
rect 8874 15744 8882 15808
rect 8946 15744 8962 15808
rect 9026 15744 9042 15808
rect 9106 15744 9122 15808
rect 9186 15744 9194 15808
rect 8874 14720 9194 15744
rect 8874 14656 8882 14720
rect 8946 14656 8962 14720
rect 9026 14656 9042 14720
rect 9106 14656 9122 14720
rect 9186 14656 9194 14720
rect 8874 13632 9194 14656
rect 8874 13568 8882 13632
rect 8946 13568 8962 13632
rect 9026 13568 9042 13632
rect 9106 13568 9122 13632
rect 9186 13568 9194 13632
rect 5395 12884 5461 12885
rect 5395 12820 5396 12884
rect 5460 12820 5461 12884
rect 5395 12819 5461 12820
rect 4909 11936 4917 12000
rect 4981 11936 4997 12000
rect 5061 11936 5077 12000
rect 5141 11936 5157 12000
rect 5221 11936 5229 12000
rect 4909 10912 5229 11936
rect 4909 10848 4917 10912
rect 4981 10848 4997 10912
rect 5061 10848 5077 10912
rect 5141 10848 5157 10912
rect 5221 10848 5229 10912
rect 4909 9854 5229 10848
rect 8874 12544 9194 13568
rect 12840 18528 13160 19552
rect 12840 18464 12848 18528
rect 12912 18464 12928 18528
rect 12992 18464 13008 18528
rect 13072 18464 13088 18528
rect 13152 18464 13160 18528
rect 12840 17440 13160 18464
rect 12840 17376 12848 17440
rect 12912 17376 12928 17440
rect 12992 17376 13008 17440
rect 13072 17376 13088 17440
rect 13152 17376 13160 17440
rect 12840 16352 13160 17376
rect 12840 16288 12848 16352
rect 12912 16288 12928 16352
rect 12992 16288 13008 16352
rect 13072 16288 13088 16352
rect 13152 16288 13160 16352
rect 12840 15264 13160 16288
rect 12840 15200 12848 15264
rect 12912 15200 12928 15264
rect 12992 15200 13008 15264
rect 13072 15200 13088 15264
rect 13152 15200 13160 15264
rect 12840 14176 13160 15200
rect 12840 14112 12848 14176
rect 12912 14112 12928 14176
rect 12992 14112 13008 14176
rect 13072 14112 13088 14176
rect 13152 14112 13160 14176
rect 9443 13156 9509 13157
rect 9443 13092 9444 13156
rect 9508 13092 9509 13156
rect 9443 13091 9509 13092
rect 8874 12480 8882 12544
rect 8946 12480 8962 12544
rect 9026 12480 9042 12544
rect 9106 12480 9122 12544
rect 9186 12480 9194 12544
rect 8874 11456 9194 12480
rect 8874 11392 8882 11456
rect 8946 11392 8962 11456
rect 9026 11392 9042 11456
rect 9106 11392 9122 11456
rect 9186 11392 9194 11456
rect 8874 10368 9194 11392
rect 8874 10304 8882 10368
rect 8946 10304 8962 10368
rect 9026 10304 9042 10368
rect 9106 10304 9122 10368
rect 9186 10304 9194 10368
rect 7235 10300 7301 10301
rect 7235 10236 7236 10300
rect 7300 10236 7301 10300
rect 7235 10235 7301 10236
rect 4909 9824 4951 9854
rect 5187 9824 5229 9854
rect 4909 9760 4917 9824
rect 5221 9760 5229 9824
rect 4909 9618 4951 9760
rect 5187 9618 5229 9760
rect 4909 8736 5229 9618
rect 5395 9076 5461 9077
rect 5395 9012 5396 9076
rect 5460 9012 5461 9076
rect 5395 9011 5461 9012
rect 4909 8672 4917 8736
rect 4981 8672 4997 8736
rect 5061 8672 5077 8736
rect 5141 8672 5157 8736
rect 5221 8672 5229 8736
rect 4909 7648 5229 8672
rect 4909 7584 4917 7648
rect 4981 7584 4997 7648
rect 5061 7584 5077 7648
rect 5141 7584 5157 7648
rect 5221 7584 5229 7648
rect 4909 6560 5229 7584
rect 4909 6496 4917 6560
rect 4981 6496 4997 6560
rect 5061 6496 5077 6560
rect 5141 6496 5157 6560
rect 5221 6496 5229 6560
rect 4909 5472 5229 6496
rect 4909 5408 4917 5472
rect 4981 5408 4997 5472
rect 5061 5408 5077 5472
rect 5141 5408 5157 5472
rect 5221 5408 5229 5472
rect 4909 4384 5229 5408
rect 4909 4320 4917 4384
rect 4981 4320 4997 4384
rect 5061 4320 5077 4384
rect 5141 4320 5157 4384
rect 5221 4320 5229 4384
rect 4909 3296 5229 4320
rect 4909 3232 4917 3296
rect 4981 3232 4997 3296
rect 5061 3232 5077 3296
rect 5141 3232 5157 3296
rect 5221 3232 5229 3296
rect 4909 2208 5229 3232
rect 4909 2144 4917 2208
rect 4981 2144 4997 2208
rect 5061 2144 5077 2208
rect 5141 2144 5157 2208
rect 5221 2144 5229 2208
rect 4909 2128 5229 2144
rect 5398 1869 5458 9011
rect 7238 7853 7298 10235
rect 8874 9280 9194 10304
rect 8874 9216 8882 9280
rect 8946 9216 8962 9280
rect 9026 9216 9042 9280
rect 9106 9216 9122 9280
rect 9186 9216 9194 9280
rect 8874 8192 9194 9216
rect 8874 8128 8882 8192
rect 8946 8128 8962 8192
rect 9026 8128 9042 8192
rect 9106 8128 9122 8192
rect 9186 8128 9194 8192
rect 7235 7852 7301 7853
rect 7235 7788 7236 7852
rect 7300 7788 7301 7852
rect 7235 7787 7301 7788
rect 8874 7104 9194 8128
rect 8874 7040 8882 7104
rect 8946 7040 8962 7104
rect 9026 7040 9042 7104
rect 9106 7040 9122 7104
rect 9186 7040 9194 7104
rect 8874 6016 9194 7040
rect 8874 5952 8882 6016
rect 8946 5952 8962 6016
rect 9026 5952 9042 6016
rect 9106 5952 9122 6016
rect 9186 5952 9194 6016
rect 8874 4928 9194 5952
rect 8874 4864 8882 4928
rect 8946 4864 8962 4928
rect 9026 4864 9042 4928
rect 9106 4864 9122 4928
rect 9186 4864 9194 4928
rect 8874 3840 9194 4864
rect 8874 3776 8882 3840
rect 8946 3776 8962 3840
rect 9026 3776 9042 3840
rect 9106 3776 9122 3840
rect 9186 3776 9194 3840
rect 8874 2752 9194 3776
rect 9446 3229 9506 13091
rect 12840 13088 13160 14112
rect 12840 13024 12848 13088
rect 12912 13024 12928 13088
rect 12992 13024 13008 13088
rect 13072 13024 13088 13088
rect 13152 13024 13160 13088
rect 12840 12000 13160 13024
rect 12840 11936 12848 12000
rect 12912 11936 12928 12000
rect 12992 11936 13008 12000
rect 13072 11936 13088 12000
rect 13152 11936 13160 12000
rect 12840 10912 13160 11936
rect 12840 10848 12848 10912
rect 12912 10848 12928 10912
rect 12992 10848 13008 10912
rect 13072 10848 13088 10912
rect 13152 10848 13160 10912
rect 12203 9892 12269 9893
rect 12203 9828 12204 9892
rect 12268 9828 12269 9892
rect 12203 9827 12269 9828
rect 12840 9854 13160 10848
rect 12206 4453 12266 9827
rect 12840 9824 12882 9854
rect 13118 9824 13160 9854
rect 12840 9760 12848 9824
rect 13152 9760 13160 9824
rect 12840 9618 12882 9760
rect 13118 9618 13160 9760
rect 12571 9076 12637 9077
rect 12571 9012 12572 9076
rect 12636 9012 12637 9076
rect 12571 9011 12637 9012
rect 12574 8533 12634 9011
rect 12840 8736 13160 9618
rect 16805 47360 17125 47376
rect 16805 47296 16813 47360
rect 16877 47296 16893 47360
rect 16957 47296 16973 47360
rect 17037 47296 17053 47360
rect 17117 47296 17125 47360
rect 16805 46272 17125 47296
rect 16805 46208 16813 46272
rect 16877 46208 16893 46272
rect 16957 46208 16973 46272
rect 17037 46208 17053 46272
rect 17117 46208 17125 46272
rect 16805 45184 17125 46208
rect 16805 45120 16813 45184
rect 16877 45120 16893 45184
rect 16957 45120 16973 45184
rect 17037 45120 17053 45184
rect 17117 45120 17125 45184
rect 16805 44096 17125 45120
rect 16805 44032 16813 44096
rect 16877 44032 16893 44096
rect 16957 44032 16973 44096
rect 17037 44032 17053 44096
rect 17117 44032 17125 44096
rect 16805 43008 17125 44032
rect 16805 42944 16813 43008
rect 16877 42944 16893 43008
rect 16957 42944 16973 43008
rect 17037 42944 17053 43008
rect 17117 42944 17125 43008
rect 16805 41920 17125 42944
rect 16805 41856 16813 41920
rect 16877 41856 16893 41920
rect 16957 41856 16973 41920
rect 17037 41856 17053 41920
rect 17117 41856 17125 41920
rect 16805 40832 17125 41856
rect 16805 40768 16813 40832
rect 16877 40768 16893 40832
rect 16957 40768 16973 40832
rect 17037 40768 17053 40832
rect 17117 40768 17125 40832
rect 16805 39744 17125 40768
rect 16805 39680 16813 39744
rect 16877 39680 16893 39744
rect 16957 39680 16973 39744
rect 17037 39680 17053 39744
rect 17117 39680 17125 39744
rect 16805 38656 17125 39680
rect 16805 38592 16813 38656
rect 16877 38592 16893 38656
rect 16957 38592 16973 38656
rect 17037 38592 17053 38656
rect 17117 38592 17125 38656
rect 16805 37568 17125 38592
rect 16805 37504 16813 37568
rect 16877 37504 16893 37568
rect 16957 37504 16973 37568
rect 17037 37504 17053 37568
rect 17117 37504 17125 37568
rect 16805 36480 17125 37504
rect 16805 36416 16813 36480
rect 16877 36416 16893 36480
rect 16957 36416 16973 36480
rect 17037 36416 17053 36480
rect 17117 36416 17125 36480
rect 16805 35392 17125 36416
rect 16805 35328 16813 35392
rect 16877 35328 16893 35392
rect 16957 35328 16973 35392
rect 17037 35328 17053 35392
rect 17117 35328 17125 35392
rect 16805 34304 17125 35328
rect 16805 34240 16813 34304
rect 16877 34240 16893 34304
rect 16957 34240 16973 34304
rect 17037 34240 17053 34304
rect 17117 34240 17125 34304
rect 16805 33216 17125 34240
rect 16805 33152 16813 33216
rect 16877 33152 16893 33216
rect 16957 33152 16973 33216
rect 17037 33152 17053 33216
rect 17117 33152 17125 33216
rect 16805 32678 17125 33152
rect 16805 32442 16847 32678
rect 17083 32442 17125 32678
rect 16805 32128 17125 32442
rect 16805 32064 16813 32128
rect 16877 32064 16893 32128
rect 16957 32064 16973 32128
rect 17037 32064 17053 32128
rect 17117 32064 17125 32128
rect 16805 31040 17125 32064
rect 16805 30976 16813 31040
rect 16877 30976 16893 31040
rect 16957 30976 16973 31040
rect 17037 30976 17053 31040
rect 17117 30976 17125 31040
rect 16805 29952 17125 30976
rect 16805 29888 16813 29952
rect 16877 29888 16893 29952
rect 16957 29888 16973 29952
rect 17037 29888 17053 29952
rect 17117 29888 17125 29952
rect 16805 28864 17125 29888
rect 16805 28800 16813 28864
rect 16877 28800 16893 28864
rect 16957 28800 16973 28864
rect 17037 28800 17053 28864
rect 17117 28800 17125 28864
rect 16805 27776 17125 28800
rect 16805 27712 16813 27776
rect 16877 27712 16893 27776
rect 16957 27712 16973 27776
rect 17037 27712 17053 27776
rect 17117 27712 17125 27776
rect 16805 26688 17125 27712
rect 16805 26624 16813 26688
rect 16877 26624 16893 26688
rect 16957 26624 16973 26688
rect 17037 26624 17053 26688
rect 17117 26624 17125 26688
rect 16805 25600 17125 26624
rect 16805 25536 16813 25600
rect 16877 25536 16893 25600
rect 16957 25536 16973 25600
rect 17037 25536 17053 25600
rect 17117 25536 17125 25600
rect 16805 24512 17125 25536
rect 16805 24448 16813 24512
rect 16877 24448 16893 24512
rect 16957 24448 16973 24512
rect 17037 24448 17053 24512
rect 17117 24448 17125 24512
rect 16805 23424 17125 24448
rect 16805 23360 16813 23424
rect 16877 23360 16893 23424
rect 16957 23360 16973 23424
rect 17037 23360 17053 23424
rect 17117 23360 17125 23424
rect 16805 22336 17125 23360
rect 16805 22272 16813 22336
rect 16877 22272 16893 22336
rect 16957 22272 16973 22336
rect 17037 22272 17053 22336
rect 17117 22272 17125 22336
rect 16805 21248 17125 22272
rect 16805 21184 16813 21248
rect 16877 21184 16893 21248
rect 16957 21184 16973 21248
rect 17037 21184 17053 21248
rect 17117 21184 17125 21248
rect 16805 20160 17125 21184
rect 16805 20096 16813 20160
rect 16877 20096 16893 20160
rect 16957 20096 16973 20160
rect 17037 20096 17053 20160
rect 17117 20096 17125 20160
rect 16805 19072 17125 20096
rect 16805 19008 16813 19072
rect 16877 19008 16893 19072
rect 16957 19008 16973 19072
rect 17037 19008 17053 19072
rect 17117 19008 17125 19072
rect 16805 17984 17125 19008
rect 16805 17920 16813 17984
rect 16877 17920 16893 17984
rect 16957 17920 16973 17984
rect 17037 17920 17053 17984
rect 17117 17920 17125 17984
rect 16805 17462 17125 17920
rect 16805 17226 16847 17462
rect 17083 17226 17125 17462
rect 16805 16896 17125 17226
rect 16805 16832 16813 16896
rect 16877 16832 16893 16896
rect 16957 16832 16973 16896
rect 17037 16832 17053 16896
rect 17117 16832 17125 16896
rect 16805 15808 17125 16832
rect 16805 15744 16813 15808
rect 16877 15744 16893 15808
rect 16957 15744 16973 15808
rect 17037 15744 17053 15808
rect 17117 15744 17125 15808
rect 16805 14720 17125 15744
rect 16805 14656 16813 14720
rect 16877 14656 16893 14720
rect 16957 14656 16973 14720
rect 17037 14656 17053 14720
rect 17117 14656 17125 14720
rect 16805 13632 17125 14656
rect 16805 13568 16813 13632
rect 16877 13568 16893 13632
rect 16957 13568 16973 13632
rect 17037 13568 17053 13632
rect 17117 13568 17125 13632
rect 16805 12544 17125 13568
rect 16805 12480 16813 12544
rect 16877 12480 16893 12544
rect 16957 12480 16973 12544
rect 17037 12480 17053 12544
rect 17117 12480 17125 12544
rect 16805 11456 17125 12480
rect 16805 11392 16813 11456
rect 16877 11392 16893 11456
rect 16957 11392 16973 11456
rect 17037 11392 17053 11456
rect 17117 11392 17125 11456
rect 16805 10368 17125 11392
rect 16805 10304 16813 10368
rect 16877 10304 16893 10368
rect 16957 10304 16973 10368
rect 17037 10304 17053 10368
rect 17117 10304 17125 10368
rect 13307 9348 13373 9349
rect 13307 9284 13308 9348
rect 13372 9284 13373 9348
rect 13307 9283 13373 9284
rect 12840 8672 12848 8736
rect 12912 8672 12928 8736
rect 12992 8672 13008 8736
rect 13072 8672 13088 8736
rect 13152 8672 13160 8736
rect 12571 8532 12637 8533
rect 12571 8468 12572 8532
rect 12636 8468 12637 8532
rect 12571 8467 12637 8468
rect 12840 7648 13160 8672
rect 13310 8397 13370 9283
rect 16805 9280 17125 10304
rect 16805 9216 16813 9280
rect 16877 9216 16893 9280
rect 16957 9216 16973 9280
rect 17037 9216 17053 9280
rect 17117 9216 17125 9280
rect 13307 8396 13373 8397
rect 13307 8332 13308 8396
rect 13372 8332 13373 8396
rect 13307 8331 13373 8332
rect 13491 8260 13557 8261
rect 13491 8196 13492 8260
rect 13556 8196 13557 8260
rect 13491 8195 13557 8196
rect 12840 7584 12848 7648
rect 12912 7584 12928 7648
rect 12992 7584 13008 7648
rect 13072 7584 13088 7648
rect 13152 7584 13160 7648
rect 12840 6560 13160 7584
rect 12840 6496 12848 6560
rect 12912 6496 12928 6560
rect 12992 6496 13008 6560
rect 13072 6496 13088 6560
rect 13152 6496 13160 6560
rect 12840 5472 13160 6496
rect 12840 5408 12848 5472
rect 12912 5408 12928 5472
rect 12992 5408 13008 5472
rect 13072 5408 13088 5472
rect 13152 5408 13160 5472
rect 12203 4452 12269 4453
rect 12203 4388 12204 4452
rect 12268 4388 12269 4452
rect 12203 4387 12269 4388
rect 12840 4384 13160 5408
rect 12840 4320 12848 4384
rect 12912 4320 12928 4384
rect 12992 4320 13008 4384
rect 13072 4320 13088 4384
rect 13152 4320 13160 4384
rect 12840 3296 13160 4320
rect 13494 4181 13554 8195
rect 16805 8192 17125 9216
rect 16805 8128 16813 8192
rect 16877 8128 16893 8192
rect 16957 8128 16973 8192
rect 17037 8128 17053 8192
rect 17117 8128 17125 8192
rect 16805 7104 17125 8128
rect 16805 7040 16813 7104
rect 16877 7040 16893 7104
rect 16957 7040 16973 7104
rect 17037 7040 17053 7104
rect 17117 7040 17125 7104
rect 16805 6016 17125 7040
rect 16805 5952 16813 6016
rect 16877 5952 16893 6016
rect 16957 5952 16973 6016
rect 17037 5952 17053 6016
rect 17117 5952 17125 6016
rect 16805 4928 17125 5952
rect 16805 4864 16813 4928
rect 16877 4864 16893 4928
rect 16957 4864 16973 4928
rect 17037 4864 17053 4928
rect 17117 4864 17125 4928
rect 13491 4180 13557 4181
rect 13491 4116 13492 4180
rect 13556 4116 13557 4180
rect 13491 4115 13557 4116
rect 12840 3232 12848 3296
rect 12912 3232 12928 3296
rect 12992 3232 13008 3296
rect 13072 3232 13088 3296
rect 13152 3232 13160 3296
rect 9443 3228 9509 3229
rect 9443 3164 9444 3228
rect 9508 3164 9509 3228
rect 9443 3163 9509 3164
rect 8874 2688 8882 2752
rect 8946 2688 8962 2752
rect 9026 2688 9042 2752
rect 9106 2688 9122 2752
rect 9186 2688 9194 2752
rect 8874 2128 9194 2688
rect 12840 2208 13160 3232
rect 12840 2144 12848 2208
rect 12912 2144 12928 2208
rect 12992 2144 13008 2208
rect 13072 2144 13088 2208
rect 13152 2144 13160 2208
rect 12840 2128 13160 2144
rect 16805 3840 17125 4864
rect 16805 3776 16813 3840
rect 16877 3776 16893 3840
rect 16957 3776 16973 3840
rect 17037 3776 17053 3840
rect 17117 3776 17125 3840
rect 16805 2752 17125 3776
rect 16805 2688 16813 2752
rect 16877 2688 16893 2752
rect 16957 2688 16973 2752
rect 17037 2688 17053 2752
rect 17117 2688 17125 2752
rect 16805 2128 17125 2688
rect 20770 46816 21090 47376
rect 20770 46752 20778 46816
rect 20842 46752 20858 46816
rect 20922 46752 20938 46816
rect 21002 46752 21018 46816
rect 21082 46752 21090 46816
rect 20770 45728 21090 46752
rect 20770 45664 20778 45728
rect 20842 45664 20858 45728
rect 20922 45664 20938 45728
rect 21002 45664 21018 45728
rect 21082 45664 21090 45728
rect 20770 44640 21090 45664
rect 20770 44576 20778 44640
rect 20842 44576 20858 44640
rect 20922 44576 20938 44640
rect 21002 44576 21018 44640
rect 21082 44576 21090 44640
rect 20770 43552 21090 44576
rect 20770 43488 20778 43552
rect 20842 43488 20858 43552
rect 20922 43488 20938 43552
rect 21002 43488 21018 43552
rect 21082 43488 21090 43552
rect 20770 42464 21090 43488
rect 20770 42400 20778 42464
rect 20842 42400 20858 42464
rect 20922 42400 20938 42464
rect 21002 42400 21018 42464
rect 21082 42400 21090 42464
rect 20770 41376 21090 42400
rect 20770 41312 20778 41376
rect 20842 41312 20858 41376
rect 20922 41312 20938 41376
rect 21002 41312 21018 41376
rect 21082 41312 21090 41376
rect 20770 40288 21090 41312
rect 20770 40224 20778 40288
rect 20842 40286 20858 40288
rect 20922 40286 20938 40288
rect 21002 40286 21018 40288
rect 21082 40224 21090 40288
rect 20770 40050 20812 40224
rect 21048 40050 21090 40224
rect 20770 39200 21090 40050
rect 20770 39136 20778 39200
rect 20842 39136 20858 39200
rect 20922 39136 20938 39200
rect 21002 39136 21018 39200
rect 21082 39136 21090 39200
rect 20770 38112 21090 39136
rect 20770 38048 20778 38112
rect 20842 38048 20858 38112
rect 20922 38048 20938 38112
rect 21002 38048 21018 38112
rect 21082 38048 21090 38112
rect 20770 37024 21090 38048
rect 20770 36960 20778 37024
rect 20842 36960 20858 37024
rect 20922 36960 20938 37024
rect 21002 36960 21018 37024
rect 21082 36960 21090 37024
rect 20770 35936 21090 36960
rect 20770 35872 20778 35936
rect 20842 35872 20858 35936
rect 20922 35872 20938 35936
rect 21002 35872 21018 35936
rect 21082 35872 21090 35936
rect 20770 34848 21090 35872
rect 20770 34784 20778 34848
rect 20842 34784 20858 34848
rect 20922 34784 20938 34848
rect 21002 34784 21018 34848
rect 21082 34784 21090 34848
rect 20770 33760 21090 34784
rect 20770 33696 20778 33760
rect 20842 33696 20858 33760
rect 20922 33696 20938 33760
rect 21002 33696 21018 33760
rect 21082 33696 21090 33760
rect 20770 32672 21090 33696
rect 20770 32608 20778 32672
rect 20842 32608 20858 32672
rect 20922 32608 20938 32672
rect 21002 32608 21018 32672
rect 21082 32608 21090 32672
rect 20770 31584 21090 32608
rect 20770 31520 20778 31584
rect 20842 31520 20858 31584
rect 20922 31520 20938 31584
rect 21002 31520 21018 31584
rect 21082 31520 21090 31584
rect 20770 30496 21090 31520
rect 20770 30432 20778 30496
rect 20842 30432 20858 30496
rect 20922 30432 20938 30496
rect 21002 30432 21018 30496
rect 21082 30432 21090 30496
rect 20770 29408 21090 30432
rect 20770 29344 20778 29408
rect 20842 29344 20858 29408
rect 20922 29344 20938 29408
rect 21002 29344 21018 29408
rect 21082 29344 21090 29408
rect 20770 28320 21090 29344
rect 20770 28256 20778 28320
rect 20842 28256 20858 28320
rect 20922 28256 20938 28320
rect 21002 28256 21018 28320
rect 21082 28256 21090 28320
rect 20770 27232 21090 28256
rect 20770 27168 20778 27232
rect 20842 27168 20858 27232
rect 20922 27168 20938 27232
rect 21002 27168 21018 27232
rect 21082 27168 21090 27232
rect 20770 26144 21090 27168
rect 20770 26080 20778 26144
rect 20842 26080 20858 26144
rect 20922 26080 20938 26144
rect 21002 26080 21018 26144
rect 21082 26080 21090 26144
rect 20770 25070 21090 26080
rect 20770 25056 20812 25070
rect 21048 25056 21090 25070
rect 20770 24992 20778 25056
rect 21082 24992 21090 25056
rect 20770 24834 20812 24992
rect 21048 24834 21090 24992
rect 20770 23968 21090 24834
rect 20770 23904 20778 23968
rect 20842 23904 20858 23968
rect 20922 23904 20938 23968
rect 21002 23904 21018 23968
rect 21082 23904 21090 23968
rect 20770 22880 21090 23904
rect 20770 22816 20778 22880
rect 20842 22816 20858 22880
rect 20922 22816 20938 22880
rect 21002 22816 21018 22880
rect 21082 22816 21090 22880
rect 20770 21792 21090 22816
rect 20770 21728 20778 21792
rect 20842 21728 20858 21792
rect 20922 21728 20938 21792
rect 21002 21728 21018 21792
rect 21082 21728 21090 21792
rect 20770 20704 21090 21728
rect 20770 20640 20778 20704
rect 20842 20640 20858 20704
rect 20922 20640 20938 20704
rect 21002 20640 21018 20704
rect 21082 20640 21090 20704
rect 20770 19616 21090 20640
rect 20770 19552 20778 19616
rect 20842 19552 20858 19616
rect 20922 19552 20938 19616
rect 21002 19552 21018 19616
rect 21082 19552 21090 19616
rect 20770 18528 21090 19552
rect 20770 18464 20778 18528
rect 20842 18464 20858 18528
rect 20922 18464 20938 18528
rect 21002 18464 21018 18528
rect 21082 18464 21090 18528
rect 20770 17440 21090 18464
rect 20770 17376 20778 17440
rect 20842 17376 20858 17440
rect 20922 17376 20938 17440
rect 21002 17376 21018 17440
rect 21082 17376 21090 17440
rect 20770 16352 21090 17376
rect 20770 16288 20778 16352
rect 20842 16288 20858 16352
rect 20922 16288 20938 16352
rect 21002 16288 21018 16352
rect 21082 16288 21090 16352
rect 20770 15264 21090 16288
rect 20770 15200 20778 15264
rect 20842 15200 20858 15264
rect 20922 15200 20938 15264
rect 21002 15200 21018 15264
rect 21082 15200 21090 15264
rect 20770 14176 21090 15200
rect 20770 14112 20778 14176
rect 20842 14112 20858 14176
rect 20922 14112 20938 14176
rect 21002 14112 21018 14176
rect 21082 14112 21090 14176
rect 20770 13088 21090 14112
rect 20770 13024 20778 13088
rect 20842 13024 20858 13088
rect 20922 13024 20938 13088
rect 21002 13024 21018 13088
rect 21082 13024 21090 13088
rect 20770 12000 21090 13024
rect 20770 11936 20778 12000
rect 20842 11936 20858 12000
rect 20922 11936 20938 12000
rect 21002 11936 21018 12000
rect 21082 11936 21090 12000
rect 20770 10912 21090 11936
rect 20770 10848 20778 10912
rect 20842 10848 20858 10912
rect 20922 10848 20938 10912
rect 21002 10848 21018 10912
rect 21082 10848 21090 10912
rect 20770 9854 21090 10848
rect 20770 9824 20812 9854
rect 21048 9824 21090 9854
rect 20770 9760 20778 9824
rect 21082 9760 21090 9824
rect 20770 9618 20812 9760
rect 21048 9618 21090 9760
rect 20770 8736 21090 9618
rect 20770 8672 20778 8736
rect 20842 8672 20858 8736
rect 20922 8672 20938 8736
rect 21002 8672 21018 8736
rect 21082 8672 21090 8736
rect 20770 7648 21090 8672
rect 20770 7584 20778 7648
rect 20842 7584 20858 7648
rect 20922 7584 20938 7648
rect 21002 7584 21018 7648
rect 21082 7584 21090 7648
rect 20770 6560 21090 7584
rect 20770 6496 20778 6560
rect 20842 6496 20858 6560
rect 20922 6496 20938 6560
rect 21002 6496 21018 6560
rect 21082 6496 21090 6560
rect 20770 5472 21090 6496
rect 20770 5408 20778 5472
rect 20842 5408 20858 5472
rect 20922 5408 20938 5472
rect 21002 5408 21018 5472
rect 21082 5408 21090 5472
rect 20770 4384 21090 5408
rect 20770 4320 20778 4384
rect 20842 4320 20858 4384
rect 20922 4320 20938 4384
rect 21002 4320 21018 4384
rect 21082 4320 21090 4384
rect 20770 3296 21090 4320
rect 20770 3232 20778 3296
rect 20842 3232 20858 3296
rect 20922 3232 20938 3296
rect 21002 3232 21018 3296
rect 21082 3232 21090 3296
rect 20770 2208 21090 3232
rect 20770 2144 20778 2208
rect 20842 2144 20858 2208
rect 20922 2144 20938 2208
rect 21002 2144 21018 2208
rect 21082 2144 21090 2208
rect 20770 2128 21090 2144
rect 5395 1868 5461 1869
rect 5395 1804 5396 1868
rect 5460 1804 5461 1868
rect 5395 1803 5461 1804
<< via4 >>
rect 4951 40224 4981 40286
rect 4981 40224 4997 40286
rect 4997 40224 5061 40286
rect 5061 40224 5077 40286
rect 5077 40224 5141 40286
rect 5141 40224 5157 40286
rect 5157 40224 5187 40286
rect 4951 40050 5187 40224
rect 8916 32442 9152 32678
rect 4951 25056 5187 25070
rect 4951 24992 4981 25056
rect 4981 24992 4997 25056
rect 4997 24992 5061 25056
rect 5061 24992 5077 25056
rect 5077 24992 5141 25056
rect 5141 24992 5157 25056
rect 5157 24992 5187 25056
rect 4951 24834 5187 24992
rect 12882 40224 12912 40286
rect 12912 40224 12928 40286
rect 12928 40224 12992 40286
rect 12992 40224 13008 40286
rect 13008 40224 13072 40286
rect 13072 40224 13088 40286
rect 13088 40224 13118 40286
rect 12882 40050 13118 40224
rect 12882 25056 13118 25070
rect 12882 24992 12912 25056
rect 12912 24992 12928 25056
rect 12928 24992 12992 25056
rect 12992 24992 13008 25056
rect 13008 24992 13072 25056
rect 13072 24992 13088 25056
rect 13088 24992 13118 25056
rect 12882 24834 13118 24992
rect 8916 17226 9152 17462
rect 4951 9824 5187 9854
rect 4951 9760 4981 9824
rect 4981 9760 4997 9824
rect 4997 9760 5061 9824
rect 5061 9760 5077 9824
rect 5077 9760 5141 9824
rect 5141 9760 5157 9824
rect 5157 9760 5187 9824
rect 4951 9618 5187 9760
rect 12882 9824 13118 9854
rect 12882 9760 12912 9824
rect 12912 9760 12928 9824
rect 12928 9760 12992 9824
rect 12992 9760 13008 9824
rect 13008 9760 13072 9824
rect 13072 9760 13088 9824
rect 13088 9760 13118 9824
rect 12882 9618 13118 9760
rect 16847 32442 17083 32678
rect 16847 17226 17083 17462
rect 20812 40224 20842 40286
rect 20842 40224 20858 40286
rect 20858 40224 20922 40286
rect 20922 40224 20938 40286
rect 20938 40224 21002 40286
rect 21002 40224 21018 40286
rect 21018 40224 21048 40286
rect 20812 40050 21048 40224
rect 20812 25056 21048 25070
rect 20812 24992 20842 25056
rect 20842 24992 20858 25056
rect 20858 24992 20922 25056
rect 20922 24992 20938 25056
rect 20938 24992 21002 25056
rect 21002 24992 21018 25056
rect 21018 24992 21048 25056
rect 20812 24834 21048 24992
rect 20812 9824 21048 9854
rect 20812 9760 20842 9824
rect 20842 9760 20858 9824
rect 20858 9760 20922 9824
rect 20922 9760 20938 9824
rect 20938 9760 21002 9824
rect 21002 9760 21018 9824
rect 21018 9760 21048 9824
rect 20812 9618 21048 9760
<< metal5 >>
rect 1104 40286 24840 40328
rect 1104 40050 4951 40286
rect 5187 40050 12882 40286
rect 13118 40050 20812 40286
rect 21048 40050 24840 40286
rect 1104 40008 24840 40050
rect 1104 32678 24840 32720
rect 1104 32442 8916 32678
rect 9152 32442 16847 32678
rect 17083 32442 24840 32678
rect 1104 32400 24840 32442
rect 1104 25070 24840 25112
rect 1104 24834 4951 25070
rect 5187 24834 12882 25070
rect 13118 24834 20812 25070
rect 21048 24834 24840 25070
rect 1104 24792 24840 24834
rect 1104 17462 24840 17504
rect 1104 17226 8916 17462
rect 9152 17226 16847 17462
rect 17083 17226 24840 17462
rect 1104 17184 24840 17226
rect 1104 9854 24840 9896
rect 1104 9618 4951 9854
rect 5187 9618 12882 9854
rect 13118 9618 20812 9854
rect 21048 9618 24840 9854
rect 1104 9576 24840 9618
use sky130_fd_sc_hd__decap_8  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1748 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7
timestamp 1607721120
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607721120
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1840 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0817_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1472 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2668 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2668 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_36
timestamp 1607721120
transform 1 0 4416 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1607721120
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1607721120
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 4232 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1607721120
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1607721120
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43
timestamp 1607721120
transform 1 0 5060 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607721120
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607721120
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0609_
timestamp 1607721120
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1607721120
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1607721120
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79
timestamp 1607721120
transform 1 0 8372 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1258_
timestamp 1607721120
transform 1 0 7452 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6900 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_1_99
timestamp 1607721120
transform 1 0 10212 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_88
timestamp 1607721120
transform 1 0 9200 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1607721120
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1607721120
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607721120
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607721120
transform 1 0 9844 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1607721120
transform 1 0 9936 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1607721120
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1607721120
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114
timestamp 1607721120
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607721120
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607721120
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607721120
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1607721120
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1607721120
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_142
timestamp 1607721120
transform 1 0 14168 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_136
timestamp 1607721120
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128
timestamp 1607721120
transform 1 0 12880 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1020_
timestamp 1607721120
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607721120
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_159
timestamp 1607721120
transform 1 0 15732 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1607721120
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607721120
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1607721120
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0606_
timestamp 1607721120
transform 1 0 14904 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_184
timestamp 1607721120
transform 1 0 18032 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607721120
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_183
timestamp 1607721120
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_171
timestamp 1607721120
transform 1 0 16836 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607721120
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607721120
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0822_
timestamp 1607721120
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204
timestamp 1607721120
transform 1 0 19872 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_192
timestamp 1607721120
transform 1 0 18768 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_208
timestamp 1607721120
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_196
timestamp 1607721120
transform 1 0 19136 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0820_
timestamp 1607721120
transform 1 0 19044 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_224
timestamp 1607721120
transform 1 0 21712 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_212
timestamp 1607721120
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_223
timestamp 1607721120
transform 1 0 21620 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1607721120
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1607721120
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607721120
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1607721120
transform 1 0 21344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0810_
timestamp 1607721120
transform 1 0 20884 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_245
timestamp 1607721120
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1607721120
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_232
timestamp 1607721120
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1607721120
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1607721120
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607721120
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607721120
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0813_
timestamp 1607721120
transform 1 0 22356 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1607721120
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_253
timestamp 1607721120
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607721120
transform -1 0 24840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607721120
transform -1 0 24840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1607721120
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607721120
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2116 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_39
timestamp 1607721120
transform 1 0 4692 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp 1607721120
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1607721120
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607721120
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 4324 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1607721120
transform 1 0 5428 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_2_78
timestamp 1607721120
transform 1 0 8280 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1607721120
transform 1 0 7176 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0610_
timestamp 1607721120
transform 1 0 7912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1607721120
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607721120
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1264_
timestamp 1607721120
transform 1 0 9660 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_112
timestamp 1607721120
transform 1 0 11408 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 12144 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1607721120
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_134
timestamp 1607721120
transform 1 0 13432 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1607721120
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_157
timestamp 1607721120
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607721120
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1607721120
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_178
timestamp 1607721120
transform 1 0 17480 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0821_
timestamp 1607721120
transform 1 0 18216 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0816_
timestamp 1607721120
transform 1 0 16652 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_207
timestamp 1607721120
transform 1 0 20148 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_195
timestamp 1607721120
transform 1 0 19044 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_227
timestamp 1607721120
transform 1 0 21988 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607721120
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1607721120
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607721120
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0809_
timestamp 1607721120
transform 1 0 22172 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_250
timestamp 1607721120
transform 1 0 24104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_238
timestamp 1607721120
transform 1 0 23000 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_254
timestamp 1607721120
transform 1 0 24472 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607721120
transform -1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1607721120
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1607721120
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607721120
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607721120
transform 1 0 1840 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1607721120
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1607721120
transform 1 0 3588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1120_
timestamp 1607721120
transform 1 0 4508 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1607721120
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1607721120
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607721120
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1259_
timestamp 1607721120
transform 1 0 7544 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_3_89
timestamp 1607721120
transform 1 0 9292 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1064_
timestamp 1607721120
transform 1 0 10028 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1607721120
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1607721120
transform 1 0 11500 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607721120
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0717_
timestamp 1607721120
transform 1 0 12420 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1607721120
transform 1 0 13708 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0837_
timestamp 1607721120
transform 1 0 14444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_165
timestamp 1607721120
transform 1 0 16284 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_154
timestamp 1607721120
transform 1 0 15272 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1607721120
transform 1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp 1607721120
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1607721120
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607721120
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 18308 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_206
timestamp 1607721120
transform 1 0 20056 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_194
timestamp 1607721120
transform 1 0 18952 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_226
timestamp 1607721120
transform 1 0 21896 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_218
timestamp 1607721120
transform 1 0 21160 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607721120
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1607721120
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_236
timestamp 1607721120
transform 1 0 22816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607721120
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_253
timestamp 1607721120
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607721120
transform -1 0 24840 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1607721120
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607721120
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0620_
timestamp 1607721120
transform 1 0 2116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1607721120
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1607721120
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1607721120
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607721120
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0618_
timestamp 1607721120
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1607721120
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_46
timestamp 1607721120
transform 1 0 5336 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1071_
timestamp 1607721120
transform 1 0 6624 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_76
timestamp 1607721120
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp 1607721120
transform 1 0 10028 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1607721120
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607721120
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1063_
timestamp 1607721120
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1607721120
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607721120
transform 1 0 10948 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607721120
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_126
timestamp 1607721120
transform 1 0 12696 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0709_
timestamp 1607721120
transform 1 0 13432 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_4_161
timestamp 1607721120
transform 1 0 15916 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607721120
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0725_
timestamp 1607721120
transform 1 0 15272 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_4_185
timestamp 1607721120
transform 1 0 18124 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_173
timestamp 1607721120
transform 1 0 17020 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1607721120
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_227
timestamp 1607721120
transform 1 0 21988 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607721120
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1607721120
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1607721120
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607721120
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_247
timestamp 1607721120
transform 1 0 23828 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_235
timestamp 1607721120
transform 1 0 22724 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0814_
timestamp 1607721120
transform 1 0 23000 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607721120
transform -1 0 24840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_14
timestamp 1607721120
transform 1 0 2392 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1607721120
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1607721120
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607721120
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1607721120
transform 1 0 2024 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1607721120
transform 1 0 4416 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3128 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1607721120
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607721120
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1074_
timestamp 1607721120
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0619_
timestamp 1607721120
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp 1607721120
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1607721120
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0710_
timestamp 1607721120
transform 1 0 8556 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_88
timestamp 1607721120
transform 1 0 9200 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0713_
timestamp 1607721120
transform 1 0 9936 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1607721120
transform 1 0 12420 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1607721120
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607721120
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1607721120
transform 1 0 12972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607721120
transform 1 0 13064 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_5_160
timestamp 1607721120
transform 1 0 15824 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1607721120
transform 1 0 14812 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1607721120
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607721120
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1607721120
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1607721120
transform 1 0 16928 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607721120
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1607721120
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1607721120
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1607721120
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1607721120
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1607721120
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607721120
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_253
timestamp 1607721120
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607721120
transform -1 0 24840 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1607721120
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1607721120
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607721120
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607721120
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607721120
transform 1 0 1380 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1607721120
transform 1 0 1472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0622_
timestamp 1607721120
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_22
timestamp 1607721120
transform 1 0 3128 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1607721120
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1607721120
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607721120
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1033_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _1032_
timestamp 1607721120
transform 1 0 3864 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1607721120
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_56
timestamp 1607721120
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1607721120
transform 1 0 5152 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_58
timestamp 1607721120
transform 1 0 6440 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607721120
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1073_
timestamp 1607721120
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_4  _1061_
timestamp 1607721120
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_78
timestamp 1607721120
transform 1 0 8280 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_75
timestamp 1607721120
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1087_
timestamp 1607721120
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1607721120
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1607721120
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1607721120
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607721120
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607721120
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0714_
timestamp 1607721120
transform 1 0 9568 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1607721120
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1607721120
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_106
timestamp 1607721120
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1607721120
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_112
timestamp 1607721120
transform 1 0 11408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607721120
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_142
timestamp 1607721120
transform 1 0 14168 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1607721120
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1607721120
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_128
timestamp 1607721120
transform 1 0 12880 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0727_
timestamp 1607721120
transform 1 0 12972 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0724_
timestamp 1607721120
transform 1 0 12880 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1607721120
transform 1 0 14904 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_157
timestamp 1607721120
transform 1 0 15548 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1607721120
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607721120
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1318_
timestamp 1607721120
transform 1 0 14996 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1607721120
transform 1 0 16284 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1607721120
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_187
timestamp 1607721120
transform 1 0 18308 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1607721120
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_170
timestamp 1607721120
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1607721120
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1607721120
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607721120
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1607721120
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_199
timestamp 1607721120
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1607721120
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_192
timestamp 1607721120
transform 1 0 18768 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_223
timestamp 1607721120
transform 1 0 21620 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1607721120
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1607721120
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1607721120
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1607721120
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607721120
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_245
timestamp 1607721120
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1607721120
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_235
timestamp 1607721120
transform 1 0 22724 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1607721120
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607721120
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_253
timestamp 1607721120
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_251
timestamp 1607721120
transform 1 0 24196 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607721120
transform -1 0 24840 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607721120
transform -1 0 24840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1607721120
transform 1 0 2944 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1607721120
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1607721120
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607721120
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0623_
timestamp 1607721120
transform 1 0 1840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1607721120
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1607721120
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607721120
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0612_
timestamp 1607721120
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1607721120
transform 1 0 5980 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1257_
timestamp 1607721120
transform 1 0 6716 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0604_
timestamp 1607721120
transform 1 0 5612 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1607721120
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_101
timestamp 1607721120
transform 1 0 10396 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1607721120
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607721120
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 9752 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_118
timestamp 1607721120
transform 1 0 11960 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1607721120
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607721120
transform 1 0 12696 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607721120
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0804_
timestamp 1607721120
transform 1 0 15272 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_8_183
timestamp 1607721120
transform 1 0 17940 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_168
timestamp 1607721120
transform 1 0 16560 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0800_
timestamp 1607721120
transform 1 0 17296 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1607721120
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_195
timestamp 1607721120
transform 1 0 19044 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1607721120
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1607721120
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1607721120
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607721120
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1607721120
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_251
timestamp 1607721120
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607721120
transform -1 0 24840 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_16
timestamp 1607721120
transform 1 0 2576 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1607721120
transform 1 0 2116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1607721120
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607721120
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1070_
timestamp 1607721120
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_33
timestamp 1607721120
transform 1 0 4140 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0615_
timestamp 1607721120
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1607721120
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1607721120
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607721120
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0616_
timestamp 1607721120
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_74
timestamp 1607721120
transform 1 0 7912 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_66
timestamp 1607721120
transform 1 0 7176 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1260_
timestamp 1607721120
transform 1 0 8004 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp 1607721120
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1607721120
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1607721120
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607721120
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1137_
timestamp 1607721120
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0708_
timestamp 1607721120
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp 1607721120
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1607721120
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1242_
timestamp 1607721120
transform 1 0 14260 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_162
timestamp 1607721120
transform 1 0 16008 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_187
timestamp 1607721120
transform 1 0 18308 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1607721120
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1607721120
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607721120
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1607721120
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1607721120
transform 1 0 16744 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_199
timestamp 1607721120
transform 1 0 19412 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_223
timestamp 1607721120
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_211
timestamp 1607721120
transform 1 0 20516 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_245
timestamp 1607721120
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1607721120
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_235
timestamp 1607721120
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607721120
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_253
timestamp 1607721120
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607721120
transform -1 0 24840 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607721120
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607721120
transform 1 0 1380 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1607721120
transform 1 0 4416 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1607721120
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_22
timestamp 1607721120
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607721120
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1607721120
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_55
timestamp 1607721120
transform 1 0 6164 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_44
timestamp 1607721120
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0641_
timestamp 1607721120
transform 1 0 5336 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_82
timestamp 1607721120
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6900 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1069_
timestamp 1607721120
transform 1 0 7176 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1607721120
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607721120
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1263_
timestamp 1607721120
transform 1 0 9660 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_10_112
timestamp 1607721120
transform 1 0 11408 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0721_
timestamp 1607721120
transform 1 0 12144 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1607721120
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_134
timestamp 1607721120
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1607721120
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_157
timestamp 1607721120
transform 1 0 15548 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607721120
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0802_
timestamp 1607721120
transform 1 0 16284 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1607721120
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_179
timestamp 1607721120
transform 1 0 17572 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1607721120
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1607721120
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1607721120
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1607721120
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607721120
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607721120
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1607721120
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_251
timestamp 1607721120
transform 1 0 24196 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607721120
transform -1 0 24840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1607721120
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607721120
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0617_
timestamp 1607721120
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1607721120
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_29
timestamp 1607721120
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_21
timestamp 1607721120
transform 1 0 3036 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1048_
timestamp 1607721120
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1607721120
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1607721120
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607721120
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1062_
timestamp 1607721120
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0640_
timestamp 1607721120
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1607721120
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_66
timestamp 1607721120
transform 1 0 7176 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1065_
timestamp 1607721120
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1607721120
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1607721120
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1136_
timestamp 1607721120
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1607721120
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1607721120
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1607721120
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607721120
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1607721120
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1607721120
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1243_
timestamp 1607721120
transform 1 0 14352 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _0722_
timestamp 1607721120
transform 1 0 12696 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1607721120
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_187
timestamp 1607721120
transform 1 0 18308 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1607721120
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1607721120
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607721120
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1607721120
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1607721120
transform 1 0 16836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_198
timestamp 1607721120
transform 1 0 19320 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1607721120
transform 1 0 19044 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_222
timestamp 1607721120
transform 1 0 21528 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_210
timestamp 1607721120
transform 1 0 20424 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1607721120
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1607721120
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_234
timestamp 1607721120
transform 1 0 22632 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607721120
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_253
timestamp 1607721120
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607721120
transform -1 0 24840 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_6
timestamp 1607721120
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607721120
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1213_
timestamp 1607721120
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1607721120
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1607721120
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1607721120
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607721120
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1119_
timestamp 1607721120
transform 1 0 4324 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1607721120
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1607721120
transform 1 0 6532 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_78
timestamp 1607721120
transform 1 0 8280 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1607721120
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1607721120
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_wb_clk_i
timestamp 1607721120
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607721120
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1607721120
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_107
timestamp 1607721120
transform 1 0 10948 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607721120
transform 1 0 11224 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1607721120
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1607721120
transform 1 0 12972 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0719_
timestamp 1607721120
transform 1 0 13708 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1607721120
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1607721120
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607721120
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1319_
timestamp 1607721120
transform 1 0 16008 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_181
timestamp 1607721120
transform 1 0 17756 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_203
timestamp 1607721120
transform 1 0 19780 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1607721120
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1607721120
transform 1 0 19504 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1607721120
transform 1 0 18492 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1607721120
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1607721120
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1607721120
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607721120
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1607721120
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_251
timestamp 1607721120
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607721120
transform -1 0 24840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1607721120
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1607721120
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607721120
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607721120
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607721120
transform 1 0 1840 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1215_
timestamp 1607721120
transform 1 0 1932 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1607721120
transform 1 0 4416 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1607721120
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1607721120
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1607721120
transform 1 0 3588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607721120
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1121_
timestamp 1607721120
transform 1 0 4508 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1607721120
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1607721120
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1607721120
transform 1 0 6808 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1607721120
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607721120
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1225_
timestamp 1607721120
transform 1 0 5336 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_77
timestamp 1607721120
transform 1 0 8188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_65
timestamp 1607721120
transform 1 0 7084 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1607721120
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1067_
timestamp 1607721120
transform 1 0 7452 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1066_
timestamp 1607721120
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1607721120
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_85
timestamp 1607721120
transform 1 0 8924 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607721120
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1262_
timestamp 1607721120
transform 1 0 9660 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1261_
timestamp 1607721120
transform 1 0 9660 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_112
timestamp 1607721120
transform 1 0 11408 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1607721120
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1607721120
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_wb_clk_i
timestamp 1607721120
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607721120
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1607721120
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1607721120
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1607721120
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_126
timestamp 1607721120
transform 1 0 12696 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1098_
timestamp 1607721120
transform 1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1097_
timestamp 1607721120
transform 1 0 13432 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_166
timestamp 1607721120
transform 1 0 16376 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1607721120
transform 1 0 15640 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1607721120
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_150
timestamp 1607721120
transform 1 0 14904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607721120
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1088_
timestamp 1607721120
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1607721120
transform 1 0 16192 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1607721120
transform 1 0 18308 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_176
timestamp 1607721120
transform 1 0 17296 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_187
timestamp 1607721120
transform 1 0 18308 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1607721120
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_168
timestamp 1607721120
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607721120
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0797_
timestamp 1607721120
transform 1 0 16468 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1607721120
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1607721120
transform 1 0 18032 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_198
timestamp 1607721120
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_198
timestamp 1607721120
transform 1 0 19320 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1607721120
transform 1 0 20056 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1607721120
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1607721120
transform 1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_218
timestamp 1607721120
transform 1 0 21160 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1607721120
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_221
timestamp 1607721120
transform 1 0 21436 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_209
timestamp 1607721120
transform 1 0 20332 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607721120
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1607721120
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_242
timestamp 1607721120
transform 1 0 23368 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_230
timestamp 1607721120
transform 1 0 22264 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1607721120
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_241
timestamp 1607721120
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_233
timestamp 1607721120
transform 1 0 22540 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607721120
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_254
timestamp 1607721120
transform 1 0 24472 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_253
timestamp 1607721120
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607721120
transform -1 0 24840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607721120
transform -1 0 24840 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1607721120
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1607721120
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607721120
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1214_
timestamp 1607721120
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_22
timestamp 1607721120
transform 1 0 3128 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1281_
timestamp 1607721120
transform 1 0 3864 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1607721120
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_49
timestamp 1607721120
transform 1 0 5612 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 6348 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607721120
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1607721120
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_65
timestamp 1607721120
transform 1 0 7084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1068_
timestamp 1607721120
transform 1 0 7820 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_97
timestamp 1607721120
transform 1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_89
timestamp 1607721120
transform 1 0 9292 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0732_
timestamp 1607721120
transform 1 0 10304 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1607721120
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1607721120
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607721120
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1099_
timestamp 1607721120
transform 1 0 13156 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1607721120
transform 1 0 14628 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0806_
timestamp 1607721120
transform 1 0 15364 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1607721120
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1607721120
transform 1 0 16652 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607721120
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1096_
timestamp 1607721120
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_199
timestamp 1607721120
transform 1 0 19412 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_188
timestamp 1607721120
transform 1 0 18400 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1607721120
transform 1 0 20148 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1607721120
transform 1 0 19136 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_222
timestamp 1607721120
transform 1 0 21528 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_210
timestamp 1607721120
transform 1 0 20424 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1607721120
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_242
timestamp 1607721120
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_234
timestamp 1607721120
transform 1 0 22632 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607721120
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_253
timestamp 1607721120
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607721120
transform -1 0 24840 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607721120
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607721120
transform 1 0 1380 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1607721120
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_22
timestamp 1607721120
transform 1 0 3128 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607721120
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1035_
timestamp 1607721120
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1607721120
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607721120
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0966_
timestamp 1607721120
transform 1 0 6624 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1607721120
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1607721120
transform 1 0 10672 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_96
timestamp 1607721120
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1607721120
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607721120
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1607721120
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_124
timestamp 1607721120
transform 1 0 12512 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607721120
transform 1 0 10764 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1607721120
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0718_
timestamp 1607721120
transform 1 0 13248 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1607721120
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607721120
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1317_
timestamp 1607721120
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_173
timestamp 1607721120
transform 1 0 17020 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1320_
timestamp 1607721120
transform 1 0 17756 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1607721120
transform 1 0 19504 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1607721120
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607721120
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1607721120
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607721120
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1607721120
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_251
timestamp 1607721120
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607721120
transform -1 0 24840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_18
timestamp 1607721120
transform 1 0 2760 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1607721120
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607721120
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0694_
timestamp 1607721120
transform 1 0 1472 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1607721120
transform 1 0 4232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1607721120
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1034_
timestamp 1607721120
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1607721120
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1607721120
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607721120
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0611_
timestamp 1607721120
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_74
timestamp 1607721120
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 1607721120
transform 1 0 7176 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1229_
timestamp 1607721120
transform 1 0 8188 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_17_96
timestamp 1607721120
transform 1 0 9936 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0706_
timestamp 1607721120
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1607721120
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1607721120
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607721120
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 1607721120
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1607721120
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1241_
timestamp 1607721120
transform 1 0 13892 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1607721120
transform 1 0 15640 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0771_
timestamp 1607721120
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1607721120
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607721120
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0793_
timestamp 1607721120
transform 1 0 18032 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_206
timestamp 1607721120
transform 1 0 20056 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1607721120
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0794_
timestamp 1607721120
transform 1 0 19412 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_218
timestamp 1607721120
transform 1 0 21160 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_245
timestamp 1607721120
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1607721120
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_230
timestamp 1607721120
transform 1 0 22264 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607721120
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_253
timestamp 1607721120
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607721120
transform -1 0 24840 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_6
timestamp 1607721120
transform 1 0 1656 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607721120
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0680_
timestamp 1607721120
transform 1 0 2392 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1607721120
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp 1607721120
transform 1 0 4416 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1607721120
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1607721120
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607721120
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1607721120
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_60
timestamp 1607721120
transform 1 0 6624 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1607721120
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0972_
timestamp 1607721120
transform 1 0 5336 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _1116_
timestamp 1607721120
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1607721120
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1607721120
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1607721120
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607721120
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 10304 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_18_113
timestamp 1607721120
transform 1 0 11500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1044_
timestamp 1607721120
transform 1 0 12512 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_140
timestamp 1607721120
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_164
timestamp 1607721120
transform 1 0 16192 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1607721120
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1607721120
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607721120
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0770_
timestamp 1607721120
transform 1 0 15824 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1607721120
transform 1 0 18216 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0799_
timestamp 1607721120
transform 1 0 16928 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1607721120
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1607721120
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1607721120
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1607721120
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1607721120
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1607721120
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607721120
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1607721120
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_251
timestamp 1607721120
transform 1 0 24196 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607721120
transform -1 0 24840 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_10
timestamp 1607721120
transform 1 0 2024 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607721120
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607721120
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607721120
transform 1 0 1380 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1145_
timestamp 1607721120
transform 1 0 1380 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1021_
timestamp 1607721120
transform 1 0 2760 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1607721120
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1607721120
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1607721120
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_25
timestamp 1607721120
transform 1 0 3404 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607721120
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1029_
timestamp 1607721120
transform 1 0 4140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0827_
timestamp 1607721120
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_45
timestamp 1607721120
transform 1 0 5244 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1607721120
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_45
timestamp 1607721120
transform 1 0 5244 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607721120
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0978_
timestamp 1607721120
transform 1 0 5980 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607721120
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_67
timestamp 1607721120
transform 1 0 7268 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_78
timestamp 1607721120
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1607721120
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0953_
timestamp 1607721120
transform 1 0 8372 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _0701_
timestamp 1607721120
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1607721120
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1607721120
transform 1 0 9660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607721120
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1230_
timestamp 1607721120
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_20_112
timestamp 1607721120
transform 1 0 11408 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1607721120
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1607721120
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1607721120
transform 1 0 11132 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1607721120
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607721120
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1283_
timestamp 1607721120
transform 1 0 12144 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0715_
timestamp 1607721120
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1607721120
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1275_
timestamp 1607721120
transform 1 0 12972 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1607721120
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1607721120
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_148
timestamp 1607721120
transform 1 0 14720 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607721120
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0782_
timestamp 1607721120
transform 1 0 15456 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_4  _0776_
timestamp 1607721120
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_186
timestamp 1607721120
transform 1 0 18216 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1607721120
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_187
timestamp 1607721120
transform 1 0 18308 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1607721120
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1607721120
transform 1 0 16652 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607721120
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0796_
timestamp 1607721120
transform 1 0 16928 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1607721120
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_198
timestamp 1607721120
transform 1 0 19320 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_198
timestamp 1607721120
transform 1 0 19320 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1607721120
transform 1 0 19044 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1607721120
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1607721120
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1607721120
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_222
timestamp 1607721120
transform 1 0 21528 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_210
timestamp 1607721120
transform 1 0 20424 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607721120
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1607721120
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_245
timestamp 1607721120
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1607721120
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_234
timestamp 1607721120
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607721120
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_251
timestamp 1607721120
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_253
timestamp 1607721120
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607721120
transform -1 0 24840 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607721120
transform -1 0 24840 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_12
timestamp 1607721120
transform 1 0 2208 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1607721120
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1607721120
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607721120
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1265_
timestamp 1607721120
transform 1 0 2944 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1057_
timestamp 1607721120
transform 1 0 1840 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_39
timestamp 1607721120
transform 1 0 4692 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1607721120
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1607721120
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607721120
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1111_
timestamp 1607721120
transform 1 0 5612 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0807_
timestamp 1607721120
transform 1 0 6808 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1607721120
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1607721120
transform 1 0 7452 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1115_
timestamp 1607721120
transform 1 0 8280 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1607721120
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_94
timestamp 1607721120
transform 1 0 9752 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1607721120
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1607721120
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_106
timestamp 1607721120
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607721120
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1607721120
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0626_
timestamp 1607721120
transform 1 0 12512 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_140
timestamp 1607721120
transform 1 0 13984 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_128
timestamp 1607721120
transform 1 0 12880 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1043_
timestamp 1607721120
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_152
timestamp 1607721120
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1244_
timestamp 1607721120
transform 1 0 15272 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_187
timestamp 1607721120
transform 1 0 18308 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1607721120
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1607721120
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607721120
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1607721120
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_198
timestamp 1607721120
transform 1 0 19320 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1607721120
transform 1 0 19044 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_222
timestamp 1607721120
transform 1 0 21528 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_210
timestamp 1607721120
transform 1 0 20424 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_245
timestamp 1607721120
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1607721120
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_234
timestamp 1607721120
transform 1 0 22632 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607721120
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_253
timestamp 1607721120
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607721120
transform -1 0 24840 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_18
timestamp 1607721120
transform 1 0 2760 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1607721120
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607721120
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0692_
timestamp 1607721120
transform 1 0 1472 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1607721120
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1607721120
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607721120
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1316_
timestamp 1607721120
transform 1 0 4784 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_59
timestamp 1607721120
transform 1 0 6532 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_83
timestamp 1607721120
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1117_
timestamp 1607721120
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1607721120
transform 1 0 10028 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1607721120
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607721120
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1114_
timestamp 1607721120
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_105
timestamp 1607721120
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 11040 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1046_
timestamp 1607721120
transform 1 0 11316 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_138
timestamp 1607721120
transform 1 0 13800 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_127
timestamp 1607721120
transform 1 0 12788 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1607721120
transform 1 0 13524 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_162
timestamp 1607721120
transform 1 0 16008 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1607721120
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1607721120
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1607721120
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607721120
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1607721120
transform 1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1321_
timestamp 1607721120
transform 1 0 16744 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1607721120
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_189
timestamp 1607721120
transform 1 0 18492 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1607721120
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1607721120
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1607721120
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607721120
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1607721120
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_251
timestamp 1607721120
transform 1 0 24196 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607721120
transform -1 0 24840 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_13
timestamp 1607721120
transform 1 0 2300 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1607721120
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607721120
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0687_
timestamp 1607721120
transform 1 0 1656 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_23_37
timestamp 1607721120
transform 1 0 4508 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1060_
timestamp 1607721120
transform 1 0 3036 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1607721120
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_52
timestamp 1607721120
transform 1 0 5888 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607721120
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1228_
timestamp 1607721120
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0826_
timestamp 1607721120
transform 1 0 5244 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1607721120
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1607721120
transform 1 0 10580 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0948_
timestamp 1607721120
transform 1 0 9292 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1607721120
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607721120
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1045_
timestamp 1607721120
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1607721120
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_139
timestamp 1607721120
transform 1 0 13892 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1607721120
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1095_
timestamp 1607721120
transform 1 0 14628 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_187
timestamp 1607721120
transform 1 0 18308 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607721120
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1607721120
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607721120
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1607721120
transform 1 0 16836 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1607721120
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_198
timestamp 1607721120
transform 1 0 19320 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1607721120
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_222
timestamp 1607721120
transform 1 0 21528 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_210
timestamp 1607721120
transform 1 0 20424 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_245
timestamp 1607721120
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1607721120
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_234
timestamp 1607721120
transform 1 0 22632 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607721120
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_253
timestamp 1607721120
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607721120
transform -1 0 24840 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_19
timestamp 1607721120
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1607721120
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607721120
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0690_
timestamp 1607721120
transform 1 0 1564 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1607721120
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1607721120
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607721120
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1023_
timestamp 1607721120
transform 1 0 4692 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1607721120
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1607721120
transform 1 0 5796 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0961_
timestamp 1607721120
transform 1 0 6716 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_24_83
timestamp 1607721120
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1607721120
transform 1 0 8004 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_96
timestamp 1607721120
transform 1 0 9936 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1607721120
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 8924 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607721120
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1273_
timestamp 1607721120
transform 1 0 10672 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1607721120
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_123
timestamp 1607721120
transform 1 0 12420 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1607721120
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0871_
timestamp 1607721120
transform 1 0 13156 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607721120
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0876_
timestamp 1607721120
transform 1 0 15272 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp 1607721120
transform 1 0 18124 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1607721120
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0783_
timestamp 1607721120
transform 1 0 17296 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1607721120
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_196
timestamp 1607721120
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1607721120
transform 1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1607721120
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1607721120
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607721120
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1607721120
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_251
timestamp 1607721120
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607721120
transform -1 0 24840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_20
timestamp 1607721120
transform 1 0 2944 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1607721120
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607721120
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0684_
timestamp 1607721120
transform 1 0 2116 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1267_
timestamp 1607721120
transform 1 0 3680 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1607721120
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1607721120
transform 1 0 5428 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 6164 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607721120
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1169_
timestamp 1607721120
transform 1 0 6808 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1607721120
transform 1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1170_
timestamp 1607721120
transform 1 0 8188 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1607721120
transform 1 0 9568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_84
timestamp 1607721120
transform 1 0 8832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1232_
timestamp 1607721120
transform 1 0 9660 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1607721120
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_112
timestamp 1607721120
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607721120
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1274_
timestamp 1607721120
transform 1 0 12420 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_25_142
timestamp 1607721120
transform 1 0 14168 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_164
timestamp 1607721120
transform 1 0 16192 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0882_
timestamp 1607721120
transform 1 0 14904 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1607721120
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607721120
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1143_
timestamp 1607721120
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1607721120
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1607721120
transform 1 0 19964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1607721120
transform 1 0 18860 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1607721120
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_217
timestamp 1607721120
transform 1 0 21068 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1607721120
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_241
timestamp 1607721120
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607721120
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_253
timestamp 1607721120
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607721120
transform -1 0 24840 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_8
timestamp 1607721120
transform 1 0 1840 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1607721120
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607721120
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607721120
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607721120
transform 1 0 1380 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1607721120
transform 1 0 1564 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0657_
timestamp 1607721120
transform 1 0 2576 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_36
timestamp 1607721120
transform 1 0 4416 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_25
timestamp 1607721120
transform 1 0 3404 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1607721120
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_22
timestamp 1607721120
transform 1 0 3128 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607721120
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1058_
timestamp 1607721120
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1607721120
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1607721120
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1607721120
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_60
timestamp 1607721120
transform 1 0 6624 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_48
timestamp 1607721120
transform 1 0 5520 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607721120
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0648_
timestamp 1607721120
transform 1 0 6256 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _0643_
timestamp 1607721120
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_73
timestamp 1607721120
transform 1 0 7820 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1166_
timestamp 1607721120
transform 1 0 7176 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1113_
timestamp 1607721120
transform 1 0 7360 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1112_
timestamp 1607721120
transform 1 0 8556 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_27_97
timestamp 1607721120
transform 1 0 10028 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1607721120
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607721120
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0936_
timestamp 1607721120
transform 1 0 9660 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1607721120
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_112
timestamp 1607721120
transform 1 0 11408 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_122
timestamp 1607721120
transform 1 0 12328 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_107
timestamp 1607721120
transform 1 0 10948 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607721120
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1199_
timestamp 1607721120
transform 1 0 12420 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1197_
timestamp 1607721120
transform 1 0 11684 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1196_
timestamp 1607721120
transform 1 0 10764 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1607721120
transform 1 0 14076 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1607721120
transform 1 0 13064 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_137
timestamp 1607721120
transform 1 0 13708 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_wb_clk_i
timestamp 1607721120
transform 1 0 14444 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_wb_clk_i
timestamp 1607721120
transform 1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1200_
timestamp 1607721120
transform 1 0 13064 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1607721120
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1607721120
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1607721120
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1607721120
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1607721120
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607721120
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1245_
timestamp 1607721120
transform 1 0 15732 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1094_
timestamp 1607721120
transform 1 0 14628 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1607721120
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_178
timestamp 1607721120
transform 1 0 17480 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607721120
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1092_
timestamp 1607721120
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1607721120
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1607721120
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_199
timestamp 1607721120
transform 1 0 19412 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_188
timestamp 1607721120
transform 1 0 18400 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1607721120
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_189
timestamp 1607721120
transform 1 0 18492 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1607721120
transform 1 0 19228 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1607721120
transform 1 0 19136 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_223
timestamp 1607721120
transform 1 0 21620 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1607721120
transform 1 0 20516 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1607721120
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1607721120
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1607721120
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607721120
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1607721120
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1607721120
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_235
timestamp 1607721120
transform 1 0 22724 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1607721120
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607721120
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_253
timestamp 1607721120
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_251
timestamp 1607721120
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607721120
transform -1 0 24840 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607721120
transform -1 0 24840 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1607721120
transform 1 0 2852 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1607721120
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607721120
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0686_
timestamp 1607721120
transform 1 0 1564 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_28_38
timestamp 1607721120
transform 1 0 4600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1607721120
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1607721120
transform 1 0 3588 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607721120
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1607721120
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_46
timestamp 1607721120
transform 1 0 5336 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607721120
transform 1 0 5428 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1607721120
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_66
timestamp 1607721120
transform 1 0 7176 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1171_
timestamp 1607721120
transform 1 0 7912 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1607721120
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1607721120
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1607721120
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607721120
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1201_
timestamp 1607721120
transform 1 0 10580 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_112
timestamp 1607721120
transform 1 0 11408 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1276_
timestamp 1607721120
transform 1 0 12144 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_28_139
timestamp 1607721120
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1607721120
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607721120
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1093_
timestamp 1607721120
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp 1607721120
transform 1 0 17848 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_170
timestamp 1607721120
transform 1 0 16744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1039_
timestamp 1607721120
transform 1 0 17480 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_205
timestamp 1607721120
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_193
timestamp 1607721120
transform 1 0 18860 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1607721120
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1607721120
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1607721120
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1607721120
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607721120
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1607721120
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_251
timestamp 1607721120
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607721120
transform -1 0 24840 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_15
timestamp 1607721120
transform 1 0 2484 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1607721120
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1607721120
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607721120
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0681_
timestamp 1607721120
transform 1 0 1840 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1266_
timestamp 1607721120
transform 1 0 3220 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1607721120
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_42
timestamp 1607721120
transform 1 0 4968 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607721120
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1607721120
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0629_
timestamp 1607721120
transform 1 0 6808 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_29_77
timestamp 1607721120
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_69
timestamp 1607721120
transform 1 0 7452 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1231_
timestamp 1607721120
transform 1 0 8280 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_97
timestamp 1607721120
transform 1 0 10028 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1607721120
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1607721120
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607721120
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1202_
timestamp 1607721120
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _1042_
timestamp 1607721120
transform 1 0 12604 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1607721120
transform 1 0 14076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_153
timestamp 1607721120
transform 1 0 15180 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1246_
timestamp 1607721120
transform 1 0 15456 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_175
timestamp 1607721120
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607721120
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0784_
timestamp 1607721120
transform 1 0 18032 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_29_202
timestamp 1607721120
transform 1 0 19688 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_191
timestamp 1607721120
transform 1 0 18676 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1607721120
transform 1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_226
timestamp 1607721120
transform 1 0 21896 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_214
timestamp 1607721120
transform 1 0 20792 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1607721120
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_238
timestamp 1607721120
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607721120
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1607721120
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607721120
transform -1 0 24840 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607721120
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607721120
transform 1 0 1380 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1607721120
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_22
timestamp 1607721120
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607721120
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1059_
timestamp 1607721120
transform 1 0 4048 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_48
timestamp 1607721120
transform 1 0 5520 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0642_
timestamp 1607721120
transform 1 0 6256 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1607721120
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_70
timestamp 1607721120
transform 1 0 7544 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0928_
timestamp 1607721120
transform 1 0 8280 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1607721120
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607721120
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0942_
timestamp 1607721120
transform 1 0 9660 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_30_122
timestamp 1607721120
transform 1 0 12328 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1607721120
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1173_
timestamp 1607721120
transform 1 0 11684 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1607721120
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_130
timestamp 1607721120
transform 1 0 13064 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0863_
timestamp 1607721120
transform 1 0 13156 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1607721120
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_158
timestamp 1607721120
transform 1 0 15640 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607721120
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1036_
timestamp 1607721120
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1607721120
transform 1 0 18308 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1322_
timestamp 1607721120
transform 1 0 16560 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1607721120
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1607721120
transform 1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607721120
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1607721120
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1607721120
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607721120
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1607721120
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_251
timestamp 1607721120
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607721120
transform -1 0 24840 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_9
timestamp 1607721120
transform 1 0 1932 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1607721120
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607721120
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1134_
timestamp 1607721120
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1607721120
transform 1 0 1656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_26
timestamp 1607721120
transform 1 0 3496 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0662_
timestamp 1607721120
transform 1 0 4232 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_55
timestamp 1607721120
transform 1 0 6164 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1607721120
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607721120
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0638_
timestamp 1607721120
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1607721120
transform 1 0 8740 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_66
timestamp 1607721120
transform 1 0 7176 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1168_
timestamp 1607721120
transform 1 0 7912 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_94
timestamp 1607721120
transform 1 0 9752 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1198_
timestamp 1607721120
transform 1 0 10488 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1607721120
transform 1 0 9476 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1607721120
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1607721120
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1607721120
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607721120
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1040_
timestamp 1607721120
transform 1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_147
timestamp 1607721120
transform 1 0 14628 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0852_
timestamp 1607721120
transform 1 0 15364 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1607721120
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1607721120
transform 1 0 16652 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607721120
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0781_
timestamp 1607721120
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1607721120
transform 1 0 19964 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1607721120
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1607721120
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1607721120
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1607721120
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1607721120
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607721120
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_253
timestamp 1607721120
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607721120
transform -1 0 24840 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_6
timestamp 1607721120
transform 1 0 1656 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607721120
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0669_
timestamp 1607721120
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1607721120
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_39
timestamp 1607721120
transform 1 0 4692 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1607721120
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1607721120
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607721120
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1146_
timestamp 1607721120
transform 1 0 4324 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607721120
transform 1 0 5428 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_32_74
timestamp 1607721120
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_66
timestamp 1607721120
transform 1 0 7176 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1172_
timestamp 1607721120
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_100
timestamp 1607721120
transform 1 0 10304 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1607721120
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607721120
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1167_
timestamp 1607721120
transform 1 0 9660 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_32_108
timestamp 1607721120
transform 1 0 11040 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1277_
timestamp 1607721120
transform 1 0 11316 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1607721120
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1607721120
transform 1 0 13064 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1203_
timestamp 1607721120
transform 1 0 13800 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1607721120
transform 1 0 15640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607721120
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1607721120
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_184
timestamp 1607721120
transform 1 0 18032 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0792_
timestamp 1607721120
transform 1 0 16744 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_32_207
timestamp 1607721120
transform 1 0 20148 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_195
timestamp 1607721120
transform 1 0 19044 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1607721120
transform 1 0 18768 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1607721120
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1607721120
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1607721120
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607721120
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1607721120
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_251
timestamp 1607721120
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607721120
transform -1 0 24840 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_19
timestamp 1607721120
transform 1 0 2852 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1607721120
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607721120
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607721120
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607721120
transform 1 0 1380 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0683_
timestamp 1607721120
transform 1 0 1564 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_34_30
timestamp 1607721120
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_22
timestamp 1607721120
transform 1 0 3128 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_31
timestamp 1607721120
transform 1 0 3956 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607721120
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1233_
timestamp 1607721120
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _0668_
timestamp 1607721120
transform 1 0 4508 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1607721120
transform 1 0 5796 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_58
timestamp 1607721120
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_50
timestamp 1607721120
transform 1 0 5704 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607721120
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0651_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6532 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _0628_
timestamp 1607721120
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_34_76
timestamp 1607721120
transform 1 0 8096 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1607721120
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_71
timestamp 1607721120
transform 1 0 7636 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0635_
timestamp 1607721120
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_102
timestamp 1607721120
transform 1 0 10488 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1607721120
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1607721120
transform 1 0 10488 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1607721120
transform 1 0 8924 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607721120
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1178_
timestamp 1607721120
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1175_
timestamp 1607721120
transform 1 0 9660 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_113
timestamp 1607721120
transform 1 0 11500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1607721120
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_114
timestamp 1607721120
transform 1 0 11592 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607721120
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1041_
timestamp 1607721120
transform 1 0 12236 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0760_
timestamp 1607721120
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1607721120
transform 1 0 11224 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_137
timestamp 1607721120
transform 1 0 13708 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1278_
timestamp 1607721120
transform 1 0 13156 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_34_161
timestamp 1607721120
transform 1 0 15916 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1607721120
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_150
timestamp 1607721120
transform 1 0 14904 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607721120
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1204_
timestamp 1607721120
transform 1 0 15272 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _0858_
timestamp 1607721120
transform 1 0 15640 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1607721120
transform 1 0 16652 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_180
timestamp 1607721120
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_172
timestamp 1607721120
transform 1 0 16928 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607721120
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1323_
timestamp 1607721120
transform 1 0 16744 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _1142_
timestamp 1607721120
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1607721120
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_189
timestamp 1607721120
transform 1 0 18492 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_204
timestamp 1607721120
transform 1 0 19872 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1607721120
transform 1 0 18860 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1607721120
transform 1 0 19596 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1607721120
transform 1 0 19228 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1607721120
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1607721120
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1607721120
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_228
timestamp 1607721120
transform 1 0 22080 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_216
timestamp 1607721120
transform 1 0 20976 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607721120
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1607721120
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_245
timestamp 1607721120
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1607721120
transform 1 0 23184 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607721120
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_251
timestamp 1607721120
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_253
timestamp 1607721120
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607721120
transform -1 0 24840 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607721120
transform -1 0 24840 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_14
timestamp 1607721120
transform 1 0 2392 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1607721120
transform 1 0 1932 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1607721120
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607721120
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1607721120
transform 1 0 2024 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_38
timestamp 1607721120
transform 1 0 4600 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1110_
timestamp 1607721120
transform 1 0 3128 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_53
timestamp 1607721120
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607721120
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0652_
timestamp 1607721120
transform 1 0 5336 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0645_
timestamp 1607721120
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_83
timestamp 1607721120
transform 1 0 8740 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_66
timestamp 1607721120
transform 1 0 7176 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1180_
timestamp 1607721120
transform 1 0 7912 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_100
timestamp 1607721120
transform 1 0 10304 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1179_
timestamp 1607721120
transform 1 0 9476 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_114
timestamp 1607721120
transform 1 0 11592 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1607721120
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607721120
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1205_
timestamp 1607721120
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0631_
timestamp 1607721120
transform 1 0 11224 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_144
timestamp 1607721120
transform 1 0 14352 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_132
timestamp 1607721120
transform 1 0 13248 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0672_
timestamp 1607721120
transform 1 0 13984 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1091_
timestamp 1607721120
transform 1 0 15088 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_35_180
timestamp 1607721120
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1607721120
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607721120
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0790_
timestamp 1607721120
transform 1 0 18032 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_35_198
timestamp 1607721120
transform 1 0 19320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1607721120
transform 1 0 20056 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_221
timestamp 1607721120
transform 1 0 21436 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_209
timestamp 1607721120
transform 1 0 20332 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1607721120
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_241
timestamp 1607721120
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1607721120
transform 1 0 22540 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607721120
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_253
timestamp 1607721120
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607721120
transform -1 0 24840 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_11
timestamp 1607721120
transform 1 0 2116 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1607721120
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607721120
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1607721120
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0673_
timestamp 1607721120
transform 1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1607721120
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_23
timestamp 1607721120
transform 1 0 3220 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607721120
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1024_
timestamp 1607721120
transform 1 0 4324 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1607721120
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_48
timestamp 1607721120
transform 1 0 5520 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0637_
timestamp 1607721120
transform 1 0 6808 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_36_69
timestamp 1607721120
transform 1 0 7452 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1176_
timestamp 1607721120
transform 1 0 8188 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_36_101
timestamp 1607721120
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_93
timestamp 1607721120
transform 1 0 9660 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_84
timestamp 1607721120
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607721120
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1210_
timestamp 1607721120
transform 1 0 10580 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_112
timestamp 1607721120
transform 1 0 11408 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1279_
timestamp 1607721120
transform 1 0 12144 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_36_139
timestamp 1607721120
transform 1 0 13892 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_162
timestamp 1607721120
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_154
timestamp 1607721120
transform 1 0 15272 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1607721120
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607721120
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1247_
timestamp 1607721120
transform 1 0 16192 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_36_183
timestamp 1607721120
transform 1 0 17940 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1607721120
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_195
timestamp 1607721120
transform 1 0 19044 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1607721120
transform 1 0 18676 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1607721120
transform 1 0 19780 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1607721120
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1607721120
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607721120
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1607721120
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_251
timestamp 1607721120
transform 1 0 24196 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607721120
transform -1 0 24840 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_10
timestamp 1607721120
transform 1 0 2024 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1607721120
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607721120
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1133_
timestamp 1607721120
transform 1 0 2760 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0930_
timestamp 1607721120
transform 1 0 1656 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_39
timestamp 1607721120
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1607721120
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0650_
timestamp 1607721120
transform 1 0 4876 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_53
timestamp 1607721120
transform 1 0 5980 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607721120
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0646_
timestamp 1607721120
transform 1 0 6808 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1607721120
transform 1 0 7452 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0654_
timestamp 1607721120
transform 1 0 8188 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_37_96
timestamp 1607721120
transform 1 0 9936 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_84
timestamp 1607721120
transform 1 0 8832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1209_
timestamp 1607721120
transform 1 0 10672 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0627_
timestamp 1607721120
transform 1 0 9568 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_123
timestamp 1607721120
transform 1 0 12420 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1607721120
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1607721120
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607721120
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1038_
timestamp 1607721120
transform 1 0 13156 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_147
timestamp 1607721120
transform 1 0 14628 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0845_
timestamp 1607721120
transform 1 0 15364 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_37_181
timestamp 1607721120
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1607721120
transform 1 0 16652 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607721120
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0785_
timestamp 1607721120
transform 1 0 18032 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_37_202
timestamp 1607721120
transform 1 0 19688 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_191
timestamp 1607721120
transform 1 0 18676 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1607721120
transform 1 0 19412 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_226
timestamp 1607721120
transform 1 0 21896 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_214
timestamp 1607721120
transform 1 0 20792 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1607721120
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_238
timestamp 1607721120
transform 1 0 23000 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607721120
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1607721120
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607721120
transform -1 0 24840 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607721120
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607721120
transform 1 0 1380 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_38_30
timestamp 1607721120
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_22
timestamp 1607721120
transform 1 0 3128 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607721120
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1109_
timestamp 1607721120
transform 1 0 4048 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_60
timestamp 1607721120
transform 1 0 6624 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_48
timestamp 1607721120
transform 1 0 5520 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_64
timestamp 1607721120
transform 1 0 6992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1349_
timestamp 1607721120
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_103
timestamp 1607721120
transform 1 0 10580 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1607721120
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1607721120
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607721120
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1174_
timestamp 1607721120
transform 1 0 9936 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1124_
timestamp 1607721120
transform 1 0 11316 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_38_142
timestamp 1607721120
transform 1 0 14168 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_127
timestamp 1607721120
transform 1 0 12788 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1607721120
transform 1 0 13524 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_38_161
timestamp 1607721120
transform 1 0 15916 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1607721120
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607721120
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1207_
timestamp 1607721120
transform 1 0 15272 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_38_178
timestamp 1607721120
transform 1 0 17480 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_169
timestamp 1607721120
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0839_
timestamp 1607721120
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0787_
timestamp 1607721120
transform 1 0 16836 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1607721120
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_190
timestamp 1607721120
transform 1 0 18584 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1148_
timestamp 1607721120
transform 1 0 19320 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1607721120
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1607721120
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607721120
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1607721120
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_251
timestamp 1607721120
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607721120
transform -1 0 24840 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_6
timestamp 1607721120
transform 1 0 1656 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_18
timestamp 1607721120
transform 1 0 2760 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1607721120
transform 1 0 1380 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607721120
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607721120
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0679_
timestamp 1607721120
transform 1 0 1472 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1607721120
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0670_
timestamp 1607721120
transform 1 0 2392 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_40_32
timestamp 1607721120
transform 1 0 4048 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1607721120
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_21
timestamp 1607721120
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_30
timestamp 1607721120
transform 1 0 3864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607721120
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1234_
timestamp 1607721120
transform 1 0 4600 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _1017_
timestamp 1607721120
transform 1 0 4140 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_40_57
timestamp 1607721120
transform 1 0 6348 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1607721120
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_47
timestamp 1607721120
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607721120
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0655_
timestamp 1607721120
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_72
timestamp 1607721120
transform 1 0 7728 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_71
timestamp 1607721120
transform 1 0 7636 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1152_
timestamp 1607721120
transform 1 0 8372 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0653_
timestamp 1607721120
transform 1 0 7084 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0624_
timestamp 1607721120
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_84
timestamp 1607721120
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1607721120
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1607721120
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607721120
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1208_
timestamp 1607721120
transform 1 0 10304 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1186_
timestamp 1607721120
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1177_
timestamp 1607721120
transform 1 0 10488 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_40_117
timestamp 1607721120
transform 1 0 11868 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1607721120
transform 1 0 11132 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1607721120
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_109
timestamp 1607721120
transform 1 0 11132 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607721120
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1607721120
transform 1 0 11960 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0633_
timestamp 1607721120
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_137
timestamp 1607721120
transform 1 0 13708 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_127
timestamp 1607721120
transform 1 0 12788 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1037_
timestamp 1607721120
transform 1 0 13524 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1607721120
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_151
timestamp 1607721120
transform 1 0 14996 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607721120
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1090_
timestamp 1607721120
transform 1 0 15272 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0840_
timestamp 1607721120
transform 1 0 15732 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1607721120
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1607721120
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_173
timestamp 1607721120
transform 1 0 17020 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607721120
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0834_
timestamp 1607721120
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0788_
timestamp 1607721120
transform 1 0 17480 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_40_203
timestamp 1607721120
transform 1 0 19780 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1607721120
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_200
timestamp 1607721120
transform 1 0 19504 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_188
timestamp 1607721120
transform 1 0 18400 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1157_
timestamp 1607721120
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1607721120
transform 1 0 19504 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1607721120
transform 1 0 20240 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1607721120
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1607721120
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1607721120
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_223
timestamp 1607721120
transform 1 0 21620 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_211
timestamp 1607721120
transform 1 0 20516 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607721120
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1607721120
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1607721120
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1607721120
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_235
timestamp 1607721120
transform 1 0 22724 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607721120
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_251
timestamp 1607721120
transform 1 0 24196 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1607721120
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607721120
transform -1 0 24840 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607721120
transform -1 0 24840 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_18
timestamp 1607721120
transform 1 0 2760 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1607721120
transform 1 0 1380 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607721120
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0671_
timestamp 1607721120
transform 1 0 2116 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1108_
timestamp 1607721120
transform 1 0 3496 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1607721120
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_53
timestamp 1607721120
transform 1 0 5980 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_42
timestamp 1607721120
transform 1 0 4968 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607721120
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1607721120
transform 1 0 5704 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1607721120
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_66
timestamp 1607721120
transform 1 0 7176 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1147_
timestamp 1607721120
transform 1 0 7268 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_41_86
timestamp 1607721120
transform 1 0 9016 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 9108 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_41_114
timestamp 1607721120
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607721120
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1184_
timestamp 1607721120
transform 1 0 12420 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1181_
timestamp 1607721120
transform 1 0 10948 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_41_138
timestamp 1607721120
transform 1 0 13800 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_130
timestamp 1607721120
transform 1 0 13064 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1280_
timestamp 1607721120
transform 1 0 14076 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1607721120
transform 1 0 15824 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1607721120
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_172
timestamp 1607721120
transform 1 0 16928 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607721120
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1153_
timestamp 1607721120
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1122_
timestamp 1607721120
transform 1 0 16560 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_199
timestamp 1607721120
transform 1 0 19412 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_188
timestamp 1607721120
transform 1 0 18400 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1607721120
transform 1 0 19136 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_223
timestamp 1607721120
transform 1 0 21620 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_211
timestamp 1607721120
transform 1 0 20516 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1607721120
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1607721120
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_235
timestamp 1607721120
transform 1 0 22724 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607721120
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_253
timestamp 1607721120
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607721120
transform -1 0 24840 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_17
timestamp 1607721120
transform 1 0 2668 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607721120
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0677_
timestamp 1607721120
transform 1 0 1380 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_42_32
timestamp 1607721120
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1607721120
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607721120
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1235_
timestamp 1607721120
transform 1 0 4416 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_42_55
timestamp 1607721120
transform 1 0 6164 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_72
timestamp 1607721120
transform 1 0 7728 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1155_
timestamp 1607721120
transform 1 0 6900 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0625_
timestamp 1607721120
transform 1 0 8464 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_100
timestamp 1607721120
transform 1 0 10304 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_84
timestamp 1607721120
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607721120
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1154_
timestamp 1607721120
transform 1 0 9660 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_124
timestamp 1607721120
transform 1 0 12512 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1123_
timestamp 1607721120
transform 1 0 11040 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_139
timestamp 1607721120
transform 1 0 13892 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1185_
timestamp 1607721120
transform 1 0 13248 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_154
timestamp 1607721120
transform 1 0 15272 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1607721120
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607721120
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1248_
timestamp 1607721120
transform 1 0 16008 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_42_181
timestamp 1607721120
transform 1 0 17756 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_205
timestamp 1607721120
transform 1 0 19964 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_193
timestamp 1607721120
transform 1 0 18860 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1607721120
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1607721120
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_213
timestamp 1607721120
transform 1 0 20700 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607721120
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1607721120
transform 1 0 23092 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_251
timestamp 1607721120
transform 1 0 24196 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607721120
transform -1 0 24840 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607721120
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607721120
transform 1 0 1380 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_43_30
timestamp 1607721120
transform 1 0 3864 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_22
timestamp 1607721120
transform 1 0 3128 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1012_
timestamp 1607721120
transform 1 0 3956 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1607721120
transform 1 0 6808 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1607721120
transform 1 0 6348 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_45
timestamp 1607721120
transform 1 0 5244 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607721120
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_79
timestamp 1607721120
transform 1 0 8372 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1150_
timestamp 1607721120
transform 1 0 7544 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_43_90
timestamp 1607721120
transform 1 0 9384 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1183_
timestamp 1607721120
transform 1 0 10120 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1607721120
transform 1 0 9108 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_119
timestamp 1607721120
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_107
timestamp 1607721120
transform 1 0 10948 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607721120
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1077_
timestamp 1607721120
transform 1 0 12420 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_43_139
timestamp 1607721120
transform 1 0 13892 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_161
timestamp 1607721120
transform 1 0 15916 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0888_
timestamp 1607721120
transform 1 0 14628 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1607721120
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_180
timestamp 1607721120
transform 1 0 17664 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_172
timestamp 1607721120
transform 1 0 16928 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607721120
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1607721120
transform 1 0 16652 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1607721120
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1607721120
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1607721120
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_245
timestamp 1607721120
transform 1 0 23644 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1607721120
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607721120
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_253
timestamp 1607721120
transform 1 0 24380 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607721120
transform -1 0 24840 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1607721120
transform 1 0 1380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607721120
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0676_
timestamp 1607721120
transform 1 0 1748 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_44_39
timestamp 1607721120
transform 1 0 4692 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1607721120
transform 1 0 3772 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_21
timestamp 1607721120
transform 1 0 3036 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607721120
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0675_
timestamp 1607721120
transform 1 0 4048 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_44_51
timestamp 1607721120
transform 1 0 5796 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0983_
timestamp 1607721120
transform 1 0 5888 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_44_83
timestamp 1607721120
transform 1 0 8740 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_66
timestamp 1607721120
transform 1 0 7176 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1156_
timestamp 1607721120
transform 1 0 7912 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_102
timestamp 1607721120
transform 1 0 10488 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1607721120
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607721120
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1187_
timestamp 1607721120
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1607721120
transform 1 0 11224 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1607721120
transform 1 0 14352 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1607721120
transform 1 0 12972 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1191_
timestamp 1607721120
transform 1 0 13708 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_44_158
timestamp 1607721120
transform 1 0 15640 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1607721120
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607721120
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1324_
timestamp 1607721120
transform 1 0 16376 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607721120
transform 1 0 15272 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_185
timestamp 1607721120
transform 1 0 18124 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1607721120
transform 1 0 19228 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1607721120
transform 1 0 21988 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1607721120
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1607721120
transform 1 0 20700 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1607721120
transform 1 0 20332 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607721120
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1607721120
transform 1 0 23092 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_251
timestamp 1607721120
transform 1 0 24196 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607721120
transform -1 0 24840 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_11
timestamp 1607721120
transform 1 0 2116 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1607721120
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607721120
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1272_
timestamp 1607721120
transform 1 0 2852 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0988_
timestamp 1607721120
transform 1 0 1748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_38
timestamp 1607721120
transform 1 0 4600 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_53
timestamp 1607721120
transform 1 0 5980 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607721120
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1162_
timestamp 1607721120
transform 1 0 5336 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0649_
timestamp 1607721120
transform 1 0 6808 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_74
timestamp 1607721120
transform 1 0 7912 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_66
timestamp 1607721120
transform 1 0 7176 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1165_
timestamp 1607721120
transform 1 0 8004 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_101
timestamp 1607721120
transform 1 0 10396 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_84
timestamp 1607721120
transform 1 0 8832 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1193_
timestamp 1607721120
transform 1 0 9568 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_114
timestamp 1607721120
transform 1 0 11592 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_109
timestamp 1607721120
transform 1 0 11132 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607721120
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0900_
timestamp 1607721120
transform 1 0 12420 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1607721120
transform 1 0 11224 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_135
timestamp 1607721120
transform 1 0 13524 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_127
timestamp 1607721120
transform 1 0 12788 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1256_
timestamp 1607721120
transform 1 0 13708 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_45_156
timestamp 1607721120
transform 1 0 15456 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0750_
timestamp 1607721120
transform 1 0 16192 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_45_187
timestamp 1607721120
transform 1 0 18308 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1607721120
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607721120
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1607721120
transform 1 0 18032 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_199
timestamp 1607721120
transform 1 0 19412 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_223
timestamp 1607721120
transform 1 0 21620 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_211
timestamp 1607721120
transform 1 0 20516 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1607721120
transform 1 0 23644 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1607721120
transform 1 0 23460 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_235
timestamp 1607721120
transform 1 0 22724 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607721120
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_253
timestamp 1607721120
transform 1 0 24380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607721120
transform -1 0 24840 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_8
timestamp 1607721120
transform 1 0 1840 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1607721120
transform 1 0 1380 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607721120
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607721120
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607721120
transform 1 0 1380 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1192_
timestamp 1607721120
transform 1 0 2576 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1607721120
transform 1 0 1564 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_34
timestamp 1607721120
transform 1 0 4232 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_22
timestamp 1607721120
transform 1 0 3128 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_23
timestamp 1607721120
transform 1 0 3220 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607721120
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1051_
timestamp 1607721120
transform 1 0 4048 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0991_
timestamp 1607721120
transform 1 0 4508 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_47_62
timestamp 1607721120
transform 1 0 6808 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1607721120
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1607721120
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_48
timestamp 1607721120
transform 1 0 5520 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607721120
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1101_
timestamp 1607721120
transform 1 0 6256 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1607721120
transform 1 0 8280 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_68
timestamp 1607721120
transform 1 0 7360 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_72
timestamp 1607721120
transform 1 0 7728 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1163_
timestamp 1607721120
transform 1 0 7452 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0636_
timestamp 1607721120
transform 1 0 8464 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_95
timestamp 1607721120
transform 1 0 9844 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_102
timestamp 1607721120
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_84
timestamp 1607721120
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607721120
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1195_
timestamp 1607721120
transform 1 0 10580 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1194_
timestamp 1607721120
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1164_
timestamp 1607721120
transform 1 0 9016 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1607721120
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_112
timestamp 1607721120
transform 1 0 11408 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1607721120
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607721120
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1182_
timestamp 1607721120
transform 1 0 11224 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1076_
timestamp 1607721120
transform 1 0 12420 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_135
timestamp 1607721120
transform 1 0 13524 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_127
timestamp 1607721120
transform 1 0 12788 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_145
timestamp 1607721120
transform 1 0 14444 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_129
timestamp 1607721120
transform 1 0 12972 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1255_
timestamp 1607721120
transform 1 0 13616 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _0893_
timestamp 1607721120
transform 1 0 13156 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_47_163
timestamp 1607721120
transform 1 0 16100 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_155
timestamp 1607721120
transform 1 0 15364 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607721120
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607721120
transform 1 0 15272 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0748_
timestamp 1607721120
transform 1 0 16192 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_47_187
timestamp 1607721120
transform 1 0 18308 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1607721120
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_184
timestamp 1607721120
transform 1 0 18032 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_173
timestamp 1607721120
transform 1 0 17020 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607721120
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1607721120
transform 1 0 18032 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1607721120
transform 1 0 17756 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_199
timestamp 1607721120
transform 1 0 19412 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1607721120
transform 1 0 20240 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_196
timestamp 1607721120
transform 1 0 19136 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_223
timestamp 1607721120
transform 1 0 21620 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_211
timestamp 1607721120
transform 1 0 20516 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_227
timestamp 1607721120
transform 1 0 21988 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1607721120
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607721120
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_245
timestamp 1607721120
transform 1 0 23644 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_243
timestamp 1607721120
transform 1 0 23460 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_235
timestamp 1607721120
transform 1 0 22724 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_239
timestamp 1607721120
transform 1 0 23092 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607721120
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_253
timestamp 1607721120
transform 1 0 24380 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_251
timestamp 1607721120
transform 1 0 24196 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607721120
transform -1 0 24840 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607721120
transform -1 0 24840 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_11
timestamp 1607721120
transform 1 0 2116 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1607721120
transform 1 0 1748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1607721120
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607721120
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1050_
timestamp 1607721120
transform 1 0 2852 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1607721120
transform 1 0 1840 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_32
timestamp 1607721120
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_23
timestamp 1607721120
transform 1 0 3220 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607721120
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0667_
timestamp 1607721120
transform 1 0 4232 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_43
timestamp 1607721120
transform 1 0 5060 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1240_
timestamp 1607721120
transform 1 0 5796 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_48_82
timestamp 1607721120
transform 1 0 8648 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_70
timestamp 1607721120
transform 1 0 7544 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0960_
timestamp 1607721120
transform 1 0 8280 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1607721120
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_90
timestamp 1607721120
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607721120
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1222_
timestamp 1607721120
transform 1 0 10028 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_48_116
timestamp 1607721120
transform 1 0 11776 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1078_
timestamp 1607721120
transform 1 0 12512 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_140
timestamp 1607721120
transform 1 0 13984 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_154
timestamp 1607721120
transform 1 0 15272 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_152
timestamp 1607721120
transform 1 0 15088 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607721120
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0751_
timestamp 1607721120
transform 1 0 15456 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_48_181
timestamp 1607721120
transform 1 0 17756 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_170
timestamp 1607721120
transform 1 0 16744 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1607721120
transform 1 0 17480 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_205
timestamp 1607721120
transform 1 0 19964 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_193
timestamp 1607721120
transform 1 0 18860 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1607721120
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1607721120
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1607721120
transform 1 0 20700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607721120
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1607721120
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_251
timestamp 1607721120
transform 1 0 24196 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607721120
transform -1 0 24840 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607721120
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1271_
timestamp 1607721120
transform 1 0 1380 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_22
timestamp 1607721120
transform 1 0 3128 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1052_
timestamp 1607721120
transform 1 0 3864 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_49_58
timestamp 1607721120
transform 1 0 6440 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_46
timestamp 1607721120
transform 1 0 5336 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607721120
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1102_
timestamp 1607721120
transform 1 0 6808 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_49_78
timestamp 1607721120
transform 1 0 8280 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_90
timestamp 1607721120
transform 1 0 9384 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1126_
timestamp 1607721120
transform 1 0 10120 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1607721120
transform 1 0 9016 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_123
timestamp 1607721120
transform 1 0 12420 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_114
timestamp 1607721120
transform 1 0 11592 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607721120
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_145
timestamp 1607721120
transform 1 0 14444 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1254_
timestamp 1607721120
transform 1 0 12696 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_162
timestamp 1607721120
transform 1 0 16008 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0744_
timestamp 1607721120
transform 1 0 15180 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_49_187
timestamp 1607721120
transform 1 0 18308 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1607721120
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_173
timestamp 1607721120
transform 1 0 17020 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607721120
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1607721120
transform 1 0 18032 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1607721120
transform 1 0 16744 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_199
timestamp 1607721120
transform 1 0 19412 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_223
timestamp 1607721120
transform 1 0 21620 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_211
timestamp 1607721120
transform 1 0 20516 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_245
timestamp 1607721120
transform 1 0 23644 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_243
timestamp 1607721120
transform 1 0 23460 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_235
timestamp 1607721120
transform 1 0 22724 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607721120
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_253
timestamp 1607721120
transform 1 0 24380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607721120
transform -1 0 24840 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607721120
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1270_
timestamp 1607721120
transform 1 0 1380 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_50_38
timestamp 1607721120
transform 1 0 4600 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_32
timestamp 1607721120
transform 1 0 4048 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1607721120
transform 1 0 3864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_22
timestamp 1607721120
transform 1 0 3128 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607721120
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0990_
timestamp 1607721120
transform 1 0 4692 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_43
timestamp 1607721120
transform 1 0 5060 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1239_
timestamp 1607721120
transform 1 0 5796 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_50_78
timestamp 1607721120
transform 1 0 8280 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_70
timestamp 1607721120
transform 1 0 7544 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1151_
timestamp 1607721120
transform 1 0 8464 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_102
timestamp 1607721120
transform 1 0 10488 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_84
timestamp 1607721120
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607721120
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1190_
timestamp 1607721120
transform 1 0 9660 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_50_110
timestamp 1607721120
transform 1 0 11224 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1080_
timestamp 1607721120
transform 1 0 11500 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_144
timestamp 1607721120
transform 1 0 14352 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_129
timestamp 1607721120
transform 1 0 12972 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1189_
timestamp 1607721120
transform 1 0 13708 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_50_152
timestamp 1607721120
transform 1 0 15088 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607721120
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607721120
transform 1 0 15272 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_185
timestamp 1607721120
transform 1 0 18124 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_173
timestamp 1607721120
transform 1 0 17020 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1607721120
transform 1 0 19228 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607721120
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607721120
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1607721120
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1607721120
transform 1 0 20332 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607721120
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_239
timestamp 1607721120
transform 1 0 23092 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_251
timestamp 1607721120
transform 1 0 24196 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607721120
transform -1 0 24840 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_12
timestamp 1607721120
transform 1 0 2208 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1607721120
transform 1 0 1380 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607721120
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1054_
timestamp 1607721120
transform 1 0 2944 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1607721120
transform 1 0 1932 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_36
timestamp 1607721120
transform 1 0 4416 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_53
timestamp 1607721120
transform 1 0 5980 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_44
timestamp 1607721120
transform 1 0 5152 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607721120
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1161_
timestamp 1607721120
transform 1 0 5336 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1607721120
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_83
timestamp 1607721120
transform 1 0 8740 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_73
timestamp 1607721120
transform 1 0 7820 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_65
timestamp 1607721120
transform 1 0 7084 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1160_
timestamp 1607721120
transform 1 0 7912 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_99
timestamp 1607721120
transform 1 0 10212 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 1607721120
transform 1 0 9844 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0901_
timestamp 1607721120
transform 1 0 10304 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_51_114
timestamp 1607721120
transform 1 0 11592 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607721120
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0745_
timestamp 1607721120
transform 1 0 12420 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_51_136
timestamp 1607721120
transform 1 0 13616 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_148
timestamp 1607721120
transform 1 0 14720 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _0752_
timestamp 1607721120
transform 1 0 15272 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1607721120
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_180
timestamp 1607721120
transform 1 0 17664 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_168
timestamp 1607721120
transform 1 0 16560 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607721120
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1607721120
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1607721120
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_220
timestamp 1607721120
transform 1 0 21344 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_245
timestamp 1607721120
transform 1 0 23644 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1607721120
transform 1 0 22448 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607721120
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_253
timestamp 1607721120
transform 1 0 24380 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607721120
transform -1 0 24840 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_3
timestamp 1607721120
transform 1 0 1380 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_11
timestamp 1607721120
transform 1 0 2116 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1607721120
transform 1 0 1748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1607721120
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607721120
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607721120
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1268_
timestamp 1607721120
transform 1 0 1472 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1607721120
transform 1 0 2852 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1607721120
transform 1 0 1840 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_23
timestamp 1607721120
transform 1 0 3220 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_40
timestamp 1607721120
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_32
timestamp 1607721120
transform 1 0 4048 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_23
timestamp 1607721120
transform 1 0 3220 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607721120
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1056_
timestamp 1607721120
transform 1 0 3956 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_53_62
timestamp 1607721120
transform 1 0 6808 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_59
timestamp 1607721120
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_47
timestamp 1607721120
transform 1 0 5428 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_58
timestamp 1607721120
transform 1 0 6440 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607721120
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1104_
timestamp 1607721120
transform 1 0 4968 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_53_68
timestamp 1607721120
transform 1 0 7360 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_76
timestamp 1607721120
transform 1 0 8096 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_wb_clk_i
timestamp 1607721120
transform 1 0 7176 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1607721120
transform 1 0 8096 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1149_
timestamp 1607721120
transform 1 0 7452 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1607721120
transform 1 0 7084 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_95
timestamp 1607721120
transform 1 0 9844 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_93
timestamp 1607721120
transform 1 0 9660 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_88
timestamp 1607721120
transform 1 0 9200 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607721120
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1159_
timestamp 1607721120
transform 1 0 10580 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1127_
timestamp 1607721120
transform 1 0 9752 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_53_121
timestamp 1607721120
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_110
timestamp 1607721120
transform 1 0 11224 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_110
timestamp 1607721120
transform 1 0 11224 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_wb_clk_i
timestamp 1607721120
transform 1 0 11960 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607721120
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1253_
timestamp 1607721120
transform 1 0 12420 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _0906_
timestamp 1607721120
transform 1 0 11960 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_53_142
timestamp 1607721120
transform 1 0 14168 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_143
timestamp 1607721120
transform 1 0 14260 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1607721120
transform 1 0 13248 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1607721120
transform 1 0 13984 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_166
timestamp 1607721120
transform 1 0 16376 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_150
timestamp 1607721120
transform 1 0 14904 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_163
timestamp 1607721120
transform 1 0 16100 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_151
timestamp 1607721120
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607721120
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1139_
timestamp 1607721120
transform 1 0 15272 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0754_
timestamp 1607721120
transform 1 0 15088 0 1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1607721120
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1607721120
transform 1 0 17848 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_178
timestamp 1607721120
transform 1 0 17480 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_186
timestamp 1607721120
transform 1 0 18216 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_174
timestamp 1607721120
transform 1 0 17112 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607721120
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1607721120
transform 1 0 16836 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1607721120
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1607721120
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_198
timestamp 1607721120
transform 1 0 19320 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_220
timestamp 1607721120
transform 1 0 21344 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607721120
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607721120
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1607721120
transform 1 0 20424 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607721120
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_245
timestamp 1607721120
transform 1 0 23644 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_232
timestamp 1607721120
transform 1 0 22448 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1607721120
transform 1 0 23092 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607721120
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_253
timestamp 1607721120
transform 1 0 24380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_251
timestamp 1607721120
transform 1 0 24196 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607721120
transform -1 0 24840 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607721120
transform -1 0 24840 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_12
timestamp 1607721120
transform 1 0 2208 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1607721120
transform 1 0 1380 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607721120
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1607721120
transform 1 0 1932 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1607721120
transform 1 0 2944 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_32
timestamp 1607721120
transform 1 0 4048 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_23
timestamp 1607721120
transform 1 0 3220 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607721120
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1100_
timestamp 1607721120
transform 1 0 4784 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_44
timestamp 1607721120
transform 1 0 5152 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1238_
timestamp 1607721120
transform 1 0 5888 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_54_79
timestamp 1607721120
transform 1 0 8372 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_71
timestamp 1607721120
transform 1 0 7636 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1125_
timestamp 1607721120
transform 1 0 8464 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_100
timestamp 1607721120
transform 1 0 10304 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_84
timestamp 1607721120
transform 1 0 8832 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607721120
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1158_
timestamp 1607721120
transform 1 0 9660 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_54_125
timestamp 1607721120
transform 1 0 12604 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_108
timestamp 1607721120
transform 1 0 11040 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1081_
timestamp 1607721120
transform 1 0 11132 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_54_145
timestamp 1607721120
transform 1 0 14444 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_wb_clk_i
timestamp 1607721120
transform 1 0 13340 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0746_
timestamp 1607721120
transform 1 0 13616 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607721120
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1330_
timestamp 1607721120
transform 1 0 15272 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_54_184
timestamp 1607721120
transform 1 0 18032 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_173
timestamp 1607721120
transform 1 0 17020 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1607721120
transform 1 0 17756 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_208
timestamp 1607721120
transform 1 0 20240 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_196
timestamp 1607721120
transform 1 0 19136 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1607721120
transform 1 0 21988 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1607721120
transform 1 0 20884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607721120
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_239
timestamp 1607721120
transform 1 0 23092 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_251
timestamp 1607721120
transform 1 0 24196 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607721120
transform -1 0 24840 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1607721120
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1607721120
transform 1 0 1380 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607721120
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1607721120
transform 1 0 1472 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1055_
timestamp 1607721120
transform 1 0 2852 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_55_35
timestamp 1607721120
transform 1 0 4324 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_62
timestamp 1607721120
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_58
timestamp 1607721120
transform 1 0 6440 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1607721120
transform 1 0 5428 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_wb_clk_i
timestamp 1607721120
transform 1 0 6164 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607721120
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1103_
timestamp 1607721120
transform 1 0 5060 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_80
timestamp 1607721120
transform 1 0 8464 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0931_
timestamp 1607721120
transform 1 0 7176 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__dfxtp_4  _1220_
timestamp 1607721120
transform 1 0 9200 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_55_119
timestamp 1607721120
transform 1 0 12052 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_107
timestamp 1607721120
transform 1 0 10948 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607721120
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1079_
timestamp 1607721120
transform 1 0 12420 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_135
timestamp 1607721120
transform 1 0 13524 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_127
timestamp 1607721120
transform 1 0 12788 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1329_
timestamp 1607721120
transform 1 0 13616 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_55_155
timestamp 1607721120
transform 1 0 15364 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0747_
timestamp 1607721120
transform 1 0 16100 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1607721120
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_182
timestamp 1607721120
transform 1 0 17848 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_170
timestamp 1607721120
transform 1 0 16744 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607721120
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1607721120
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1607721120
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_220
timestamp 1607721120
transform 1 0 21344 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_245
timestamp 1607721120
transform 1 0 23644 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1607721120
transform 1 0 22448 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607721120
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_253
timestamp 1607721120
transform 1 0 24380 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607721120
transform -1 0 24840 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_12
timestamp 1607721120
transform 1 0 2208 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1607721120
transform 1 0 1380 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607721120
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1607721120
transform 1 0 1932 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1607721120
transform 1 0 2944 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_35
timestamp 1607721120
transform 1 0 4324 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_23
timestamp 1607721120
transform 1 0 3220 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607721120
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1607721120
transform 1 0 4048 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_47
timestamp 1607721120
transform 1 0 5428 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1607721120
transform 1 0 5704 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1237_
timestamp 1607721120
transform 1 0 5980 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_80
timestamp 1607721120
transform 1 0 8464 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_72
timestamp 1607721120
transform 1 0 7728 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1607721120
transform 1 0 8556 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_100
timestamp 1607721120
transform 1 0 10304 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_84
timestamp 1607721120
transform 1 0 8832 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607721120
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1188_
timestamp 1607721120
transform 1 0 9660 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_56_125
timestamp 1607721120
transform 1 0 12604 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_108
timestamp 1607721120
transform 1 0 11040 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1082_
timestamp 1607721120
transform 1 0 11132 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_145
timestamp 1607721120
transform 1 0 14444 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1607721120
transform 1 0 13340 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1140_
timestamp 1607721120
transform 1 0 13616 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607721120
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0758_
timestamp 1607721120
transform 1 0 15272 0 -1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1607721120
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1607721120
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_204
timestamp 1607721120
transform 1 0 19872 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_192
timestamp 1607721120
transform 1 0 18768 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_227
timestamp 1607721120
transform 1 0 21988 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1607721120
transform 1 0 20884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_212
timestamp 1607721120
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607721120
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1607721120
transform 1 0 23092 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_251
timestamp 1607721120
transform 1 0 24196 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607721120
transform -1 0 24840 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_11
timestamp 1607721120
transform 1 0 2116 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_3
timestamp 1607721120
transform 1 0 1380 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607721120
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1269_
timestamp 1607721120
transform 1 0 2208 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_31
timestamp 1607721120
transform 1 0 3956 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0996_
timestamp 1607721120
transform 1 0 4692 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_57_62
timestamp 1607721120
transform 1 0 6808 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_53
timestamp 1607721120
transform 1 0 5980 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607721120
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_68
timestamp 1607721120
transform 1 0 7360 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1217_
timestamp 1607721120
transform 1 0 7452 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_88
timestamp 1607721120
transform 1 0 9200 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1128_
timestamp 1607721120
transform 1 0 9936 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_57_120
timestamp 1607721120
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_112
timestamp 1607721120
transform 1 0 11408 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607721120
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1252_
timestamp 1607721120
transform 1 0 12420 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_142
timestamp 1607721120
transform 1 0 14168 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_161
timestamp 1607721120
transform 1 0 15916 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_153
timestamp 1607721120
transform 1 0 15180 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0842_
timestamp 1607721120
transform 1 0 16008 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1607721120
transform 1 0 14904 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1607721120
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_171
timestamp 1607721120
transform 1 0 16836 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607721120
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1607721120
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1607721120
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_220
timestamp 1607721120
transform 1 0 21344 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_245
timestamp 1607721120
transform 1 0 23644 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_232
timestamp 1607721120
transform 1 0 22448 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607721120
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_253
timestamp 1607721120
transform 1 0 24380 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607721120
transform -1 0 24840 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1607721120
transform 1 0 1380 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607721120
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _1007_
timestamp 1607721120
transform 1 0 1932 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_58_32
timestamp 1607721120
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_23
timestamp 1607721120
transform 1 0 3220 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607721120
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1607721120
transform 1 0 4784 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_43
timestamp 1607721120
transform 1 0 5060 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1236_
timestamp 1607721120
transform 1 0 5796 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_58_82
timestamp 1607721120
transform 1 0 8648 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_70
timestamp 1607721120
transform 1 0 7544 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1129_
timestamp 1607721120
transform 1 0 8280 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_98
timestamp 1607721120
transform 1 0 10120 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1607721120
transform 1 0 9660 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_90
timestamp 1607721120
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607721120
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1607721120
transform 1 0 9752 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1607721120
transform 1 0 12236 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_106
timestamp 1607721120
transform 1 0 10856 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0912_
timestamp 1607721120
transform 1 0 10948 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_58_145
timestamp 1607721120
transform 1 0 14444 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_132
timestamp 1607721120
transform 1 0 13248 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 12972 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 13616 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_58_166
timestamp 1607721120
transform 1 0 16376 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_154
timestamp 1607721120
transform 1 0 15272 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607721120
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_187
timestamp 1607721120
transform 1 0 18308 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1315_
timestamp 1607721120
transform 1 0 16560 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_199
timestamp 1607721120
transform 1 0 19412 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1607721120
transform 1 0 21988 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1607721120
transform 1 0 20884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_211
timestamp 1607721120
transform 1 0 20516 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607721120
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1607721120
transform 1 0 23092 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_251
timestamp 1607721120
transform 1 0 24196 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607721120
transform -1 0 24840 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607721120
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607721120
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607721120
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607721120
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607721120
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _1002_
timestamp 1607721120
transform 1 0 2484 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 1607721120
transform 1 0 4876 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607721120
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_29
timestamp 1607721120
transform 1 0 3772 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607721120
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1105_
timestamp 1607721120
transform 1 0 4508 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_4  _1018_
timestamp 1607721120
transform 1 0 4048 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_59_53
timestamp 1607721120
transform 1 0 5980 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607721120
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1282_
timestamp 1607721120
transform 1 0 5612 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1132_
timestamp 1607721120
transform 1 0 6808 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_83
timestamp 1607721120
transform 1 0 8740 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_68
timestamp 1607721120
transform 1 0 7360 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_78
timestamp 1607721120
transform 1 0 8280 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1030_
timestamp 1607721120
transform 1 0 8096 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_60_93
timestamp 1607721120
transform 1 0 9660 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_91
timestamp 1607721120
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_102
timestamp 1607721120
transform 1 0 10488 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607721120
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1249_
timestamp 1607721120
transform 1 0 9936 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1086_
timestamp 1607721120
transform 1 0 9016 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_123
timestamp 1607721120
transform 1 0 12420 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_115
timestamp 1607721120
transform 1 0 11684 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_114
timestamp 1607721120
transform 1 0 11592 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_110
timestamp 1607721120
transform 1 0 11224 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607721120
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0739_
timestamp 1607721120
transform 1 0 12420 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1607721120
transform 1 0 11316 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1607721120
transform 1 0 12512 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_145
timestamp 1607721120
transform 1 0 14444 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_128
timestamp 1607721120
transform 1 0 12880 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_143
timestamp 1607721120
transform 1 0 14260 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_132
timestamp 1607721120
transform 1 0 13248 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0759_
timestamp 1607721120
transform 1 0 13616 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1607721120
transform 1 0 13984 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_165
timestamp 1607721120
transform 1 0 16284 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_157
timestamp 1607721120
transform 1 0 15548 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_162
timestamp 1607721120
transform 1 0 16008 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_151
timestamp 1607721120
transform 1 0 14996 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607721120
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0841_
timestamp 1607721120
transform 1 0 15180 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1607721120
transform 1 0 15272 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_187
timestamp 1607721120
transform 1 0 18308 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_182
timestamp 1607721120
transform 1 0 17848 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_174
timestamp 1607721120
transform 1 0 17112 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607721120
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1314_
timestamp 1607721120
transform 1 0 16560 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _0847_
timestamp 1607721120
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_199
timestamp 1607721120
transform 1 0 19412 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1607721120
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1607721120
transform 1 0 18860 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0843_
timestamp 1607721120
transform 1 0 19596 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1607721120
transform 1 0 21988 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1607721120
transform 1 0 20884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_211
timestamp 1607721120
transform 1 0 20516 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_220
timestamp 1607721120
transform 1 0 21344 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607721120
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1607721120
transform 1 0 23092 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_245
timestamp 1607721120
transform 1 0 23644 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_232
timestamp 1607721120
transform 1 0 22448 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607721120
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_251
timestamp 1607721120
transform 1 0 24196 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_253
timestamp 1607721120
transform 1 0 24380 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607721120
transform -1 0 24840 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607721120
transform -1 0 24840 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_15
timestamp 1607721120
transform 1 0 2484 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607721120
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607721120
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_29
timestamp 1607721120
transform 1 0 3772 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_23
timestamp 1607721120
transform 1 0 3220 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1106_
timestamp 1607721120
transform 1 0 4508 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1607721120
transform 1 0 3496 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_53
timestamp 1607721120
transform 1 0 5980 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607721120
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1607721120
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_74
timestamp 1607721120
transform 1 0 7912 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_66
timestamp 1607721120
transform 1 0 7176 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1131_
timestamp 1607721120
transform 1 0 8004 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_61_103
timestamp 1607721120
transform 1 0 10580 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_99
timestamp 1607721120
transform 1 0 10212 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_91
timestamp 1607721120
transform 1 0 9476 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1607721120
transform 1 0 10304 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_114
timestamp 1607721120
transform 1 0 11592 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607721120
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1325_
timestamp 1607721120
transform 1 0 12420 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1607721120
transform 1 0 11316 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_142
timestamp 1607721120
transform 1 0 14168 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1328_
timestamp 1607721120
transform 1 0 14904 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_61_181
timestamp 1607721120
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1607721120
transform 1 0 16652 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607721120
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0831_
timestamp 1607721120
transform 1 0 18032 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_61_203
timestamp 1607721120
transform 1 0 19780 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_191
timestamp 1607721120
transform 1 0 18676 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_227
timestamp 1607721120
transform 1 0 21988 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_215
timestamp 1607721120
transform 1 0 20884 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_245
timestamp 1607721120
transform 1 0 23644 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1607721120
transform 1 0 23460 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1607721120
transform 1 0 23092 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607721120
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_253
timestamp 1607721120
transform 1 0 24380 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607721120
transform -1 0 24840 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_19
timestamp 1607721120
transform 1 0 2852 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1607721120
transform 1 0 2484 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607721120
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607721120
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1607721120
transform 1 0 2944 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1607721120
transform 1 0 4048 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_23
timestamp 1607721120
transform 1 0 3220 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607721120
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1025_
timestamp 1607721120
transform 1 0 4600 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_62_55
timestamp 1607721120
transform 1 0 6164 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_63
timestamp 1607721120
transform 1 0 6900 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1218_
timestamp 1607721120
transform 1 0 7084 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_99
timestamp 1607721120
transform 1 0 10212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_93
timestamp 1607721120
transform 1 0 9660 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_84
timestamp 1607721120
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607721120
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0923_
timestamp 1607721120
transform 1 0 10304 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_62_114
timestamp 1607721120
transform 1 0 11592 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0769_
timestamp 1607721120
transform 1 0 12328 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_136
timestamp 1607721120
transform 1 0 13616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_163
timestamp 1607721120
transform 1 0 16100 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1607721120
transform 1 0 15088 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_148
timestamp 1607721120
transform 1 0 14720 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607721120
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0734_
timestamp 1607721120
transform 1 0 15272 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_178
timestamp 1607721120
transform 1 0 17480 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0756_
timestamp 1607721120
transform 1 0 16836 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_202
timestamp 1607721120
transform 1 0 19688 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_190
timestamp 1607721120
transform 1 0 18584 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1607721120
transform 1 0 21988 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1607721120
transform 1 0 20884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607721120
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1607721120
transform 1 0 23092 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_251
timestamp 1607721120
transform 1 0 24196 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607721120
transform -1 0 24840 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_15
timestamp 1607721120
transform 1 0 2484 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607721120
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607721120
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1285_
timestamp 1607721120
transform 1 0 2760 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_63_37
timestamp 1607721120
transform 1 0 4508 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_60
timestamp 1607721120
transform 1 0 6624 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_52
timestamp 1607721120
transform 1 0 5888 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607721120
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1026_
timestamp 1607721120
transform 1 0 6808 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1015_
timestamp 1607721120
transform 1 0 5244 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_63_81
timestamp 1607721120
transform 1 0 8556 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1607721120
transform 1 0 7452 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0830_
timestamp 1607721120
transform 1 0 8188 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 9292 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1085_
timestamp 1607721120
transform 1 0 9568 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_63_123
timestamp 1607721120
transform 1 0 12420 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_119
timestamp 1607721120
transform 1 0 12052 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_108
timestamp 1607721120
transform 1 0 11040 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 11776 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607721120
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0755_
timestamp 1607721120
transform 1 0 12604 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_63_132
timestamp 1607721120
transform 1 0 13248 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0762_
timestamp 1607721120
transform 1 0 13984 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_63_154
timestamp 1607721120
transform 1 0 15272 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0853_
timestamp 1607721120
transform 1 0 16008 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1607721120
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_171
timestamp 1607721120
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607721120
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1607721120
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1607721120
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_220
timestamp 1607721120
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_245
timestamp 1607721120
transform 1 0 23644 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_232
timestamp 1607721120
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607721120
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_253
timestamp 1607721120
transform 1 0 24380 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607721120
transform -1 0 24840 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_11
timestamp 1607721120
transform 1 0 2116 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_3
timestamp 1607721120
transform 1 0 1380 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607721120
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _1019_
timestamp 1607721120
transform 1 0 2392 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_64_38
timestamp 1607721120
transform 1 0 4600 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_32
timestamp 1607721120
transform 1 0 4048 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_23
timestamp 1607721120
transform 1 0 3220 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607721120
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1284_
timestamp 1607721120
transform 1 0 4692 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_58
timestamp 1607721120
transform 1 0 6440 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_66
timestamp 1607721120
transform 1 0 7176 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1130_
timestamp 1607721120
transform 1 0 7360 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1607721120
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_84
timestamp 1607721120
transform 1 0 8832 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607721120
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1084_
timestamp 1607721120
transform 1 0 9752 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_110
timestamp 1607721120
transform 1 0 11224 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0918_
timestamp 1607721120
transform 1 0 11960 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_64_143
timestamp 1607721120
transform 1 0 14260 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1607721120
transform 1 0 13248 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1607721120
transform 1 0 13984 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_166
timestamp 1607721120
transform 1 0 16376 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_158
timestamp 1607721120
transform 1 0 15640 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_151
timestamp 1607721120
transform 1 0 14996 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607721120
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0867_
timestamp 1607721120
transform 1 0 15272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_186
timestamp 1607721120
transform 1 0 18216 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1313_
timestamp 1607721120
transform 1 0 16468 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_198
timestamp 1607721120
transform 1 0 19320 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_227
timestamp 1607721120
transform 1 0 21988 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1607721120
transform 1 0 20884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1607721120
transform 1 0 20424 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607721120
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1607721120
transform 1 0 23092 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_251
timestamp 1607721120
transform 1 0 24196 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607721120
transform -1 0 24840 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_15
timestamp 1607721120
transform 1 0 2484 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607721120
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607721120
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1607721120
transform 1 0 2852 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_39
timestamp 1607721120
transform 1 0 4692 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_22
timestamp 1607721120
transform 1 0 3128 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1013_
timestamp 1607721120
transform 1 0 3864 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_65_53
timestamp 1607721120
transform 1 0 5980 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_47
timestamp 1607721120
transform 1 0 5428 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607721120
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0973_
timestamp 1607721120
transform 1 0 6808 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0848_
timestamp 1607721120
transform 1 0 5612 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_79
timestamp 1607721120
transform 1 0 8372 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_71
timestamp 1607721120
transform 1 0 7636 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1219_
timestamp 1607721120
transform 1 0 8464 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_99
timestamp 1607721120
transform 1 0 10212 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_123
timestamp 1607721120
transform 1 0 12420 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_114
timestamp 1607721120
transform 1 0 11592 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1607721120
transform 1 0 10948 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607721120
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607721120
transform 1 0 11224 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_142
timestamp 1607721120
transform 1 0 14168 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_127
timestamp 1607721120
transform 1 0 12788 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0765_
timestamp 1607721120
transform 1 0 12880 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_65_154
timestamp 1607721120
transform 1 0 15272 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0854_
timestamp 1607721120
transform 1 0 16008 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0833_
timestamp 1607721120
transform 1 0 14904 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_187
timestamp 1607721120
transform 1 0 18308 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_171
timestamp 1607721120
transform 1 0 16836 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607721120
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1607721120
transform 1 0 18032 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_199
timestamp 1607721120
transform 1 0 19412 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_223
timestamp 1607721120
transform 1 0 21620 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_211
timestamp 1607721120
transform 1 0 20516 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_245
timestamp 1607721120
transform 1 0 23644 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1607721120
transform 1 0 23460 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_235
timestamp 1607721120
transform 1 0 22724 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607721120
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_253
timestamp 1607721120
transform 1 0 24380 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607721120
transform -1 0 24840 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_19
timestamp 1607721120
transform 1 0 2852 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_9
timestamp 1607721120
transform 1 0 1932 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1607721120
transform 1 0 1380 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_15
timestamp 1607721120
transform 1 0 2484 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1607721120
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607721120
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607721120
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _1014_
timestamp 1607721120
transform 1 0 2024 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0957_
timestamp 1607721120
transform 1 0 2852 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_36
timestamp 1607721120
transform 1 0 4416 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_39
timestamp 1607721120
transform 1 0 4692 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_23
timestamp 1607721120
transform 1 0 3220 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607721120
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1010_
timestamp 1607721120
transform 1 0 4048 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1008_
timestamp 1607721120
transform 1 0 3588 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_67_62
timestamp 1607721120
transform 1 0 6808 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_53
timestamp 1607721120
transform 1 0 5980 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_57
timestamp 1607721120
transform 1 0 6348 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_47
timestamp 1607721120
transform 1 0 5428 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607721120
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0984_
timestamp 1607721120
transform 1 0 5152 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0979_
timestamp 1607721120
transform 1 0 5520 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_67_74
timestamp 1607721120
transform 1 0 7912 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_74
timestamp 1607721120
transform 1 0 7912 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1607721120
transform 1 0 8648 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0967_
timestamp 1607721120
transform 1 0 7084 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0962_
timestamp 1607721120
transform 1 0 7084 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0832_
timestamp 1607721120
transform 1 0 8648 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_103
timestamp 1607721120
transform 1 0 10580 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_86
timestamp 1607721120
transform 1 0 9016 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_97
timestamp 1607721120
transform 1 0 10028 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_91
timestamp 1607721120
transform 1 0 9476 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_85
timestamp 1607721120
transform 1 0 8924 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607721120
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0937_
timestamp 1607721120
transform 1 0 9752 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1607721120
transform 1 0 9660 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_123
timestamp 1607721120
transform 1 0 12420 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_114
timestamp 1607721120
transform 1 0 11592 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_105
timestamp 1607721120
transform 1 0 10764 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607721120
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1327_
timestamp 1607721120
transform 1 0 12604 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1251_
timestamp 1607721120
transform 1 0 10948 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1607721120
transform 1 0 11316 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_144
timestamp 1607721120
transform 1 0 14352 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_145
timestamp 1607721120
transform 1 0 14444 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_134
timestamp 1607721120
transform 1 0 13432 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_126
timestamp 1607721120
transform 1 0 12696 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0889_
timestamp 1607721120
transform 1 0 13616 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_67_161
timestamp 1607721120
transform 1 0 15916 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_163
timestamp 1607721120
transform 1 0 16100 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607721120
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0864_
timestamp 1607721120
transform 1 0 15088 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0859_
timestamp 1607721120
transform 1 0 15272 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1607721120
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_181
timestamp 1607721120
transform 1 0 17756 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_173
timestamp 1607721120
transform 1 0 17020 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_178
timestamp 1607721120
transform 1 0 17480 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607721120
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1607721120
transform 1 0 16652 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0850_
timestamp 1607721120
transform 1 0 16836 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1607721120
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1607721120
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_202
timestamp 1607721120
transform 1 0 19688 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_190
timestamp 1607721120
transform 1 0 18584 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_220
timestamp 1607721120
transform 1 0 21344 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_227
timestamp 1607721120
transform 1 0 21988 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1607721120
transform 1 0 20884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607721120
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_245
timestamp 1607721120
transform 1 0 23644 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_232
timestamp 1607721120
transform 1 0 22448 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_239
timestamp 1607721120
transform 1 0 23092 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607721120
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_253
timestamp 1607721120
transform 1 0 24380 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_251
timestamp 1607721120
transform 1 0 24196 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607721120
transform -1 0 24840 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607721120
transform -1 0 24840 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1607721120
transform 1 0 2484 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607721120
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607721120
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0987_
timestamp 1607721120
transform 1 0 2852 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1607721120
transform 1 0 4048 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_23
timestamp 1607721120
transform 1 0 3220 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607721120
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0997_
timestamp 1607721120
transform 1 0 4416 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_62
timestamp 1607721120
transform 1 0 6808 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_45
timestamp 1607721120
transform 1 0 5244 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0828_
timestamp 1607721120
transform 1 0 5980 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_68_73
timestamp 1607721120
transform 1 0 7820 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_wb_clk_i
timestamp 1607721120
transform 1 0 7544 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0954_
timestamp 1607721120
transform 1 0 8004 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_101
timestamp 1607721120
transform 1 0 10396 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_93
timestamp 1607721120
transform 1 0 9660 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_84
timestamp 1607721120
transform 1 0 8832 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607721120
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1250_
timestamp 1607721120
transform 1 0 10488 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_68_121
timestamp 1607721120
transform 1 0 12236 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_145
timestamp 1607721120
transform 1 0 14444 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_132
timestamp 1607721120
transform 1 0 13248 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_wb_clk_i
timestamp 1607721120
transform 1 0 12972 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0883_
timestamp 1607721120
transform 1 0 13616 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_161
timestamp 1607721120
transform 1 0 15916 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607721120
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0763_
timestamp 1607721120
transform 1 0 15272 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_68_169
timestamp 1607721120
transform 1 0 16652 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1312_
timestamp 1607721120
transform 1 0 16744 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_201
timestamp 1607721120
transform 1 0 19596 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_189
timestamp 1607721120
transform 1 0 18492 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_227
timestamp 1607721120
transform 1 0 21988 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_215
timestamp 1607721120
transform 1 0 20884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_213
timestamp 1607721120
transform 1 0 20700 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607721120
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1607721120
transform 1 0 23092 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_251
timestamp 1607721120
transform 1 0 24196 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607721120
transform -1 0 24840 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_3
timestamp 1607721120
transform 1 0 1380 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607721120
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1286_
timestamp 1607721120
transform 1 0 2116 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_69_38
timestamp 1607721120
transform 1 0 4600 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_30
timestamp 1607721120
transform 1 0 3864 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0992_
timestamp 1607721120
transform 1 0 4784 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_62
timestamp 1607721120
transform 1 0 6808 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_60
timestamp 1607721120
transform 1 0 6624 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_49
timestamp 1607721120
transform 1 0 5612 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_wb_clk_i
timestamp 1607721120
transform 1 0 6348 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607721120
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_80
timestamp 1607721120
transform 1 0 8464 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_70
timestamp 1607721120
transform 1 0 7544 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0943_
timestamp 1607721120
transform 1 0 7636 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_97
timestamp 1607721120
transform 1 0 10028 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0932_
timestamp 1607721120
transform 1 0 9200 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_123
timestamp 1607721120
transform 1 0 12420 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_114
timestamp 1607721120
transform 1 0 11592 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607721120
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0919_
timestamp 1607721120
transform 1 0 10764 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_141
timestamp 1607721120
transform 1 0 14076 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0767_
timestamp 1607721120
transform 1 0 12788 0 1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_69_154
timestamp 1607721120
transform 1 0 15272 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_149
timestamp 1607721120
transform 1 0 14812 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0860_
timestamp 1607721120
transform 1 0 16008 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0849_
timestamp 1607721120
transform 1 0 14904 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_171
timestamp 1607721120
transform 1 0 16836 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607721120
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0856_
timestamp 1607721120
transform 1 0 18032 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_69_203
timestamp 1607721120
transform 1 0 19780 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_191
timestamp 1607721120
transform 1 0 18676 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_227
timestamp 1607721120
transform 1 0 21988 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_215
timestamp 1607721120
transform 1 0 20884 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_245
timestamp 1607721120
transform 1 0 23644 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_243
timestamp 1607721120
transform 1 0 23460 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_239
timestamp 1607721120
transform 1 0 23092 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607721120
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_253
timestamp 1607721120
transform 1 0 24380 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607721120
transform -1 0 24840 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_11
timestamp 1607721120
transform 1 0 2116 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1607721120
transform 1 0 1380 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607721120
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0999_
timestamp 1607721120
transform 1 0 1748 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0969_
timestamp 1607721120
transform 1 0 2852 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_32
timestamp 1607721120
transform 1 0 4048 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_23
timestamp 1607721120
transform 1 0 3220 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607721120
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1003_
timestamp 1607721120
transform 1 0 4416 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_70_57
timestamp 1607721120
transform 1 0 6348 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_45
timestamp 1607721120
transform 1 0 5244 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0974_
timestamp 1607721120
transform 1 0 6440 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_67
timestamp 1607721120
transform 1 0 7268 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0949_
timestamp 1607721120
transform 1 0 8004 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_99
timestamp 1607721120
transform 1 0 10212 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_93
timestamp 1607721120
transform 1 0 9660 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_84
timestamp 1607721120
transform 1 0 8832 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607721120
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0829_
timestamp 1607721120
transform 1 0 9844 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_116
timestamp 1607721120
transform 1 0 11776 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1326_
timestamp 1607721120
transform 1 0 12512 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _0902_
timestamp 1607721120
transform 1 0 10948 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_143
timestamp 1607721120
transform 1 0 14260 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_162
timestamp 1607721120
transform 1 0 16008 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_154
timestamp 1607721120
transform 1 0 15272 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1607721120
transform 1 0 14996 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607721120
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0861_
timestamp 1607721120
transform 1 0 15364 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1311_
timestamp 1607721120
transform 1 0 16744 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_201
timestamp 1607721120
transform 1 0 19596 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_189
timestamp 1607721120
transform 1 0 18492 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1607721120
transform 1 0 21988 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_215
timestamp 1607721120
transform 1 0 20884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_213
timestamp 1607721120
transform 1 0 20700 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607721120
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_239
timestamp 1607721120
transform 1 0 23092 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_251
timestamp 1607721120
transform 1 0 24196 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607721120
transform -1 0 24840 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_19
timestamp 1607721120
transform 1 0 2852 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_15
timestamp 1607721120
transform 1 0 2484 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607721120
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607721120
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _1009_
timestamp 1607721120
transform 1 0 2944 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_71_29
timestamp 1607721120
transform 1 0 3772 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1004_
timestamp 1607721120
transform 1 0 4508 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_71_62
timestamp 1607721120
transform 1 0 6808 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_58
timestamp 1607721120
transform 1 0 6440 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_46
timestamp 1607721120
transform 1 0 5336 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607721120
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_83
timestamp 1607721120
transform 1 0 8740 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1293_
timestamp 1607721120
transform 1 0 6992 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_71_97
timestamp 1607721120
transform 1 0 10028 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_91
timestamp 1607721120
transform 1 0 9476 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0885_
timestamp 1607721120
transform 1 0 9660 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_123
timestamp 1607721120
transform 1 0 12420 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_114
timestamp 1607721120
transform 1 0 11592 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607721120
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0913_
timestamp 1607721120
transform 1 0 10764 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_71_136
timestamp 1607721120
transform 1 0 13616 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0894_
timestamp 1607721120
transform 1 0 12788 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0872_
timestamp 1607721120
transform 1 0 14352 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_71_153
timestamp 1607721120
transform 1 0 15180 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0865_
timestamp 1607721120
transform 1 0 15916 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1607721120
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_182
timestamp 1607721120
transform 1 0 17848 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_170
timestamp 1607721120
transform 1 0 16744 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607721120
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_208
timestamp 1607721120
transform 1 0 20240 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_196
timestamp 1607721120
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_220
timestamp 1607721120
transform 1 0 21344 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_245
timestamp 1607721120
transform 1 0 23644 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_232
timestamp 1607721120
transform 1 0 22448 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607721120
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_253
timestamp 1607721120
transform 1 0 24380 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607721120
transform -1 0 24840 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_15
timestamp 1607721120
transform 1 0 2484 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607721120
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_15
timestamp 1607721120
transform 1 0 2484 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607721120
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607721120
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607721120
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1287_
timestamp 1607721120
transform 1 0 2668 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1000_
timestamp 1607721120
transform 1 0 2576 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_73_36
timestamp 1607721120
transform 1 0 4416 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_32
timestamp 1607721120
transform 1 0 4048 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_23
timestamp 1607721120
transform 1 0 3220 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607721120
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1288_
timestamp 1607721120
transform 1 0 4232 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_73_62
timestamp 1607721120
transform 1 0 6808 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_53
timestamp 1607721120
transform 1 0 5980 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1607721120
transform 1 0 5980 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607721120
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0985_
timestamp 1607721120
transform 1 0 5152 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_79
timestamp 1607721120
transform 1 0 8372 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_69
timestamp 1607721120
transform 1 0 7452 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1607721120
transform 1 0 7084 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1294_
timestamp 1607721120
transform 1 0 7544 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _0968_
timestamp 1607721120
transform 1 0 7544 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_73_101
timestamp 1607721120
transform 1 0 10396 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_89
timestamp 1607721120
transform 1 0 9292 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_102
timestamp 1607721120
transform 1 0 10488 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_91
timestamp 1607721120
transform 1 0 9476 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607721120
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0950_
timestamp 1607721120
transform 1 0 9660 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_73_123
timestamp 1607721120
transform 1 0 12420 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_114
timestamp 1607721120
transform 1 0 11592 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_123
timestamp 1607721120
transform 1 0 12420 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607721120
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0924_
timestamp 1607721120
transform 1 0 10764 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0907_
timestamp 1607721120
transform 1 0 11592 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_73_136
timestamp 1607721120
transform 1 0 13616 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_145
timestamp 1607721120
transform 1 0 14444 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_135
timestamp 1607721120
transform 1 0 13524 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_131
timestamp 1607721120
transform 1 0 13156 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_wb_clk_i
timestamp 1607721120
transform 1 0 13248 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0904_
timestamp 1607721120
transform 1 0 12972 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0878_
timestamp 1607721120
transform 1 0 14352 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0877_
timestamp 1607721120
transform 1 0 13616 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_73_153
timestamp 1607721120
transform 1 0 15180 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_162
timestamp 1607721120
transform 1 0 16008 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_154
timestamp 1607721120
transform 1 0 15272 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607721120
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0874_
timestamp 1607721120
transform 1 0 15364 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0873_
timestamp 1607721120
transform 1 0 15916 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_73_182
timestamp 1607721120
transform 1 0 17848 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_170
timestamp 1607721120
transform 1 0 16744 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607721120
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1310_
timestamp 1607721120
transform 1 0 16744 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0879_
timestamp 1607721120
transform 1 0 18032 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_200
timestamp 1607721120
transform 1 0 19504 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_188
timestamp 1607721120
transform 1 0 18400 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_201
timestamp 1607721120
transform 1 0 19596 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_189
timestamp 1607721120
transform 1 0 18492 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_224
timestamp 1607721120
transform 1 0 21712 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_212
timestamp 1607721120
transform 1 0 20608 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1607721120
transform 1 0 21988 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_215
timestamp 1607721120
transform 1 0 20884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_213
timestamp 1607721120
transform 1 0 20700 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607721120
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_245
timestamp 1607721120
transform 1 0 23644 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_236
timestamp 1607721120
transform 1 0 22816 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1607721120
transform 1 0 23092 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607721120
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_253
timestamp 1607721120
transform 1 0 24380 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_251
timestamp 1607721120
transform 1 0 24196 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607721120
transform -1 0 24840 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607721120
transform -1 0 24840 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_11
timestamp 1607721120
transform 1 0 2116 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1607721120
transform 1 0 1380 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607721120
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0975_
timestamp 1607721120
transform 1 0 1748 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1607721120
transform 1 0 2852 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_40
timestamp 1607721120
transform 1 0 4784 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_32
timestamp 1607721120
transform 1 0 4048 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_23
timestamp 1607721120
transform 1 0 3220 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607721120
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0981_
timestamp 1607721120
transform 1 0 4140 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1291_
timestamp 1607721120
transform 1 0 5520 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_74_75
timestamp 1607721120
transform 1 0 8004 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_67
timestamp 1607721120
transform 1 0 7268 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0956_
timestamp 1607721120
transform 1 0 8188 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_74_84
timestamp 1607721120
transform 1 0 8832 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607721120
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1297_
timestamp 1607721120
transform 1 0 9660 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_74_112
timestamp 1607721120
transform 1 0 11408 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1299_
timestamp 1607721120
transform 1 0 12144 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_139
timestamp 1607721120
transform 1 0 13892 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_162
timestamp 1607721120
transform 1 0 16008 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_154
timestamp 1607721120
transform 1 0 15272 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_151
timestamp 1607721120
transform 1 0 14996 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607721120
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0866_
timestamp 1607721120
transform 1 0 15364 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1309_
timestamp 1607721120
transform 1 0 16744 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_201
timestamp 1607721120
transform 1 0 19596 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_189
timestamp 1607721120
transform 1 0 18492 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_227
timestamp 1607721120
transform 1 0 21988 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_215
timestamp 1607721120
transform 1 0 20884 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_213
timestamp 1607721120
transform 1 0 20700 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607721120
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_239
timestamp 1607721120
transform 1 0 23092 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_251
timestamp 1607721120
transform 1 0 24196 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607721120
transform -1 0 24840 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_15
timestamp 1607721120
transform 1 0 2484 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1607721120
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607721120
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1607721120
transform 1 0 4140 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_23
timestamp 1607721120
transform 1 0 3220 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1005_
timestamp 1607721120
transform 1 0 3496 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_75_62
timestamp 1607721120
transform 1 0 6808 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_53
timestamp 1607721120
transform 1 0 5980 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_45
timestamp 1607721120
transform 1 0 5244 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607721120
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0970_
timestamp 1607721120
transform 1 0 5336 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_75_77
timestamp 1607721120
transform 1 0 8188 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0964_
timestamp 1607721120
transform 1 0 7544 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_75_92
timestamp 1607721120
transform 1 0 9568 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0946_
timestamp 1607721120
transform 1 0 8924 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0938_
timestamp 1607721120
transform 1 0 10304 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1607721120
transform 1 0 12236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_109
timestamp 1607721120
transform 1 0 11132 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607721120
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1302_
timestamp 1607721120
transform 1 0 12420 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_75_142
timestamp 1607721120
transform 1 0 14168 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1304_
timestamp 1607721120
transform 1 0 14904 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_75_181
timestamp 1607721120
transform 1 0 17756 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1607721120
transform 1 0 16652 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607721120
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0880_
timestamp 1607721120
transform 1 0 18032 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_203
timestamp 1607721120
transform 1 0 19780 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_191
timestamp 1607721120
transform 1 0 18676 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_227
timestamp 1607721120
transform 1 0 21988 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_215
timestamp 1607721120
transform 1 0 20884 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_245
timestamp 1607721120
transform 1 0 23644 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_243
timestamp 1607721120
transform 1 0 23460 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_239
timestamp 1607721120
transform 1 0 23092 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607721120
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_253
timestamp 1607721120
transform 1 0 24380 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607721120
transform -1 0 24840 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607721120
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607721120
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1607721120
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_38
timestamp 1607721120
transform 1 0 4600 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_32
timestamp 1607721120
transform 1 0 4048 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607721120
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607721120
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0998_
timestamp 1607721120
transform 1 0 4692 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_76_61
timestamp 1607721120
transform 1 0 6716 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_56
timestamp 1607721120
transform 1 0 6256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_48
timestamp 1607721120
transform 1 0 5520 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1607721120
transform 1 0 6348 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_78
timestamp 1607721120
transform 1 0 8280 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0963_
timestamp 1607721120
transform 1 0 7452 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_76_97
timestamp 1607721120
transform 1 0 10028 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_93
timestamp 1607721120
transform 1 0 9660 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_90
timestamp 1607721120
transform 1 0 9384 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607721120
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0934_
timestamp 1607721120
transform 1 0 10120 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_76_122
timestamp 1607721120
transform 1 0 12328 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_105
timestamp 1607721120
transform 1 0 10764 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0920_
timestamp 1607721120
transform 1 0 11500 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_76_142
timestamp 1607721120
transform 1 0 14168 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_130
timestamp 1607721120
transform 1 0 13064 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0908_
timestamp 1607721120
transform 1 0 13340 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_76_154
timestamp 1607721120
transform 1 0 15272 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_150
timestamp 1607721120
transform 1 0 14904 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607721120
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1308_
timestamp 1607721120
transform 1 0 16008 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_76_181
timestamp 1607721120
transform 1 0 17756 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_205
timestamp 1607721120
transform 1 0 19964 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_193
timestamp 1607721120
transform 1 0 18860 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_227
timestamp 1607721120
transform 1 0 21988 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_215
timestamp 1607721120
transform 1 0 20884 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_213
timestamp 1607721120
transform 1 0 20700 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607721120
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_239
timestamp 1607721120
transform 1 0 23092 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_251
timestamp 1607721120
transform 1 0 24196 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607721120
transform -1 0 24840 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_15
timestamp 1607721120
transform 1 0 2484 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1607721120
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1607721120
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0994_
timestamp 1607721120
transform 1 0 2852 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_77_26
timestamp 1607721120
transform 1 0 3496 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1289_
timestamp 1607721120
transform 1 0 4232 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_77_62
timestamp 1607721120
transform 1 0 6808 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_77_53
timestamp 1607721120
transform 1 0 5980 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607721120
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_70
timestamp 1607721120
transform 1 0 7544 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1295_
timestamp 1607721120
transform 1 0 7636 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_77_98
timestamp 1607721120
transform 1 0 10120 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_90
timestamp 1607721120
transform 1 0 9384 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0933_
timestamp 1607721120
transform 1 0 10304 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_77_123
timestamp 1607721120
transform 1 0 12420 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_121
timestamp 1607721120
transform 1 0 12236 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_109
timestamp 1607721120
transform 1 0 11132 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607721120
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0916_
timestamp 1607721120
transform 1 0 12512 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_77_131
timestamp 1607721120
transform 1 0 13156 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0891_
timestamp 1607721120
transform 1 0 13892 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_77_163
timestamp 1607721120
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_77_146
timestamp 1607721120
transform 1 0 14536 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0884_
timestamp 1607721120
transform 1 0 15272 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1607721120
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_175
timestamp 1607721120
transform 1 0 17204 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607721120
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0909_
timestamp 1607721120
transform 1 0 16836 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1607721120
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1607721120
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_220
timestamp 1607721120
transform 1 0 21344 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_245
timestamp 1607721120
transform 1 0 23644 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_232
timestamp 1607721120
transform 1 0 22448 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607721120
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_253
timestamp 1607721120
transform 1 0 24380 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1607721120
transform -1 0 24840 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1607721120
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1607721120
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1607721120
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_78_32
timestamp 1607721120
transform 1 0 4048 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1607721120
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607721120
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0980_
timestamp 1607721120
transform 1 0 4600 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_78_47
timestamp 1607721120
transform 1 0 5428 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1292_
timestamp 1607721120
transform 1 0 6164 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_78_74
timestamp 1607721120
transform 1 0 7912 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_102
timestamp 1607721120
transform 1 0 10488 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_86
timestamp 1607721120
transform 1 0 9016 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607721120
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0944_
timestamp 1607721120
transform 1 0 9660 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_78_119
timestamp 1607721120
transform 1 0 12052 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0925_
timestamp 1607721120
transform 1 0 11224 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_78_136
timestamp 1607721120
transform 1 0 13616 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0914_
timestamp 1607721120
transform 1 0 12788 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_78_162
timestamp 1607721120
transform 1 0 16008 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_154
timestamp 1607721120
transform 1 0 15272 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_152
timestamp 1607721120
transform 1 0 15088 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_148
timestamp 1607721120
transform 1 0 14720 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607721120
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1307_
timestamp 1607721120
transform 1 0 16100 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_78_182
timestamp 1607721120
transform 1 0 17848 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_206
timestamp 1607721120
transform 1 0 20056 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_194
timestamp 1607721120
transform 1 0 18952 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_227
timestamp 1607721120
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_215
timestamp 1607721120
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607721120
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_239
timestamp 1607721120
transform 1 0 23092 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_251
timestamp 1607721120
transform 1 0 24196 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1607721120
transform -1 0 24840 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1607721120
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1607721120
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1607721120
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1607721120
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1607721120
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1607721120
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_40
timestamp 1607721120
transform 1 0 4784 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_32
timestamp 1607721120
transform 1 0 4048 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_27
timestamp 1607721120
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_39
timestamp 1607721120
transform 1 0 4692 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1607721120
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607721120
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1290_
timestamp 1607721120
transform 1 0 4876 0 -1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_80_60
timestamp 1607721120
transform 1 0 6624 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_59
timestamp 1607721120
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_51
timestamp 1607721120
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607721120
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0993_
timestamp 1607721120
transform 1 0 4968 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0976_
timestamp 1607721120
transform 1 0 6808 0 1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_80_76
timestamp 1607721120
transform 1 0 8096 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_72
timestamp 1607721120
transform 1 0 7728 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_77
timestamp 1607721120
transform 1 0 8188 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_69
timestamp 1607721120
transform 1 0 7452 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0955_
timestamp 1607721120
transform 1 0 8280 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0951_
timestamp 1607721120
transform 1 0 8188 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_80_101
timestamp 1607721120
transform 1 0 10396 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_93
timestamp 1607721120
transform 1 0 9660 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_84
timestamp 1607721120
transform 1 0 8832 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_87
timestamp 1607721120
transform 1 0 9108 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607721120
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1300_
timestamp 1607721120
transform 1 0 10672 0 -1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1298_
timestamp 1607721120
transform 1 0 9844 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1607721120
transform 1 0 12420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_114
timestamp 1607721120
transform 1 0 11592 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607721120
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1301_
timestamp 1607721120
transform 1 0 12420 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_80_145
timestamp 1607721120
transform 1 0 14444 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_135
timestamp 1607721120
transform 1 0 13524 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_142
timestamp 1607721120
transform 1 0 14168 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0903_
timestamp 1607721120
transform 1 0 13616 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_80_162
timestamp 1607721120
transform 1 0 16008 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_154
timestamp 1607721120
transform 1 0 15272 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607721120
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1306_
timestamp 1607721120
transform 1 0 16100 0 -1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1303_
timestamp 1607721120
transform 1 0 14904 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_80_182
timestamp 1607721120
transform 1 0 17848 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_181
timestamp 1607721120
transform 1 0 17756 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1607721120
transform 1 0 16652 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607721120
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0886_
timestamp 1607721120
transform 1 0 18032 0 1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_80_206
timestamp 1607721120
transform 1 0 20056 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_194
timestamp 1607721120
transform 1 0 18952 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_203
timestamp 1607721120
transform 1 0 19780 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_191
timestamp 1607721120
transform 1 0 18676 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_227
timestamp 1607721120
transform 1 0 21988 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_215
timestamp 1607721120
transform 1 0 20884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_227
timestamp 1607721120
transform 1 0 21988 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_215
timestamp 1607721120
transform 1 0 20884 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607721120
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_239
timestamp 1607721120
transform 1 0 23092 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_245
timestamp 1607721120
transform 1 0 23644 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_243
timestamp 1607721120
transform 1 0 23460 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_239
timestamp 1607721120
transform 1 0 23092 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607721120
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_251
timestamp 1607721120
transform 1 0 24196 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_253
timestamp 1607721120
transform 1 0 24380 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1607721120
transform -1 0 24840 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1607721120
transform -1 0 24840 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1607721120
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1607721120
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1607721120
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_39
timestamp 1607721120
transform 1 0 4692 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1607721120
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_62
timestamp 1607721120
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_53
timestamp 1607721120
transform 1 0 5980 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_45
timestamp 1607721120
transform 1 0 5244 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607721120
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0986_
timestamp 1607721120
transform 1 0 5336 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_81_74
timestamp 1607721120
transform 1 0 7912 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1296_
timestamp 1607721120
transform 1 0 8648 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_81_101
timestamp 1607721120
transform 1 0 10396 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_121
timestamp 1607721120
transform 1 0 12236 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1607721120
transform 1 0 11500 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607721120
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0915_
timestamp 1607721120
transform 1 0 11132 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0910_
timestamp 1607721120
transform 1 0 12420 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_81_130
timestamp 1607721120
transform 1 0 13064 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1305_
timestamp 1607721120
transform 1 0 13800 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_81_157
timestamp 1607721120
transform 1 0 15548 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0895_
timestamp 1607721120
transform 1 0 16284 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1607721120
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_182
timestamp 1607721120
transform 1 0 17848 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_174
timestamp 1607721120
transform 1 0 17112 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607721120
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_208
timestamp 1607721120
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1607721120
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_220
timestamp 1607721120
transform 1 0 21344 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_245
timestamp 1607721120
transform 1 0 23644 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_232
timestamp 1607721120
transform 1 0 22448 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607721120
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_253
timestamp 1607721120
transform 1 0 24380 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1607721120
transform -1 0 24840 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1607721120
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1607721120
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1607721120
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1607721120
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1607721120
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607721120
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_56
timestamp 1607721120
transform 1 0 6256 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1607721120
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607721120
transform 1 0 6808 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_75
timestamp 1607721120
transform 1 0 8004 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_63
timestamp 1607721120
transform 1 0 6900 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_101
timestamp 1607721120
transform 1 0 10396 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_87
timestamp 1607721120
transform 1 0 9108 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607721120
transform 1 0 9660 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0940_
timestamp 1607721120
transform 1 0 9752 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_82_116
timestamp 1607721120
transform 1 0 11776 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607721120
transform 1 0 12512 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0926_
timestamp 1607721120
transform 1 0 11132 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0921_
timestamp 1607721120
transform 1 0 12604 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1607721120
transform 1 0 13248 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0896_
timestamp 1607721120
transform 1 0 13984 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1607721120
transform 1 0 16284 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_147
timestamp 1607721120
transform 1 0 14628 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607721120
transform 1 0 15364 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0890_
timestamp 1607721120
transform 1 0 15456 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_82_187
timestamp 1607721120
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_185
timestamp 1607721120
transform 1 0 18124 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_177
timestamp 1607721120
transform 1 0 17388 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607721120
transform 1 0 18216 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_199
timestamp 1607721120
transform 1 0 19412 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_218
timestamp 1607721120
transform 1 0 21160 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_211
timestamp 1607721120
transform 1 0 20516 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607721120
transform 1 0 21068 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_249
timestamp 1607721120
transform 1 0 24012 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_242
timestamp 1607721120
transform 1 0 23368 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_230
timestamp 1607721120
transform 1 0 22264 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607721120
transform 1 0 23920 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1607721120
transform -1 0 24840 0 -1 47328
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 2728 800 2848 6 cen
port 0 nsew default tristate
rlabel metal3 s 0 8168 800 8288 6 set_out[0]
port 1 nsew default tristate
rlabel metal3 s 0 13744 800 13864 6 set_out[1]
port 2 nsew default tristate
rlabel metal3 s 0 19320 800 19440 6 set_out[2]
port 3 nsew default tristate
rlabel metal3 s 0 24896 800 25016 6 set_out[3]
port 4 nsew default tristate
rlabel metal3 s 0 30472 800 30592 6 shift_out[0]
port 5 nsew default tristate
rlabel metal3 s 0 36048 800 36168 6 shift_out[1]
port 6 nsew default tristate
rlabel metal3 s 0 41624 800 41744 6 shift_out[2]
port 7 nsew default tristate
rlabel metal3 s 0 47200 800 47320 6 shift_out[3]
port 8 nsew default tristate
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 9 nsew default input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 10 nsew default input
rlabel metal2 s 386 49200 442 50000 6 wbs_ack_o
port 11 nsew default tristate
rlabel metal2 s 14646 0 14702 800 6 wbs_addr_i[0]
port 12 nsew default input
rlabel metal2 s 18234 0 18290 800 6 wbs_addr_i[10]
port 13 nsew default input
rlabel metal2 s 18602 0 18658 800 6 wbs_addr_i[11]
port 14 nsew default input
rlabel metal2 s 18970 0 19026 800 6 wbs_addr_i[12]
port 15 nsew default input
rlabel metal2 s 19338 0 19394 800 6 wbs_addr_i[13]
port 16 nsew default input
rlabel metal2 s 19706 0 19762 800 6 wbs_addr_i[14]
port 17 nsew default input
rlabel metal2 s 20074 0 20130 800 6 wbs_addr_i[15]
port 18 nsew default input
rlabel metal2 s 20350 0 20406 800 6 wbs_addr_i[16]
port 19 nsew default input
rlabel metal2 s 20718 0 20774 800 6 wbs_addr_i[17]
port 20 nsew default input
rlabel metal2 s 21086 0 21142 800 6 wbs_addr_i[18]
port 21 nsew default input
rlabel metal2 s 21454 0 21510 800 6 wbs_addr_i[19]
port 22 nsew default input
rlabel metal2 s 15014 0 15070 800 6 wbs_addr_i[1]
port 23 nsew default input
rlabel metal2 s 21822 0 21878 800 6 wbs_addr_i[20]
port 24 nsew default input
rlabel metal2 s 22190 0 22246 800 6 wbs_addr_i[21]
port 25 nsew default input
rlabel metal2 s 22558 0 22614 800 6 wbs_addr_i[22]
port 26 nsew default input
rlabel metal2 s 22926 0 22982 800 6 wbs_addr_i[23]
port 27 nsew default input
rlabel metal2 s 23202 0 23258 800 6 wbs_addr_i[24]
port 28 nsew default input
rlabel metal2 s 23570 0 23626 800 6 wbs_addr_i[25]
port 29 nsew default input
rlabel metal2 s 23938 0 23994 800 6 wbs_addr_i[26]
port 30 nsew default input
rlabel metal2 s 24306 0 24362 800 6 wbs_addr_i[27]
port 31 nsew default input
rlabel metal2 s 24674 0 24730 800 6 wbs_addr_i[28]
port 32 nsew default input
rlabel metal2 s 25042 0 25098 800 6 wbs_addr_i[29]
port 33 nsew default input
rlabel metal2 s 15382 0 15438 800 6 wbs_addr_i[2]
port 34 nsew default input
rlabel metal2 s 25410 0 25466 800 6 wbs_addr_i[30]
port 35 nsew default input
rlabel metal2 s 25778 0 25834 800 6 wbs_addr_i[31]
port 36 nsew default input
rlabel metal2 s 15750 0 15806 800 6 wbs_addr_i[3]
port 37 nsew default input
rlabel metal2 s 16118 0 16174 800 6 wbs_addr_i[4]
port 38 nsew default input
rlabel metal2 s 16486 0 16542 800 6 wbs_addr_i[5]
port 39 nsew default input
rlabel metal2 s 16854 0 16910 800 6 wbs_addr_i[6]
port 40 nsew default input
rlabel metal2 s 17222 0 17278 800 6 wbs_addr_i[7]
port 41 nsew default input
rlabel metal2 s 17498 0 17554 800 6 wbs_addr_i[8]
port 42 nsew default input
rlabel metal2 s 17866 0 17922 800 6 wbs_addr_i[9]
port 43 nsew default input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 44 nsew default input
rlabel metal2 s 3238 0 3294 800 6 wbs_data_i[0]
port 45 nsew default input
rlabel metal2 s 6826 0 6882 800 6 wbs_data_i[10]
port 46 nsew default input
rlabel metal2 s 7194 0 7250 800 6 wbs_data_i[11]
port 47 nsew default input
rlabel metal2 s 7562 0 7618 800 6 wbs_data_i[12]
port 48 nsew default input
rlabel metal2 s 7930 0 7986 800 6 wbs_data_i[13]
port 49 nsew default input
rlabel metal2 s 8298 0 8354 800 6 wbs_data_i[14]
port 50 nsew default input
rlabel metal2 s 8666 0 8722 800 6 wbs_data_i[15]
port 51 nsew default input
rlabel metal2 s 8942 0 8998 800 6 wbs_data_i[16]
port 52 nsew default input
rlabel metal2 s 9310 0 9366 800 6 wbs_data_i[17]
port 53 nsew default input
rlabel metal2 s 9678 0 9734 800 6 wbs_data_i[18]
port 54 nsew default input
rlabel metal2 s 10046 0 10102 800 6 wbs_data_i[19]
port 55 nsew default input
rlabel metal2 s 3606 0 3662 800 6 wbs_data_i[1]
port 56 nsew default input
rlabel metal2 s 10414 0 10470 800 6 wbs_data_i[20]
port 57 nsew default input
rlabel metal2 s 10782 0 10838 800 6 wbs_data_i[21]
port 58 nsew default input
rlabel metal2 s 11150 0 11206 800 6 wbs_data_i[22]
port 59 nsew default input
rlabel metal2 s 11518 0 11574 800 6 wbs_data_i[23]
port 60 nsew default input
rlabel metal2 s 11794 0 11850 800 6 wbs_data_i[24]
port 61 nsew default input
rlabel metal2 s 12162 0 12218 800 6 wbs_data_i[25]
port 62 nsew default input
rlabel metal2 s 12530 0 12586 800 6 wbs_data_i[26]
port 63 nsew default input
rlabel metal2 s 12898 0 12954 800 6 wbs_data_i[27]
port 64 nsew default input
rlabel metal2 s 13266 0 13322 800 6 wbs_data_i[28]
port 65 nsew default input
rlabel metal2 s 13634 0 13690 800 6 wbs_data_i[29]
port 66 nsew default input
rlabel metal2 s 3974 0 4030 800 6 wbs_data_i[2]
port 67 nsew default input
rlabel metal2 s 14002 0 14058 800 6 wbs_data_i[30]
port 68 nsew default input
rlabel metal2 s 14370 0 14426 800 6 wbs_data_i[31]
port 69 nsew default input
rlabel metal2 s 4342 0 4398 800 6 wbs_data_i[3]
port 70 nsew default input
rlabel metal2 s 4710 0 4766 800 6 wbs_data_i[4]
port 71 nsew default input
rlabel metal2 s 5078 0 5134 800 6 wbs_data_i[5]
port 72 nsew default input
rlabel metal2 s 5446 0 5502 800 6 wbs_data_i[6]
port 73 nsew default input
rlabel metal2 s 5814 0 5870 800 6 wbs_data_i[7]
port 74 nsew default input
rlabel metal2 s 6090 0 6146 800 6 wbs_data_i[8]
port 75 nsew default input
rlabel metal2 s 6458 0 6514 800 6 wbs_data_i[9]
port 76 nsew default input
rlabel metal2 s 1122 49200 1178 50000 6 wbs_data_o[0]
port 77 nsew default tristate
rlabel metal2 s 9034 49200 9090 50000 6 wbs_data_o[10]
port 78 nsew default tristate
rlabel metal2 s 9770 49200 9826 50000 6 wbs_data_o[11]
port 79 nsew default tristate
rlabel metal2 s 10598 49200 10654 50000 6 wbs_data_o[12]
port 80 nsew default tristate
rlabel metal2 s 11426 49200 11482 50000 6 wbs_data_o[13]
port 81 nsew default tristate
rlabel metal2 s 12162 49200 12218 50000 6 wbs_data_o[14]
port 82 nsew default tristate
rlabel metal2 s 12990 49200 13046 50000 6 wbs_data_o[15]
port 83 nsew default tristate
rlabel metal2 s 13726 49200 13782 50000 6 wbs_data_o[16]
port 84 nsew default tristate
rlabel metal2 s 14554 49200 14610 50000 6 wbs_data_o[17]
port 85 nsew default tristate
rlabel metal2 s 15290 49200 15346 50000 6 wbs_data_o[18]
port 86 nsew default tristate
rlabel metal2 s 16118 49200 16174 50000 6 wbs_data_o[19]
port 87 nsew default tristate
rlabel metal2 s 1950 49200 2006 50000 6 wbs_data_o[1]
port 88 nsew default tristate
rlabel metal2 s 16946 49200 17002 50000 6 wbs_data_o[20]
port 89 nsew default tristate
rlabel metal2 s 17682 49200 17738 50000 6 wbs_data_o[21]
port 90 nsew default tristate
rlabel metal2 s 18510 49200 18566 50000 6 wbs_data_o[22]
port 91 nsew default tristate
rlabel metal2 s 19246 49200 19302 50000 6 wbs_data_o[23]
port 92 nsew default tristate
rlabel metal2 s 20074 49200 20130 50000 6 wbs_data_o[24]
port 93 nsew default tristate
rlabel metal2 s 20810 49200 20866 50000 6 wbs_data_o[25]
port 94 nsew default tristate
rlabel metal2 s 21638 49200 21694 50000 6 wbs_data_o[26]
port 95 nsew default tristate
rlabel metal2 s 22466 49200 22522 50000 6 wbs_data_o[27]
port 96 nsew default tristate
rlabel metal2 s 23202 49200 23258 50000 6 wbs_data_o[28]
port 97 nsew default tristate
rlabel metal2 s 24030 49200 24086 50000 6 wbs_data_o[29]
port 98 nsew default tristate
rlabel metal2 s 2686 49200 2742 50000 6 wbs_data_o[2]
port 99 nsew default tristate
rlabel metal2 s 24766 49200 24822 50000 6 wbs_data_o[30]
port 100 nsew default tristate
rlabel metal2 s 25594 49200 25650 50000 6 wbs_data_o[31]
port 101 nsew default tristate
rlabel metal2 s 3514 49200 3570 50000 6 wbs_data_o[3]
port 102 nsew default tristate
rlabel metal2 s 4250 49200 4306 50000 6 wbs_data_o[4]
port 103 nsew default tristate
rlabel metal2 s 5078 49200 5134 50000 6 wbs_data_o[5]
port 104 nsew default tristate
rlabel metal2 s 5906 49200 5962 50000 6 wbs_data_o[6]
port 105 nsew default tristate
rlabel metal2 s 6642 49200 6698 50000 6 wbs_data_o[7]
port 106 nsew default tristate
rlabel metal2 s 7470 49200 7526 50000 6 wbs_data_o[8]
port 107 nsew default tristate
rlabel metal2 s 8206 49200 8262 50000 6 wbs_data_o[9]
port 108 nsew default tristate
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 109 nsew default input
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[1]
port 110 nsew default input
rlabel metal2 s 2594 0 2650 800 6 wbs_sel_i[2]
port 111 nsew default input
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[3]
port 112 nsew default input
rlabel metal2 s 754 0 810 800 6 wbs_stb_i
port 113 nsew default input
rlabel metal2 s 1490 0 1546 800 6 wbs_we_i
port 114 nsew default input
rlabel metal5 s 1104 9576 24840 9896 6 VPWR
port 115 nsew default input
rlabel metal5 s 1104 17184 24840 17504 6 VGND
port 116 nsew default input
<< properties >>
string FIXED_BBOX 0 0 25838 50000
<< end >>
