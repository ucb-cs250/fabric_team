VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO baked_disjoint_switch_box
  CLASS BLOCK ;
  FOREIGN baked_disjoint_switch_box ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END cen
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 694.230 696.000 694.510 700.000 ;
    END
  END cset
  PIN cset_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END cset_out
  PIN east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 1.400 700.000 2.000 ;
    END
  END east[0]
  PIN east[100]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 359.760 700.000 360.360 ;
    END
  END east[100]
  PIN east[101]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 363.160 700.000 363.760 ;
    END
  END east[101]
  PIN east[102]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END east[102]
  PIN east[103]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 370.640 700.000 371.240 ;
    END
  END east[103]
  PIN east[104]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 374.040 700.000 374.640 ;
    END
  END east[104]
  PIN east[105]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 378.120 700.000 378.720 ;
    END
  END east[105]
  PIN east[106]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 381.520 700.000 382.120 ;
    END
  END east[106]
  PIN east[107]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 384.920 700.000 385.520 ;
    END
  END east[107]
  PIN east[108]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 388.320 700.000 388.920 ;
    END
  END east[108]
  PIN east[109]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 392.400 700.000 393.000 ;
    END
  END east[109]
  PIN east[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 36.760 700.000 37.360 ;
    END
  END east[10]
  PIN east[110]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 395.800 700.000 396.400 ;
    END
  END east[110]
  PIN east[111]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 399.200 700.000 399.800 ;
    END
  END east[111]
  PIN east[112]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 403.280 700.000 403.880 ;
    END
  END east[112]
  PIN east[113]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 406.680 700.000 407.280 ;
    END
  END east[113]
  PIN east[114]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 410.080 700.000 410.680 ;
    END
  END east[114]
  PIN east[115]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 413.480 700.000 414.080 ;
    END
  END east[115]
  PIN east[116]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 417.560 700.000 418.160 ;
    END
  END east[116]
  PIN east[117]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 420.960 700.000 421.560 ;
    END
  END east[117]
  PIN east[118]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 424.360 700.000 424.960 ;
    END
  END east[118]
  PIN east[119]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 427.760 700.000 428.360 ;
    END
  END east[119]
  PIN east[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 40.840 700.000 41.440 ;
    END
  END east[11]
  PIN east[120]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 431.840 700.000 432.440 ;
    END
  END east[120]
  PIN east[121]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 435.240 700.000 435.840 ;
    END
  END east[121]
  PIN east[122]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 438.640 700.000 439.240 ;
    END
  END east[122]
  PIN east[123]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 442.720 700.000 443.320 ;
    END
  END east[123]
  PIN east[124]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 446.120 700.000 446.720 ;
    END
  END east[124]
  PIN east[125]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 449.520 700.000 450.120 ;
    END
  END east[125]
  PIN east[126]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 452.920 700.000 453.520 ;
    END
  END east[126]
  PIN east[127]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 457.000 700.000 457.600 ;
    END
  END east[127]
  PIN east[128]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 460.400 700.000 461.000 ;
    END
  END east[128]
  PIN east[129]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 463.800 700.000 464.400 ;
    END
  END east[129]
  PIN east[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 44.240 700.000 44.840 ;
    END
  END east[12]
  PIN east[130]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 467.880 700.000 468.480 ;
    END
  END east[130]
  PIN east[131]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 471.280 700.000 471.880 ;
    END
  END east[131]
  PIN east[132]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 474.680 700.000 475.280 ;
    END
  END east[132]
  PIN east[133]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 478.080 700.000 478.680 ;
    END
  END east[133]
  PIN east[134]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 482.160 700.000 482.760 ;
    END
  END east[134]
  PIN east[135]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 485.560 700.000 486.160 ;
    END
  END east[135]
  PIN east[136]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 488.960 700.000 489.560 ;
    END
  END east[136]
  PIN east[137]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 492.360 700.000 492.960 ;
    END
  END east[137]
  PIN east[138]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 496.440 700.000 497.040 ;
    END
  END east[138]
  PIN east[139]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 499.840 700.000 500.440 ;
    END
  END east[139]
  PIN east[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 47.640 700.000 48.240 ;
    END
  END east[13]
  PIN east[140]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 503.240 700.000 503.840 ;
    END
  END east[140]
  PIN east[141]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 507.320 700.000 507.920 ;
    END
  END east[141]
  PIN east[142]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 510.720 700.000 511.320 ;
    END
  END east[142]
  PIN east[143]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 514.120 700.000 514.720 ;
    END
  END east[143]
  PIN east[144]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 517.520 700.000 518.120 ;
    END
  END east[144]
  PIN east[145]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 521.600 700.000 522.200 ;
    END
  END east[145]
  PIN east[146]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 525.000 700.000 525.600 ;
    END
  END east[146]
  PIN east[147]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 528.400 700.000 529.000 ;
    END
  END east[147]
  PIN east[148]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 531.800 700.000 532.400 ;
    END
  END east[148]
  PIN east[149]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 535.880 700.000 536.480 ;
    END
  END east[149]
  PIN east[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 51.040 700.000 51.640 ;
    END
  END east[14]
  PIN east[150]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 539.280 700.000 539.880 ;
    END
  END east[150]
  PIN east[151]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 542.680 700.000 543.280 ;
    END
  END east[151]
  PIN east[152]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 546.760 700.000 547.360 ;
    END
  END east[152]
  PIN east[153]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 550.160 700.000 550.760 ;
    END
  END east[153]
  PIN east[154]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 553.560 700.000 554.160 ;
    END
  END east[154]
  PIN east[155]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 556.960 700.000 557.560 ;
    END
  END east[155]
  PIN east[156]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 561.040 700.000 561.640 ;
    END
  END east[156]
  PIN east[157]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 564.440 700.000 565.040 ;
    END
  END east[157]
  PIN east[158]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 567.840 700.000 568.440 ;
    END
  END east[158]
  PIN east[159]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 571.920 700.000 572.520 ;
    END
  END east[159]
  PIN east[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 55.120 700.000 55.720 ;
    END
  END east[15]
  PIN east[160]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 575.320 700.000 575.920 ;
    END
  END east[160]
  PIN east[161]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 578.720 700.000 579.320 ;
    END
  END east[161]
  PIN east[162]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 582.120 700.000 582.720 ;
    END
  END east[162]
  PIN east[163]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 586.200 700.000 586.800 ;
    END
  END east[163]
  PIN east[164]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 589.600 700.000 590.200 ;
    END
  END east[164]
  PIN east[165]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 593.000 700.000 593.600 ;
    END
  END east[165]
  PIN east[166]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 596.400 700.000 597.000 ;
    END
  END east[166]
  PIN east[167]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 600.480 700.000 601.080 ;
    END
  END east[167]
  PIN east[168]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 603.880 700.000 604.480 ;
    END
  END east[168]
  PIN east[169]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 607.280 700.000 607.880 ;
    END
  END east[169]
  PIN east[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 58.520 700.000 59.120 ;
    END
  END east[16]
  PIN east[170]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 611.360 700.000 611.960 ;
    END
  END east[170]
  PIN east[171]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 614.760 700.000 615.360 ;
    END
  END east[171]
  PIN east[172]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 618.160 700.000 618.760 ;
    END
  END east[172]
  PIN east[173]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 621.560 700.000 622.160 ;
    END
  END east[173]
  PIN east[174]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 625.640 700.000 626.240 ;
    END
  END east[174]
  PIN east[175]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 629.040 700.000 629.640 ;
    END
  END east[175]
  PIN east[176]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 632.440 700.000 633.040 ;
    END
  END east[176]
  PIN east[177]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 636.520 700.000 637.120 ;
    END
  END east[177]
  PIN east[178]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 639.920 700.000 640.520 ;
    END
  END east[178]
  PIN east[179]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 643.320 700.000 643.920 ;
    END
  END east[179]
  PIN east[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 61.920 700.000 62.520 ;
    END
  END east[17]
  PIN east[180]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 646.720 700.000 647.320 ;
    END
  END east[180]
  PIN east[181]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 650.800 700.000 651.400 ;
    END
  END east[181]
  PIN east[182]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 654.200 700.000 654.800 ;
    END
  END east[182]
  PIN east[183]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 657.600 700.000 658.200 ;
    END
  END east[183]
  PIN east[184]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 661.000 700.000 661.600 ;
    END
  END east[184]
  PIN east[185]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 665.080 700.000 665.680 ;
    END
  END east[185]
  PIN east[186]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 668.480 700.000 669.080 ;
    END
  END east[186]
  PIN east[187]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 671.880 700.000 672.480 ;
    END
  END east[187]
  PIN east[188]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 675.960 700.000 676.560 ;
    END
  END east[188]
  PIN east[189]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 679.360 700.000 679.960 ;
    END
  END east[189]
  PIN east[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 65.320 700.000 65.920 ;
    END
  END east[18]
  PIN east[190]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 682.760 700.000 683.360 ;
    END
  END east[190]
  PIN east[191]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 686.160 700.000 686.760 ;
    END
  END east[191]
  PIN east[192]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 690.240 700.000 690.840 ;
    END
  END east[192]
  PIN east[193]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 693.640 700.000 694.240 ;
    END
  END east[193]
  PIN east[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 69.400 700.000 70.000 ;
    END
  END east[19]
  PIN east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 4.800 700.000 5.400 ;
    END
  END east[1]
  PIN east[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 72.800 700.000 73.400 ;
    END
  END east[20]
  PIN east[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 76.200 700.000 76.800 ;
    END
  END east[21]
  PIN east[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 80.280 700.000 80.880 ;
    END
  END east[22]
  PIN east[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 83.680 700.000 84.280 ;
    END
  END east[23]
  PIN east[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 87.080 700.000 87.680 ;
    END
  END east[24]
  PIN east[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 90.480 700.000 91.080 ;
    END
  END east[25]
  PIN east[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 94.560 700.000 95.160 ;
    END
  END east[26]
  PIN east[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 97.960 700.000 98.560 ;
    END
  END east[27]
  PIN east[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 101.360 700.000 101.960 ;
    END
  END east[28]
  PIN east[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 105.440 700.000 106.040 ;
    END
  END east[29]
  PIN east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 8.200 700.000 8.800 ;
    END
  END east[2]
  PIN east[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 108.840 700.000 109.440 ;
    END
  END east[30]
  PIN east[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 112.240 700.000 112.840 ;
    END
  END east[31]
  PIN east[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 115.640 700.000 116.240 ;
    END
  END east[32]
  PIN east[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 119.720 700.000 120.320 ;
    END
  END east[33]
  PIN east[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 123.120 700.000 123.720 ;
    END
  END east[34]
  PIN east[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 126.520 700.000 127.120 ;
    END
  END east[35]
  PIN east[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 129.920 700.000 130.520 ;
    END
  END east[36]
  PIN east[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 134.000 700.000 134.600 ;
    END
  END east[37]
  PIN east[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 137.400 700.000 138.000 ;
    END
  END east[38]
  PIN east[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 140.800 700.000 141.400 ;
    END
  END east[39]
  PIN east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 11.600 700.000 12.200 ;
    END
  END east[3]
  PIN east[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 144.880 700.000 145.480 ;
    END
  END east[40]
  PIN east[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 148.280 700.000 148.880 ;
    END
  END east[41]
  PIN east[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 151.680 700.000 152.280 ;
    END
  END east[42]
  PIN east[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 155.080 700.000 155.680 ;
    END
  END east[43]
  PIN east[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 159.160 700.000 159.760 ;
    END
  END east[44]
  PIN east[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 162.560 700.000 163.160 ;
    END
  END east[45]
  PIN east[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 165.960 700.000 166.560 ;
    END
  END east[46]
  PIN east[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 170.040 700.000 170.640 ;
    END
  END east[47]
  PIN east[48]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 173.440 700.000 174.040 ;
    END
  END east[48]
  PIN east[49]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 176.840 700.000 177.440 ;
    END
  END east[49]
  PIN east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 15.680 700.000 16.280 ;
    END
  END east[4]
  PIN east[50]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 180.240 700.000 180.840 ;
    END
  END east[50]
  PIN east[51]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 184.320 700.000 184.920 ;
    END
  END east[51]
  PIN east[52]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.720 700.000 188.320 ;
    END
  END east[52]
  PIN east[53]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 191.120 700.000 191.720 ;
    END
  END east[53]
  PIN east[54]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 194.520 700.000 195.120 ;
    END
  END east[54]
  PIN east[55]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 198.600 700.000 199.200 ;
    END
  END east[55]
  PIN east[56]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 202.000 700.000 202.600 ;
    END
  END east[56]
  PIN east[57]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 205.400 700.000 206.000 ;
    END
  END east[57]
  PIN east[58]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 209.480 700.000 210.080 ;
    END
  END east[58]
  PIN east[59]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 212.880 700.000 213.480 ;
    END
  END east[59]
  PIN east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 19.080 700.000 19.680 ;
    END
  END east[5]
  PIN east[60]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 216.280 700.000 216.880 ;
    END
  END east[60]
  PIN east[61]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 219.680 700.000 220.280 ;
    END
  END east[61]
  PIN east[62]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 223.760 700.000 224.360 ;
    END
  END east[62]
  PIN east[63]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 227.160 700.000 227.760 ;
    END
  END east[63]
  PIN east[64]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 230.560 700.000 231.160 ;
    END
  END east[64]
  PIN east[65]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 234.640 700.000 235.240 ;
    END
  END east[65]
  PIN east[66]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.040 700.000 238.640 ;
    END
  END east[66]
  PIN east[67]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 241.440 700.000 242.040 ;
    END
  END east[67]
  PIN east[68]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.840 700.000 245.440 ;
    END
  END east[68]
  PIN east[69]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 248.920 700.000 249.520 ;
    END
  END east[69]
  PIN east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 22.480 700.000 23.080 ;
    END
  END east[6]
  PIN east[70]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 252.320 700.000 252.920 ;
    END
  END east[70]
  PIN east[71]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 255.720 700.000 256.320 ;
    END
  END east[71]
  PIN east[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 259.120 700.000 259.720 ;
    END
  END east[72]
  PIN east[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 263.200 700.000 263.800 ;
    END
  END east[73]
  PIN east[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 266.600 700.000 267.200 ;
    END
  END east[74]
  PIN east[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 270.000 700.000 270.600 ;
    END
  END east[75]
  PIN east[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 274.080 700.000 274.680 ;
    END
  END east[76]
  PIN east[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 277.480 700.000 278.080 ;
    END
  END east[77]
  PIN east[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 280.880 700.000 281.480 ;
    END
  END east[78]
  PIN east[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 284.280 700.000 284.880 ;
    END
  END east[79]
  PIN east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 25.880 700.000 26.480 ;
    END
  END east[7]
  PIN east[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 288.360 700.000 288.960 ;
    END
  END east[80]
  PIN east[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 291.760 700.000 292.360 ;
    END
  END east[81]
  PIN east[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.160 700.000 295.760 ;
    END
  END east[82]
  PIN east[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 298.560 700.000 299.160 ;
    END
  END east[83]
  PIN east[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 302.640 700.000 303.240 ;
    END
  END east[84]
  PIN east[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 306.040 700.000 306.640 ;
    END
  END east[85]
  PIN east[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 309.440 700.000 310.040 ;
    END
  END east[86]
  PIN east[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 313.520 700.000 314.120 ;
    END
  END east[87]
  PIN east[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.920 700.000 317.520 ;
    END
  END east[88]
  PIN east[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 320.320 700.000 320.920 ;
    END
  END east[89]
  PIN east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 29.960 700.000 30.560 ;
    END
  END east[8]
  PIN east[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 323.720 700.000 324.320 ;
    END
  END east[90]
  PIN east[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 327.800 700.000 328.400 ;
    END
  END east[91]
  PIN east[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 331.200 700.000 331.800 ;
    END
  END east[92]
  PIN east[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 334.600 700.000 335.200 ;
    END
  END east[93]
  PIN east[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 338.680 700.000 339.280 ;
    END
  END east[94]
  PIN east[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 342.080 700.000 342.680 ;
    END
  END east[95]
  PIN east[96]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 345.480 700.000 346.080 ;
    END
  END east[96]
  PIN east[97]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 348.880 700.000 349.480 ;
    END
  END east[97]
  PIN east[98]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 352.960 700.000 353.560 ;
    END
  END east[98]
  PIN east[99]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 356.360 700.000 356.960 ;
    END
  END east[99]
  PIN east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 33.360 700.000 33.960 ;
    END
  END east[9]
  PIN north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 696.000 1.750 700.000 ;
    END
  END north[0]
  PIN north[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 356.590 696.000 356.870 700.000 ;
    END
  END north[100]
  PIN north[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 360.270 696.000 360.550 700.000 ;
    END
  END north[101]
  PIN north[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 363.950 696.000 364.230 700.000 ;
    END
  END north[102]
  PIN north[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 367.170 696.000 367.450 700.000 ;
    END
  END north[103]
  PIN north[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 370.850 696.000 371.130 700.000 ;
    END
  END north[104]
  PIN north[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 696.000 374.810 700.000 ;
    END
  END north[105]
  PIN north[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 377.750 696.000 378.030 700.000 ;
    END
  END north[106]
  PIN north[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 381.430 696.000 381.710 700.000 ;
    END
  END north[107]
  PIN north[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 385.110 696.000 385.390 700.000 ;
    END
  END north[108]
  PIN north[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 388.790 696.000 389.070 700.000 ;
    END
  END north[109]
  PIN north[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 696.000 37.170 700.000 ;
    END
  END north[10]
  PIN north[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 392.010 696.000 392.290 700.000 ;
    END
  END north[110]
  PIN north[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 395.690 696.000 395.970 700.000 ;
    END
  END north[111]
  PIN north[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 399.370 696.000 399.650 700.000 ;
    END
  END north[112]
  PIN north[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 696.000 403.330 700.000 ;
    END
  END north[113]
  PIN north[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 406.270 696.000 406.550 700.000 ;
    END
  END north[114]
  PIN north[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 409.950 696.000 410.230 700.000 ;
    END
  END north[115]
  PIN north[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 413.630 696.000 413.910 700.000 ;
    END
  END north[116]
  PIN north[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 696.000 417.130 700.000 ;
    END
  END north[117]
  PIN north[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 420.530 696.000 420.810 700.000 ;
    END
  END north[118]
  PIN north[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 424.210 696.000 424.490 700.000 ;
    END
  END north[119]
  PIN north[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 696.000 40.390 700.000 ;
    END
  END north[11]
  PIN north[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 427.890 696.000 428.170 700.000 ;
    END
  END north[120]
  PIN north[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 431.110 696.000 431.390 700.000 ;
    END
  END north[121]
  PIN north[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 434.790 696.000 435.070 700.000 ;
    END
  END north[122]
  PIN north[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 438.470 696.000 438.750 700.000 ;
    END
  END north[123]
  PIN north[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 442.150 696.000 442.430 700.000 ;
    END
  END north[124]
  PIN north[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 445.370 696.000 445.650 700.000 ;
    END
  END north[125]
  PIN north[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 449.050 696.000 449.330 700.000 ;
    END
  END north[126]
  PIN north[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 452.730 696.000 453.010 700.000 ;
    END
  END north[127]
  PIN north[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 455.950 696.000 456.230 700.000 ;
    END
  END north[128]
  PIN north[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 459.630 696.000 459.910 700.000 ;
    END
  END north[129]
  PIN north[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 696.000 44.070 700.000 ;
    END
  END north[12]
  PIN north[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 696.000 463.590 700.000 ;
    END
  END north[130]
  PIN north[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 466.990 696.000 467.270 700.000 ;
    END
  END north[131]
  PIN north[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 470.210 696.000 470.490 700.000 ;
    END
  END north[132]
  PIN north[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 473.890 696.000 474.170 700.000 ;
    END
  END north[133]
  PIN north[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 477.570 696.000 477.850 700.000 ;
    END
  END north[134]
  PIN north[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 480.790 696.000 481.070 700.000 ;
    END
  END north[135]
  PIN north[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 484.470 696.000 484.750 700.000 ;
    END
  END north[136]
  PIN north[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 488.150 696.000 488.430 700.000 ;
    END
  END north[137]
  PIN north[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 491.830 696.000 492.110 700.000 ;
    END
  END north[138]
  PIN north[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 495.050 696.000 495.330 700.000 ;
    END
  END north[139]
  PIN north[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 696.000 47.750 700.000 ;
    END
  END north[13]
  PIN north[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 498.730 696.000 499.010 700.000 ;
    END
  END north[140]
  PIN north[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 502.410 696.000 502.690 700.000 ;
    END
  END north[141]
  PIN north[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 506.090 696.000 506.370 700.000 ;
    END
  END north[142]
  PIN north[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 509.310 696.000 509.590 700.000 ;
    END
  END north[143]
  PIN north[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 512.990 696.000 513.270 700.000 ;
    END
  END north[144]
  PIN north[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 516.670 696.000 516.950 700.000 ;
    END
  END north[145]
  PIN north[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 519.890 696.000 520.170 700.000 ;
    END
  END north[146]
  PIN north[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 523.570 696.000 523.850 700.000 ;
    END
  END north[147]
  PIN north[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 527.250 696.000 527.530 700.000 ;
    END
  END north[148]
  PIN north[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 530.930 696.000 531.210 700.000 ;
    END
  END north[149]
  PIN north[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 696.000 51.430 700.000 ;
    END
  END north[14]
  PIN north[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 534.150 696.000 534.430 700.000 ;
    END
  END north[150]
  PIN north[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 537.830 696.000 538.110 700.000 ;
    END
  END north[151]
  PIN north[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 541.510 696.000 541.790 700.000 ;
    END
  END north[152]
  PIN north[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 545.190 696.000 545.470 700.000 ;
    END
  END north[153]
  PIN north[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 548.410 696.000 548.690 700.000 ;
    END
  END north[154]
  PIN north[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 552.090 696.000 552.370 700.000 ;
    END
  END north[155]
  PIN north[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 555.770 696.000 556.050 700.000 ;
    END
  END north[156]
  PIN north[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 558.990 696.000 559.270 700.000 ;
    END
  END north[157]
  PIN north[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 562.670 696.000 562.950 700.000 ;
    END
  END north[158]
  PIN north[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 566.350 696.000 566.630 700.000 ;
    END
  END north[159]
  PIN north[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 696.000 54.650 700.000 ;
    END
  END north[15]
  PIN north[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 570.030 696.000 570.310 700.000 ;
    END
  END north[160]
  PIN north[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 573.250 696.000 573.530 700.000 ;
    END
  END north[161]
  PIN north[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 576.930 696.000 577.210 700.000 ;
    END
  END north[162]
  PIN north[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 580.610 696.000 580.890 700.000 ;
    END
  END north[163]
  PIN north[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 584.290 696.000 584.570 700.000 ;
    END
  END north[164]
  PIN north[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 587.510 696.000 587.790 700.000 ;
    END
  END north[165]
  PIN north[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 591.190 696.000 591.470 700.000 ;
    END
  END north[166]
  PIN north[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 594.870 696.000 595.150 700.000 ;
    END
  END north[167]
  PIN north[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 696.000 598.370 700.000 ;
    END
  END north[168]
  PIN north[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 601.770 696.000 602.050 700.000 ;
    END
  END north[169]
  PIN north[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 696.000 58.330 700.000 ;
    END
  END north[16]
  PIN north[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.450 696.000 605.730 700.000 ;
    END
  END north[170]
  PIN north[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 609.130 696.000 609.410 700.000 ;
    END
  END north[171]
  PIN north[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 612.350 696.000 612.630 700.000 ;
    END
  END north[172]
  PIN north[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 616.030 696.000 616.310 700.000 ;
    END
  END north[173]
  PIN north[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 619.710 696.000 619.990 700.000 ;
    END
  END north[174]
  PIN north[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 623.390 696.000 623.670 700.000 ;
    END
  END north[175]
  PIN north[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 626.610 696.000 626.890 700.000 ;
    END
  END north[176]
  PIN north[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 630.290 696.000 630.570 700.000 ;
    END
  END north[177]
  PIN north[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 633.970 696.000 634.250 700.000 ;
    END
  END north[178]
  PIN north[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 637.190 696.000 637.470 700.000 ;
    END
  END north[179]
  PIN north[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 696.000 62.010 700.000 ;
    END
  END north[17]
  PIN north[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 640.870 696.000 641.150 700.000 ;
    END
  END north[180]
  PIN north[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 644.550 696.000 644.830 700.000 ;
    END
  END north[181]
  PIN north[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 648.230 696.000 648.510 700.000 ;
    END
  END north[182]
  PIN north[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 651.450 696.000 651.730 700.000 ;
    END
  END north[183]
  PIN north[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 655.130 696.000 655.410 700.000 ;
    END
  END north[184]
  PIN north[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 658.810 696.000 659.090 700.000 ;
    END
  END north[185]
  PIN north[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 696.000 662.770 700.000 ;
    END
  END north[186]
  PIN north[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 665.710 696.000 665.990 700.000 ;
    END
  END north[187]
  PIN north[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 669.390 696.000 669.670 700.000 ;
    END
  END north[188]
  PIN north[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 673.070 696.000 673.350 700.000 ;
    END
  END north[189]
  PIN north[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 696.000 65.690 700.000 ;
    END
  END north[18]
  PIN north[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 676.290 696.000 676.570 700.000 ;
    END
  END north[190]
  PIN north[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 679.970 696.000 680.250 700.000 ;
    END
  END north[191]
  PIN north[192]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 683.650 696.000 683.930 700.000 ;
    END
  END north[192]
  PIN north[193]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 687.330 696.000 687.610 700.000 ;
    END
  END north[193]
  PIN north[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 696.000 68.910 700.000 ;
    END
  END north[19]
  PIN north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 696.000 4.970 700.000 ;
    END
  END north[1]
  PIN north[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 696.000 72.590 700.000 ;
    END
  END north[20]
  PIN north[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.990 696.000 76.270 700.000 ;
    END
  END north[21]
  PIN north[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 696.000 79.490 700.000 ;
    END
  END north[22]
  PIN north[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 696.000 83.170 700.000 ;
    END
  END north[23]
  PIN north[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 696.000 86.850 700.000 ;
    END
  END north[24]
  PIN north[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 696.000 90.530 700.000 ;
    END
  END north[25]
  PIN north[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 696.000 93.750 700.000 ;
    END
  END north[26]
  PIN north[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 696.000 97.430 700.000 ;
    END
  END north[27]
  PIN north[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 696.000 101.110 700.000 ;
    END
  END north[28]
  PIN north[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 696.000 104.790 700.000 ;
    END
  END north[29]
  PIN north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 696.000 8.650 700.000 ;
    END
  END north[2]
  PIN north[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 107.730 696.000 108.010 700.000 ;
    END
  END north[30]
  PIN north[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 696.000 111.690 700.000 ;
    END
  END north[31]
  PIN north[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 696.000 115.370 700.000 ;
    END
  END north[32]
  PIN north[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 118.310 696.000 118.590 700.000 ;
    END
  END north[33]
  PIN north[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 696.000 122.270 700.000 ;
    END
  END north[34]
  PIN north[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 125.670 696.000 125.950 700.000 ;
    END
  END north[35]
  PIN north[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 129.350 696.000 129.630 700.000 ;
    END
  END north[36]
  PIN north[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 696.000 132.850 700.000 ;
    END
  END north[37]
  PIN north[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 696.000 136.530 700.000 ;
    END
  END north[38]
  PIN north[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 696.000 140.210 700.000 ;
    END
  END north[39]
  PIN north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 696.000 12.330 700.000 ;
    END
  END north[3]
  PIN north[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 696.000 143.890 700.000 ;
    END
  END north[40]
  PIN north[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 146.830 696.000 147.110 700.000 ;
    END
  END north[41]
  PIN north[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 150.510 696.000 150.790 700.000 ;
    END
  END north[42]
  PIN north[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 696.000 154.470 700.000 ;
    END
  END north[43]
  PIN north[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 696.000 157.690 700.000 ;
    END
  END north[44]
  PIN north[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 161.090 696.000 161.370 700.000 ;
    END
  END north[45]
  PIN north[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 164.770 696.000 165.050 700.000 ;
    END
  END north[46]
  PIN north[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 168.450 696.000 168.730 700.000 ;
    END
  END north[47]
  PIN north[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 171.670 696.000 171.950 700.000 ;
    END
  END north[48]
  PIN north[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 175.350 696.000 175.630 700.000 ;
    END
  END north[49]
  PIN north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 696.000 15.550 700.000 ;
    END
  END north[4]
  PIN north[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 179.030 696.000 179.310 700.000 ;
    END
  END north[50]
  PIN north[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 182.710 696.000 182.990 700.000 ;
    END
  END north[51]
  PIN north[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 185.930 696.000 186.210 700.000 ;
    END
  END north[52]
  PIN north[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 696.000 189.890 700.000 ;
    END
  END north[53]
  PIN north[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 696.000 193.570 700.000 ;
    END
  END north[54]
  PIN north[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 196.510 696.000 196.790 700.000 ;
    END
  END north[55]
  PIN north[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 200.190 696.000 200.470 700.000 ;
    END
  END north[56]
  PIN north[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 203.870 696.000 204.150 700.000 ;
    END
  END north[57]
  PIN north[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 207.550 696.000 207.830 700.000 ;
    END
  END north[58]
  PIN north[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 210.770 696.000 211.050 700.000 ;
    END
  END north[59]
  PIN north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 696.000 19.230 700.000 ;
    END
  END north[5]
  PIN north[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 214.450 696.000 214.730 700.000 ;
    END
  END north[60]
  PIN north[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 696.000 218.410 700.000 ;
    END
  END north[61]
  PIN north[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 221.810 696.000 222.090 700.000 ;
    END
  END north[62]
  PIN north[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 225.030 696.000 225.310 700.000 ;
    END
  END north[63]
  PIN north[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 228.710 696.000 228.990 700.000 ;
    END
  END north[64]
  PIN north[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 232.390 696.000 232.670 700.000 ;
    END
  END north[65]
  PIN north[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 235.610 696.000 235.890 700.000 ;
    END
  END north[66]
  PIN north[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 239.290 696.000 239.570 700.000 ;
    END
  END north[67]
  PIN north[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 696.000 243.250 700.000 ;
    END
  END north[68]
  PIN north[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 696.000 246.930 700.000 ;
    END
  END north[69]
  PIN north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 696.000 22.910 700.000 ;
    END
  END north[6]
  PIN north[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 249.870 696.000 250.150 700.000 ;
    END
  END north[70]
  PIN north[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 253.550 696.000 253.830 700.000 ;
    END
  END north[71]
  PIN north[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 257.230 696.000 257.510 700.000 ;
    END
  END north[72]
  PIN north[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 260.450 696.000 260.730 700.000 ;
    END
  END north[73]
  PIN north[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 696.000 264.410 700.000 ;
    END
  END north[74]
  PIN north[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 267.810 696.000 268.090 700.000 ;
    END
  END north[75]
  PIN north[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 271.490 696.000 271.770 700.000 ;
    END
  END north[76]
  PIN north[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 274.710 696.000 274.990 700.000 ;
    END
  END north[77]
  PIN north[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 278.390 696.000 278.670 700.000 ;
    END
  END north[78]
  PIN north[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 282.070 696.000 282.350 700.000 ;
    END
  END north[79]
  PIN north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 696.000 26.590 700.000 ;
    END
  END north[7]
  PIN north[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 285.750 696.000 286.030 700.000 ;
    END
  END north[80]
  PIN north[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 696.000 289.250 700.000 ;
    END
  END north[81]
  PIN north[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 292.650 696.000 292.930 700.000 ;
    END
  END north[82]
  PIN north[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 296.330 696.000 296.610 700.000 ;
    END
  END north[83]
  PIN north[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 299.550 696.000 299.830 700.000 ;
    END
  END north[84]
  PIN north[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 303.230 696.000 303.510 700.000 ;
    END
  END north[85]
  PIN north[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 306.910 696.000 307.190 700.000 ;
    END
  END north[86]
  PIN north[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 310.590 696.000 310.870 700.000 ;
    END
  END north[87]
  PIN north[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 313.810 696.000 314.090 700.000 ;
    END
  END north[88]
  PIN north[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 317.490 696.000 317.770 700.000 ;
    END
  END north[89]
  PIN north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 696.000 29.810 700.000 ;
    END
  END north[8]
  PIN north[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 321.170 696.000 321.450 700.000 ;
    END
  END north[90]
  PIN north[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 696.000 325.130 700.000 ;
    END
  END north[91]
  PIN north[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 328.070 696.000 328.350 700.000 ;
    END
  END north[92]
  PIN north[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 331.750 696.000 332.030 700.000 ;
    END
  END north[93]
  PIN north[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 335.430 696.000 335.710 700.000 ;
    END
  END north[94]
  PIN north[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 338.650 696.000 338.930 700.000 ;
    END
  END north[95]
  PIN north[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 342.330 696.000 342.610 700.000 ;
    END
  END north[96]
  PIN north[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 346.010 696.000 346.290 700.000 ;
    END
  END north[97]
  PIN north[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 696.000 349.970 700.000 ;
    END
  END north[98]
  PIN north[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 352.910 696.000 353.190 700.000 ;
    END
  END north[99]
  PIN north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 696.000 33.490 700.000 ;
    END
  END north[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 696.000 697.040 700.000 697.640 ;
    END
  END rst
  PIN set_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.910 696.000 698.190 700.000 ;
    END
  END set_soft
  PIN shift_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END shift_in
  PIN shift_in_soft
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END shift_in_soft
  PIN shift_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.550 696.000 690.830 700.000 ;
    END
  END shift_out
  PIN south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END south[0]
  PIN south[100]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END south[100]
  PIN south[101]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END south[101]
  PIN south[102]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END south[102]
  PIN south[103]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END south[103]
  PIN south[104]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END south[104]
  PIN south[105]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END south[105]
  PIN south[106]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END south[106]
  PIN south[107]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END south[107]
  PIN south[108]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END south[108]
  PIN south[109]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END south[109]
  PIN south[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END south[10]
  PIN south[110]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END south[110]
  PIN south[111]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END south[111]
  PIN south[112]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END south[112]
  PIN south[113]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END south[113]
  PIN south[114]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END south[114]
  PIN south[115]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END south[115]
  PIN south[116]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END south[116]
  PIN south[117]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END south[117]
  PIN south[118]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END south[118]
  PIN south[119]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END south[119]
  PIN south[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END south[11]
  PIN south[120]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END south[120]
  PIN south[121]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END south[121]
  PIN south[122]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END south[122]
  PIN south[123]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END south[123]
  PIN south[124]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END south[124]
  PIN south[125]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END south[125]
  PIN south[126]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END south[126]
  PIN south[127]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END south[127]
  PIN south[128]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END south[128]
  PIN south[129]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END south[129]
  PIN south[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END south[12]
  PIN south[130]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END south[130]
  PIN south[131]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END south[131]
  PIN south[132]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END south[132]
  PIN south[133]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END south[133]
  PIN south[134]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END south[134]
  PIN south[135]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END south[135]
  PIN south[136]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END south[136]
  PIN south[137]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END south[137]
  PIN south[138]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END south[138]
  PIN south[139]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END south[139]
  PIN south[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END south[13]
  PIN south[140]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END south[140]
  PIN south[141]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END south[141]
  PIN south[142]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END south[142]
  PIN south[143]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END south[143]
  PIN south[144]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END south[144]
  PIN south[145]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END south[145]
  PIN south[146]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END south[146]
  PIN south[147]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END south[147]
  PIN south[148]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END south[148]
  PIN south[149]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END south[149]
  PIN south[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END south[14]
  PIN south[150]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END south[150]
  PIN south[151]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END south[151]
  PIN south[152]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END south[152]
  PIN south[153]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END south[153]
  PIN south[154]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END south[154]
  PIN south[155]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END south[155]
  PIN south[156]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END south[156]
  PIN south[157]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END south[157]
  PIN south[158]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END south[158]
  PIN south[159]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END south[159]
  PIN south[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END south[15]
  PIN south[160]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END south[160]
  PIN south[161]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END south[161]
  PIN south[162]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END south[162]
  PIN south[163]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END south[163]
  PIN south[164]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END south[164]
  PIN south[165]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END south[165]
  PIN south[166]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END south[166]
  PIN south[167]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END south[167]
  PIN south[168]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END south[168]
  PIN south[169]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END south[169]
  PIN south[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END south[16]
  PIN south[170]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END south[170]
  PIN south[171]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END south[171]
  PIN south[172]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END south[172]
  PIN south[173]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END south[173]
  PIN south[174]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END south[174]
  PIN south[175]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END south[175]
  PIN south[176]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END south[176]
  PIN south[177]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END south[177]
  PIN south[178]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END south[178]
  PIN south[179]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END south[179]
  PIN south[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END south[17]
  PIN south[180]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END south[180]
  PIN south[181]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END south[181]
  PIN south[182]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END south[182]
  PIN south[183]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 648.230 0.000 648.510 4.000 ;
    END
  END south[183]
  PIN south[184]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END south[184]
  PIN south[185]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END south[185]
  PIN south[186]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END south[186]
  PIN south[187]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END south[187]
  PIN south[188]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END south[188]
  PIN south[189]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END south[189]
  PIN south[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END south[18]
  PIN south[190]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END south[190]
  PIN south[191]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END south[191]
  PIN south[192]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END south[192]
  PIN south[193]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END south[193]
  PIN south[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END south[19]
  PIN south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END south[1]
  PIN south[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END south[20]
  PIN south[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END south[21]
  PIN south[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END south[22]
  PIN south[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END south[23]
  PIN south[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END south[24]
  PIN south[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END south[25]
  PIN south[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END south[26]
  PIN south[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END south[27]
  PIN south[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END south[28]
  PIN south[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END south[29]
  PIN south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END south[2]
  PIN south[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END south[30]
  PIN south[31]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END south[31]
  PIN south[32]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END south[32]
  PIN south[33]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END south[33]
  PIN south[34]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END south[34]
  PIN south[35]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END south[35]
  PIN south[36]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END south[36]
  PIN south[37]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END south[37]
  PIN south[38]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END south[38]
  PIN south[39]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END south[39]
  PIN south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END south[3]
  PIN south[40]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END south[40]
  PIN south[41]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END south[41]
  PIN south[42]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END south[42]
  PIN south[43]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END south[43]
  PIN south[44]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END south[44]
  PIN south[45]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END south[45]
  PIN south[46]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END south[46]
  PIN south[47]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END south[47]
  PIN south[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END south[48]
  PIN south[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END south[49]
  PIN south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END south[4]
  PIN south[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END south[50]
  PIN south[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END south[51]
  PIN south[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END south[52]
  PIN south[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END south[53]
  PIN south[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END south[54]
  PIN south[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END south[55]
  PIN south[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END south[56]
  PIN south[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END south[57]
  PIN south[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END south[58]
  PIN south[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END south[59]
  PIN south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END south[5]
  PIN south[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END south[60]
  PIN south[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END south[61]
  PIN south[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END south[62]
  PIN south[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END south[63]
  PIN south[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END south[64]
  PIN south[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END south[65]
  PIN south[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END south[66]
  PIN south[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END south[67]
  PIN south[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END south[68]
  PIN south[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END south[69]
  PIN south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END south[6]
  PIN south[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END south[70]
  PIN south[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END south[71]
  PIN south[72]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END south[72]
  PIN south[73]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END south[73]
  PIN south[74]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END south[74]
  PIN south[75]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END south[75]
  PIN south[76]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END south[76]
  PIN south[77]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END south[77]
  PIN south[78]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END south[78]
  PIN south[79]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END south[79]
  PIN south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END south[7]
  PIN south[80]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END south[80]
  PIN south[81]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END south[81]
  PIN south[82]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END south[82]
  PIN south[83]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END south[83]
  PIN south[84]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END south[84]
  PIN south[85]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END south[85]
  PIN south[86]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END south[86]
  PIN south[87]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END south[87]
  PIN south[88]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END south[88]
  PIN south[89]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END south[89]
  PIN south[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END south[8]
  PIN south[90]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END south[90]
  PIN south[91]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END south[91]
  PIN south[92]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END south[92]
  PIN south[93]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END south[93]
  PIN south[94]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END south[94]
  PIN south[95]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END south[95]
  PIN south[96]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END south[96]
  PIN south[97]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END south[97]
  PIN south[98]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END south[98]
  PIN south[99]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END south[99]
  PIN south[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END south[9]
  PIN west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END west[0]
  PIN west[100]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END west[100]
  PIN west[101]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END west[101]
  PIN west[102]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END west[102]
  PIN west[103]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END west[103]
  PIN west[104]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END west[104]
  PIN west[105]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END west[105]
  PIN west[106]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END west[106]
  PIN west[107]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END west[107]
  PIN west[108]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END west[108]
  PIN west[109]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END west[109]
  PIN west[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END west[10]
  PIN west[110]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END west[110]
  PIN west[111]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END west[111]
  PIN west[112]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END west[112]
  PIN west[113]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END west[113]
  PIN west[114]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END west[114]
  PIN west[115]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END west[115]
  PIN west[116]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END west[116]
  PIN west[117]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END west[117]
  PIN west[118]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END west[118]
  PIN west[119]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END west[119]
  PIN west[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END west[11]
  PIN west[120]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END west[120]
  PIN west[121]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END west[121]
  PIN west[122]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END west[122]
  PIN west[123]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END west[123]
  PIN west[124]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END west[124]
  PIN west[125]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END west[125]
  PIN west[126]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END west[126]
  PIN west[127]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END west[127]
  PIN west[128]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END west[128]
  PIN west[129]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END west[129]
  PIN west[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END west[12]
  PIN west[130]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END west[130]
  PIN west[131]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END west[131]
  PIN west[132]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END west[132]
  PIN west[133]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END west[133]
  PIN west[134]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END west[134]
  PIN west[135]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END west[135]
  PIN west[136]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END west[136]
  PIN west[137]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END west[137]
  PIN west[138]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END west[138]
  PIN west[139]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END west[139]
  PIN west[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END west[13]
  PIN west[140]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END west[140]
  PIN west[141]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END west[141]
  PIN west[142]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END west[142]
  PIN west[143]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END west[143]
  PIN west[144]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END west[144]
  PIN west[145]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 521.600 4.000 522.200 ;
    END
  END west[145]
  PIN west[146]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END west[146]
  PIN west[147]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 528.400 4.000 529.000 ;
    END
  END west[147]
  PIN west[148]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END west[148]
  PIN west[149]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END west[149]
  PIN west[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END west[14]
  PIN west[150]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END west[150]
  PIN west[151]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END west[151]
  PIN west[152]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END west[152]
  PIN west[153]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END west[153]
  PIN west[154]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END west[154]
  PIN west[155]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END west[155]
  PIN west[156]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END west[156]
  PIN west[157]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END west[157]
  PIN west[158]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END west[158]
  PIN west[159]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END west[159]
  PIN west[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END west[15]
  PIN west[160]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END west[160]
  PIN west[161]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END west[161]
  PIN west[162]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END west[162]
  PIN west[163]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END west[163]
  PIN west[164]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END west[164]
  PIN west[165]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END west[165]
  PIN west[166]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END west[166]
  PIN west[167]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END west[167]
  PIN west[168]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END west[168]
  PIN west[169]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END west[169]
  PIN west[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END west[16]
  PIN west[170]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END west[170]
  PIN west[171]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END west[171]
  PIN west[172]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END west[172]
  PIN west[173]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END west[173]
  PIN west[174]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END west[174]
  PIN west[175]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END west[175]
  PIN west[176]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END west[176]
  PIN west[177]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END west[177]
  PIN west[178]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END west[178]
  PIN west[179]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END west[179]
  PIN west[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END west[17]
  PIN west[180]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END west[180]
  PIN west[181]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END west[181]
  PIN west[182]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END west[182]
  PIN west[183]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END west[183]
  PIN west[184]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END west[184]
  PIN west[185]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END west[185]
  PIN west[186]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END west[186]
  PIN west[187]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END west[187]
  PIN west[188]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END west[188]
  PIN west[189]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 679.360 4.000 679.960 ;
    END
  END west[189]
  PIN west[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END west[18]
  PIN west[190]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END west[190]
  PIN west[191]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END west[191]
  PIN west[192]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END west[192]
  PIN west[193]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END west[193]
  PIN west[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END west[19]
  PIN west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END west[1]
  PIN west[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END west[20]
  PIN west[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END west[21]
  PIN west[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END west[22]
  PIN west[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END west[23]
  PIN west[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END west[24]
  PIN west[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END west[25]
  PIN west[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END west[26]
  PIN west[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END west[27]
  PIN west[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END west[28]
  PIN west[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END west[29]
  PIN west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END west[2]
  PIN west[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END west[30]
  PIN west[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END west[31]
  PIN west[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END west[32]
  PIN west[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END west[33]
  PIN west[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END west[34]
  PIN west[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END west[35]
  PIN west[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END west[36]
  PIN west[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END west[37]
  PIN west[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END west[38]
  PIN west[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END west[39]
  PIN west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END west[3]
  PIN west[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END west[40]
  PIN west[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END west[41]
  PIN west[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END west[42]
  PIN west[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END west[43]
  PIN west[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END west[44]
  PIN west[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END west[45]
  PIN west[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END west[46]
  PIN west[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END west[47]
  PIN west[48]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END west[48]
  PIN west[49]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END west[49]
  PIN west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END west[4]
  PIN west[50]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END west[50]
  PIN west[51]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END west[51]
  PIN west[52]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END west[52]
  PIN west[53]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END west[53]
  PIN west[54]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END west[54]
  PIN west[55]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END west[55]
  PIN west[56]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END west[56]
  PIN west[57]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END west[57]
  PIN west[58]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END west[58]
  PIN west[59]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END west[59]
  PIN west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END west[5]
  PIN west[60]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END west[60]
  PIN west[61]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END west[61]
  PIN west[62]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END west[62]
  PIN west[63]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END west[63]
  PIN west[64]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END west[64]
  PIN west[65]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END west[65]
  PIN west[66]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END west[66]
  PIN west[67]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END west[67]
  PIN west[68]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END west[68]
  PIN west[69]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END west[69]
  PIN west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END west[6]
  PIN west[70]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END west[70]
  PIN west[71]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END west[71]
  PIN west[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END west[72]
  PIN west[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END west[73]
  PIN west[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END west[74]
  PIN west[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END west[75]
  PIN west[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END west[76]
  PIN west[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END west[77]
  PIN west[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END west[78]
  PIN west[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END west[79]
  PIN west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END west[7]
  PIN west[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END west[80]
  PIN west[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END west[81]
  PIN west[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END west[82]
  PIN west[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END west[83]
  PIN west[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END west[84]
  PIN west[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END west[85]
  PIN west[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END west[86]
  PIN west[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END west[87]
  PIN west[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END west[88]
  PIN west[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END west[89]
  PIN west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END west[8]
  PIN west[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END west[90]
  PIN west[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END west[91]
  PIN west[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END west[92]
  PIN west[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END west[93]
  PIN west[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END west[94]
  PIN west[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END west[95]
  PIN west[96]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END west[96]
  PIN west[97]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END west[97]
  PIN west[98]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END west[98]
  PIN west[99]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END west[99]
  PIN west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END west[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.065 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 0.070 4.800 698.210 690.840 ;
      LAYER met2 ;
        RECT 0.100 695.720 1.190 697.525 ;
        RECT 2.030 695.720 4.410 697.525 ;
        RECT 5.250 695.720 8.090 697.525 ;
        RECT 8.930 695.720 11.770 697.525 ;
        RECT 12.610 695.720 14.990 697.525 ;
        RECT 15.830 695.720 18.670 697.525 ;
        RECT 19.510 695.720 22.350 697.525 ;
        RECT 23.190 695.720 26.030 697.525 ;
        RECT 26.870 695.720 29.250 697.525 ;
        RECT 30.090 695.720 32.930 697.525 ;
        RECT 33.770 695.720 36.610 697.525 ;
        RECT 37.450 695.720 39.830 697.525 ;
        RECT 40.670 695.720 43.510 697.525 ;
        RECT 44.350 695.720 47.190 697.525 ;
        RECT 48.030 695.720 50.870 697.525 ;
        RECT 51.710 695.720 54.090 697.525 ;
        RECT 54.930 695.720 57.770 697.525 ;
        RECT 58.610 695.720 61.450 697.525 ;
        RECT 62.290 695.720 65.130 697.525 ;
        RECT 65.970 695.720 68.350 697.525 ;
        RECT 69.190 695.720 72.030 697.525 ;
        RECT 72.870 695.720 75.710 697.525 ;
        RECT 76.550 695.720 78.930 697.525 ;
        RECT 79.770 695.720 82.610 697.525 ;
        RECT 83.450 695.720 86.290 697.525 ;
        RECT 87.130 695.720 89.970 697.525 ;
        RECT 90.810 695.720 93.190 697.525 ;
        RECT 94.030 695.720 96.870 697.525 ;
        RECT 97.710 695.720 100.550 697.525 ;
        RECT 101.390 695.720 104.230 697.525 ;
        RECT 105.070 695.720 107.450 697.525 ;
        RECT 108.290 695.720 111.130 697.525 ;
        RECT 111.970 695.720 114.810 697.525 ;
        RECT 115.650 695.720 118.030 697.525 ;
        RECT 118.870 695.720 121.710 697.525 ;
        RECT 122.550 695.720 125.390 697.525 ;
        RECT 126.230 695.720 129.070 697.525 ;
        RECT 129.910 695.720 132.290 697.525 ;
        RECT 133.130 695.720 135.970 697.525 ;
        RECT 136.810 695.720 139.650 697.525 ;
        RECT 140.490 695.720 143.330 697.525 ;
        RECT 144.170 695.720 146.550 697.525 ;
        RECT 147.390 695.720 150.230 697.525 ;
        RECT 151.070 695.720 153.910 697.525 ;
        RECT 154.750 695.720 157.130 697.525 ;
        RECT 157.970 695.720 160.810 697.525 ;
        RECT 161.650 695.720 164.490 697.525 ;
        RECT 165.330 695.720 168.170 697.525 ;
        RECT 169.010 695.720 171.390 697.525 ;
        RECT 172.230 695.720 175.070 697.525 ;
        RECT 175.910 695.720 178.750 697.525 ;
        RECT 179.590 695.720 182.430 697.525 ;
        RECT 183.270 695.720 185.650 697.525 ;
        RECT 186.490 695.720 189.330 697.525 ;
        RECT 190.170 695.720 193.010 697.525 ;
        RECT 193.850 695.720 196.230 697.525 ;
        RECT 197.070 695.720 199.910 697.525 ;
        RECT 200.750 695.720 203.590 697.525 ;
        RECT 204.430 695.720 207.270 697.525 ;
        RECT 208.110 695.720 210.490 697.525 ;
        RECT 211.330 695.720 214.170 697.525 ;
        RECT 215.010 695.720 217.850 697.525 ;
        RECT 218.690 695.720 221.530 697.525 ;
        RECT 222.370 695.720 224.750 697.525 ;
        RECT 225.590 695.720 228.430 697.525 ;
        RECT 229.270 695.720 232.110 697.525 ;
        RECT 232.950 695.720 235.330 697.525 ;
        RECT 236.170 695.720 239.010 697.525 ;
        RECT 239.850 695.720 242.690 697.525 ;
        RECT 243.530 695.720 246.370 697.525 ;
        RECT 247.210 695.720 249.590 697.525 ;
        RECT 250.430 695.720 253.270 697.525 ;
        RECT 254.110 695.720 256.950 697.525 ;
        RECT 257.790 695.720 260.170 697.525 ;
        RECT 261.010 695.720 263.850 697.525 ;
        RECT 264.690 695.720 267.530 697.525 ;
        RECT 268.370 695.720 271.210 697.525 ;
        RECT 272.050 695.720 274.430 697.525 ;
        RECT 275.270 695.720 278.110 697.525 ;
        RECT 278.950 695.720 281.790 697.525 ;
        RECT 282.630 695.720 285.470 697.525 ;
        RECT 286.310 695.720 288.690 697.525 ;
        RECT 289.530 695.720 292.370 697.525 ;
        RECT 293.210 695.720 296.050 697.525 ;
        RECT 296.890 695.720 299.270 697.525 ;
        RECT 300.110 695.720 302.950 697.525 ;
        RECT 303.790 695.720 306.630 697.525 ;
        RECT 307.470 695.720 310.310 697.525 ;
        RECT 311.150 695.720 313.530 697.525 ;
        RECT 314.370 695.720 317.210 697.525 ;
        RECT 318.050 695.720 320.890 697.525 ;
        RECT 321.730 695.720 324.570 697.525 ;
        RECT 325.410 695.720 327.790 697.525 ;
        RECT 328.630 695.720 331.470 697.525 ;
        RECT 332.310 695.720 335.150 697.525 ;
        RECT 335.990 695.720 338.370 697.525 ;
        RECT 339.210 695.720 342.050 697.525 ;
        RECT 342.890 695.720 345.730 697.525 ;
        RECT 346.570 695.720 349.410 697.525 ;
        RECT 350.250 695.720 352.630 697.525 ;
        RECT 353.470 695.720 356.310 697.525 ;
        RECT 357.150 695.720 359.990 697.525 ;
        RECT 360.830 695.720 363.670 697.525 ;
        RECT 364.510 695.720 366.890 697.525 ;
        RECT 367.730 695.720 370.570 697.525 ;
        RECT 371.410 695.720 374.250 697.525 ;
        RECT 375.090 695.720 377.470 697.525 ;
        RECT 378.310 695.720 381.150 697.525 ;
        RECT 381.990 695.720 384.830 697.525 ;
        RECT 385.670 695.720 388.510 697.525 ;
        RECT 389.350 695.720 391.730 697.525 ;
        RECT 392.570 695.720 395.410 697.525 ;
        RECT 396.250 695.720 399.090 697.525 ;
        RECT 399.930 695.720 402.770 697.525 ;
        RECT 403.610 695.720 405.990 697.525 ;
        RECT 406.830 695.720 409.670 697.525 ;
        RECT 410.510 695.720 413.350 697.525 ;
        RECT 414.190 695.720 416.570 697.525 ;
        RECT 417.410 695.720 420.250 697.525 ;
        RECT 421.090 695.720 423.930 697.525 ;
        RECT 424.770 695.720 427.610 697.525 ;
        RECT 428.450 695.720 430.830 697.525 ;
        RECT 431.670 695.720 434.510 697.525 ;
        RECT 435.350 695.720 438.190 697.525 ;
        RECT 439.030 695.720 441.870 697.525 ;
        RECT 442.710 695.720 445.090 697.525 ;
        RECT 445.930 695.720 448.770 697.525 ;
        RECT 449.610 695.720 452.450 697.525 ;
        RECT 453.290 695.720 455.670 697.525 ;
        RECT 456.510 695.720 459.350 697.525 ;
        RECT 460.190 695.720 463.030 697.525 ;
        RECT 463.870 695.720 466.710 697.525 ;
        RECT 467.550 695.720 469.930 697.525 ;
        RECT 470.770 695.720 473.610 697.525 ;
        RECT 474.450 695.720 477.290 697.525 ;
        RECT 478.130 695.720 480.510 697.525 ;
        RECT 481.350 695.720 484.190 697.525 ;
        RECT 485.030 695.720 487.870 697.525 ;
        RECT 488.710 695.720 491.550 697.525 ;
        RECT 492.390 695.720 494.770 697.525 ;
        RECT 495.610 695.720 498.450 697.525 ;
        RECT 499.290 695.720 502.130 697.525 ;
        RECT 502.970 695.720 505.810 697.525 ;
        RECT 506.650 695.720 509.030 697.525 ;
        RECT 509.870 695.720 512.710 697.525 ;
        RECT 513.550 695.720 516.390 697.525 ;
        RECT 517.230 695.720 519.610 697.525 ;
        RECT 520.450 695.720 523.290 697.525 ;
        RECT 524.130 695.720 526.970 697.525 ;
        RECT 527.810 695.720 530.650 697.525 ;
        RECT 531.490 695.720 533.870 697.525 ;
        RECT 534.710 695.720 537.550 697.525 ;
        RECT 538.390 695.720 541.230 697.525 ;
        RECT 542.070 695.720 544.910 697.525 ;
        RECT 545.750 695.720 548.130 697.525 ;
        RECT 548.970 695.720 551.810 697.525 ;
        RECT 552.650 695.720 555.490 697.525 ;
        RECT 556.330 695.720 558.710 697.525 ;
        RECT 559.550 695.720 562.390 697.525 ;
        RECT 563.230 695.720 566.070 697.525 ;
        RECT 566.910 695.720 569.750 697.525 ;
        RECT 570.590 695.720 572.970 697.525 ;
        RECT 573.810 695.720 576.650 697.525 ;
        RECT 577.490 695.720 580.330 697.525 ;
        RECT 581.170 695.720 584.010 697.525 ;
        RECT 584.850 695.720 587.230 697.525 ;
        RECT 588.070 695.720 590.910 697.525 ;
        RECT 591.750 695.720 594.590 697.525 ;
        RECT 595.430 695.720 597.810 697.525 ;
        RECT 598.650 695.720 601.490 697.525 ;
        RECT 602.330 695.720 605.170 697.525 ;
        RECT 606.010 695.720 608.850 697.525 ;
        RECT 609.690 695.720 612.070 697.525 ;
        RECT 612.910 695.720 615.750 697.525 ;
        RECT 616.590 695.720 619.430 697.525 ;
        RECT 620.270 695.720 623.110 697.525 ;
        RECT 623.950 695.720 626.330 697.525 ;
        RECT 627.170 695.720 630.010 697.525 ;
        RECT 630.850 695.720 633.690 697.525 ;
        RECT 634.530 695.720 636.910 697.525 ;
        RECT 637.750 695.720 640.590 697.525 ;
        RECT 641.430 695.720 644.270 697.525 ;
        RECT 645.110 695.720 647.950 697.525 ;
        RECT 648.790 695.720 651.170 697.525 ;
        RECT 652.010 695.720 654.850 697.525 ;
        RECT 655.690 695.720 658.530 697.525 ;
        RECT 659.370 695.720 662.210 697.525 ;
        RECT 663.050 695.720 665.430 697.525 ;
        RECT 666.270 695.720 669.110 697.525 ;
        RECT 669.950 695.720 672.790 697.525 ;
        RECT 673.630 695.720 676.010 697.525 ;
        RECT 676.850 695.720 679.690 697.525 ;
        RECT 680.530 695.720 683.370 697.525 ;
        RECT 684.210 695.720 687.050 697.525 ;
        RECT 687.890 695.720 690.270 697.525 ;
        RECT 691.110 695.720 693.950 697.525 ;
        RECT 694.790 695.720 697.630 697.525 ;
        RECT 0.100 4.280 698.180 695.720 ;
        RECT 0.100 1.515 1.190 4.280 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 8.090 4.280 ;
        RECT 8.930 1.515 11.770 4.280 ;
        RECT 12.610 1.515 14.990 4.280 ;
        RECT 15.830 1.515 18.670 4.280 ;
        RECT 19.510 1.515 22.350 4.280 ;
        RECT 23.190 1.515 25.570 4.280 ;
        RECT 26.410 1.515 29.250 4.280 ;
        RECT 30.090 1.515 32.930 4.280 ;
        RECT 33.770 1.515 36.150 4.280 ;
        RECT 36.990 1.515 39.830 4.280 ;
        RECT 40.670 1.515 43.510 4.280 ;
        RECT 44.350 1.515 46.730 4.280 ;
        RECT 47.570 1.515 50.410 4.280 ;
        RECT 51.250 1.515 54.090 4.280 ;
        RECT 54.930 1.515 57.310 4.280 ;
        RECT 58.150 1.515 60.990 4.280 ;
        RECT 61.830 1.515 64.670 4.280 ;
        RECT 65.510 1.515 68.350 4.280 ;
        RECT 69.190 1.515 71.570 4.280 ;
        RECT 72.410 1.515 75.250 4.280 ;
        RECT 76.090 1.515 78.930 4.280 ;
        RECT 79.770 1.515 82.150 4.280 ;
        RECT 82.990 1.515 85.830 4.280 ;
        RECT 86.670 1.515 89.510 4.280 ;
        RECT 90.350 1.515 92.730 4.280 ;
        RECT 93.570 1.515 96.410 4.280 ;
        RECT 97.250 1.515 100.090 4.280 ;
        RECT 100.930 1.515 103.310 4.280 ;
        RECT 104.150 1.515 106.990 4.280 ;
        RECT 107.830 1.515 110.670 4.280 ;
        RECT 111.510 1.515 113.890 4.280 ;
        RECT 114.730 1.515 117.570 4.280 ;
        RECT 118.410 1.515 121.250 4.280 ;
        RECT 122.090 1.515 124.930 4.280 ;
        RECT 125.770 1.515 128.150 4.280 ;
        RECT 128.990 1.515 131.830 4.280 ;
        RECT 132.670 1.515 135.510 4.280 ;
        RECT 136.350 1.515 138.730 4.280 ;
        RECT 139.570 1.515 142.410 4.280 ;
        RECT 143.250 1.515 146.090 4.280 ;
        RECT 146.930 1.515 149.310 4.280 ;
        RECT 150.150 1.515 152.990 4.280 ;
        RECT 153.830 1.515 156.670 4.280 ;
        RECT 157.510 1.515 159.890 4.280 ;
        RECT 160.730 1.515 163.570 4.280 ;
        RECT 164.410 1.515 167.250 4.280 ;
        RECT 168.090 1.515 170.470 4.280 ;
        RECT 171.310 1.515 174.150 4.280 ;
        RECT 174.990 1.515 177.830 4.280 ;
        RECT 178.670 1.515 181.510 4.280 ;
        RECT 182.350 1.515 184.730 4.280 ;
        RECT 185.570 1.515 188.410 4.280 ;
        RECT 189.250 1.515 192.090 4.280 ;
        RECT 192.930 1.515 195.310 4.280 ;
        RECT 196.150 1.515 198.990 4.280 ;
        RECT 199.830 1.515 202.670 4.280 ;
        RECT 203.510 1.515 205.890 4.280 ;
        RECT 206.730 1.515 209.570 4.280 ;
        RECT 210.410 1.515 213.250 4.280 ;
        RECT 214.090 1.515 216.470 4.280 ;
        RECT 217.310 1.515 220.150 4.280 ;
        RECT 220.990 1.515 223.830 4.280 ;
        RECT 224.670 1.515 227.050 4.280 ;
        RECT 227.890 1.515 230.730 4.280 ;
        RECT 231.570 1.515 234.410 4.280 ;
        RECT 235.250 1.515 238.090 4.280 ;
        RECT 238.930 1.515 241.310 4.280 ;
        RECT 242.150 1.515 244.990 4.280 ;
        RECT 245.830 1.515 248.670 4.280 ;
        RECT 249.510 1.515 251.890 4.280 ;
        RECT 252.730 1.515 255.570 4.280 ;
        RECT 256.410 1.515 259.250 4.280 ;
        RECT 260.090 1.515 262.470 4.280 ;
        RECT 263.310 1.515 266.150 4.280 ;
        RECT 266.990 1.515 269.830 4.280 ;
        RECT 270.670 1.515 273.050 4.280 ;
        RECT 273.890 1.515 276.730 4.280 ;
        RECT 277.570 1.515 280.410 4.280 ;
        RECT 281.250 1.515 283.630 4.280 ;
        RECT 284.470 1.515 287.310 4.280 ;
        RECT 288.150 1.515 290.990 4.280 ;
        RECT 291.830 1.515 294.670 4.280 ;
        RECT 295.510 1.515 297.890 4.280 ;
        RECT 298.730 1.515 301.570 4.280 ;
        RECT 302.410 1.515 305.250 4.280 ;
        RECT 306.090 1.515 308.470 4.280 ;
        RECT 309.310 1.515 312.150 4.280 ;
        RECT 312.990 1.515 315.830 4.280 ;
        RECT 316.670 1.515 319.050 4.280 ;
        RECT 319.890 1.515 322.730 4.280 ;
        RECT 323.570 1.515 326.410 4.280 ;
        RECT 327.250 1.515 329.630 4.280 ;
        RECT 330.470 1.515 333.310 4.280 ;
        RECT 334.150 1.515 336.990 4.280 ;
        RECT 337.830 1.515 340.210 4.280 ;
        RECT 341.050 1.515 343.890 4.280 ;
        RECT 344.730 1.515 347.570 4.280 ;
        RECT 348.410 1.515 351.250 4.280 ;
        RECT 352.090 1.515 354.470 4.280 ;
        RECT 355.310 1.515 358.150 4.280 ;
        RECT 358.990 1.515 361.830 4.280 ;
        RECT 362.670 1.515 365.050 4.280 ;
        RECT 365.890 1.515 368.730 4.280 ;
        RECT 369.570 1.515 372.410 4.280 ;
        RECT 373.250 1.515 375.630 4.280 ;
        RECT 376.470 1.515 379.310 4.280 ;
        RECT 380.150 1.515 382.990 4.280 ;
        RECT 383.830 1.515 386.210 4.280 ;
        RECT 387.050 1.515 389.890 4.280 ;
        RECT 390.730 1.515 393.570 4.280 ;
        RECT 394.410 1.515 396.790 4.280 ;
        RECT 397.630 1.515 400.470 4.280 ;
        RECT 401.310 1.515 404.150 4.280 ;
        RECT 404.990 1.515 407.370 4.280 ;
        RECT 408.210 1.515 411.050 4.280 ;
        RECT 411.890 1.515 414.730 4.280 ;
        RECT 415.570 1.515 418.410 4.280 ;
        RECT 419.250 1.515 421.630 4.280 ;
        RECT 422.470 1.515 425.310 4.280 ;
        RECT 426.150 1.515 428.990 4.280 ;
        RECT 429.830 1.515 432.210 4.280 ;
        RECT 433.050 1.515 435.890 4.280 ;
        RECT 436.730 1.515 439.570 4.280 ;
        RECT 440.410 1.515 442.790 4.280 ;
        RECT 443.630 1.515 446.470 4.280 ;
        RECT 447.310 1.515 450.150 4.280 ;
        RECT 450.990 1.515 453.370 4.280 ;
        RECT 454.210 1.515 457.050 4.280 ;
        RECT 457.890 1.515 460.730 4.280 ;
        RECT 461.570 1.515 463.950 4.280 ;
        RECT 464.790 1.515 467.630 4.280 ;
        RECT 468.470 1.515 471.310 4.280 ;
        RECT 472.150 1.515 474.990 4.280 ;
        RECT 475.830 1.515 478.210 4.280 ;
        RECT 479.050 1.515 481.890 4.280 ;
        RECT 482.730 1.515 485.570 4.280 ;
        RECT 486.410 1.515 488.790 4.280 ;
        RECT 489.630 1.515 492.470 4.280 ;
        RECT 493.310 1.515 496.150 4.280 ;
        RECT 496.990 1.515 499.370 4.280 ;
        RECT 500.210 1.515 503.050 4.280 ;
        RECT 503.890 1.515 506.730 4.280 ;
        RECT 507.570 1.515 509.950 4.280 ;
        RECT 510.790 1.515 513.630 4.280 ;
        RECT 514.470 1.515 517.310 4.280 ;
        RECT 518.150 1.515 520.530 4.280 ;
        RECT 521.370 1.515 524.210 4.280 ;
        RECT 525.050 1.515 527.890 4.280 ;
        RECT 528.730 1.515 531.570 4.280 ;
        RECT 532.410 1.515 534.790 4.280 ;
        RECT 535.630 1.515 538.470 4.280 ;
        RECT 539.310 1.515 542.150 4.280 ;
        RECT 542.990 1.515 545.370 4.280 ;
        RECT 546.210 1.515 549.050 4.280 ;
        RECT 549.890 1.515 552.730 4.280 ;
        RECT 553.570 1.515 555.950 4.280 ;
        RECT 556.790 1.515 559.630 4.280 ;
        RECT 560.470 1.515 563.310 4.280 ;
        RECT 564.150 1.515 566.530 4.280 ;
        RECT 567.370 1.515 570.210 4.280 ;
        RECT 571.050 1.515 573.890 4.280 ;
        RECT 574.730 1.515 577.110 4.280 ;
        RECT 577.950 1.515 580.790 4.280 ;
        RECT 581.630 1.515 584.470 4.280 ;
        RECT 585.310 1.515 588.150 4.280 ;
        RECT 588.990 1.515 591.370 4.280 ;
        RECT 592.210 1.515 595.050 4.280 ;
        RECT 595.890 1.515 598.730 4.280 ;
        RECT 599.570 1.515 601.950 4.280 ;
        RECT 602.790 1.515 605.630 4.280 ;
        RECT 606.470 1.515 609.310 4.280 ;
        RECT 610.150 1.515 612.530 4.280 ;
        RECT 613.370 1.515 616.210 4.280 ;
        RECT 617.050 1.515 619.890 4.280 ;
        RECT 620.730 1.515 623.110 4.280 ;
        RECT 623.950 1.515 626.790 4.280 ;
        RECT 627.630 1.515 630.470 4.280 ;
        RECT 631.310 1.515 633.690 4.280 ;
        RECT 634.530 1.515 637.370 4.280 ;
        RECT 638.210 1.515 641.050 4.280 ;
        RECT 641.890 1.515 644.730 4.280 ;
        RECT 645.570 1.515 647.950 4.280 ;
        RECT 648.790 1.515 651.630 4.280 ;
        RECT 652.470 1.515 655.310 4.280 ;
        RECT 656.150 1.515 658.530 4.280 ;
        RECT 659.370 1.515 662.210 4.280 ;
        RECT 663.050 1.515 665.890 4.280 ;
        RECT 666.730 1.515 669.110 4.280 ;
        RECT 669.950 1.515 672.790 4.280 ;
        RECT 673.630 1.515 676.470 4.280 ;
        RECT 677.310 1.515 679.690 4.280 ;
        RECT 680.530 1.515 683.370 4.280 ;
        RECT 684.210 1.515 687.050 4.280 ;
        RECT 687.890 1.515 690.270 4.280 ;
        RECT 691.110 1.515 693.950 4.280 ;
        RECT 694.790 1.515 697.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 696.640 695.600 697.505 ;
        RECT 4.000 694.640 696.130 696.640 ;
        RECT 4.400 693.240 695.600 694.640 ;
        RECT 4.000 691.240 696.130 693.240 ;
        RECT 4.400 689.840 695.600 691.240 ;
        RECT 4.000 687.160 696.130 689.840 ;
        RECT 4.400 685.760 695.600 687.160 ;
        RECT 4.000 683.760 696.130 685.760 ;
        RECT 4.400 682.360 695.600 683.760 ;
        RECT 4.000 680.360 696.130 682.360 ;
        RECT 4.400 678.960 695.600 680.360 ;
        RECT 4.000 676.960 696.130 678.960 ;
        RECT 4.400 675.560 695.600 676.960 ;
        RECT 4.000 672.880 696.130 675.560 ;
        RECT 4.400 671.480 695.600 672.880 ;
        RECT 4.000 669.480 696.130 671.480 ;
        RECT 4.400 668.080 695.600 669.480 ;
        RECT 4.000 666.080 696.130 668.080 ;
        RECT 4.400 664.680 695.600 666.080 ;
        RECT 4.000 662.000 696.130 664.680 ;
        RECT 4.400 660.600 695.600 662.000 ;
        RECT 4.000 658.600 696.130 660.600 ;
        RECT 4.400 657.200 695.600 658.600 ;
        RECT 4.000 655.200 696.130 657.200 ;
        RECT 4.400 653.800 695.600 655.200 ;
        RECT 4.000 651.800 696.130 653.800 ;
        RECT 4.400 650.400 695.600 651.800 ;
        RECT 4.000 647.720 696.130 650.400 ;
        RECT 4.400 646.320 695.600 647.720 ;
        RECT 4.000 644.320 696.130 646.320 ;
        RECT 4.400 642.920 695.600 644.320 ;
        RECT 4.000 640.920 696.130 642.920 ;
        RECT 4.400 639.520 695.600 640.920 ;
        RECT 4.000 637.520 696.130 639.520 ;
        RECT 4.400 636.120 695.600 637.520 ;
        RECT 4.000 633.440 696.130 636.120 ;
        RECT 4.400 632.040 695.600 633.440 ;
        RECT 4.000 630.040 696.130 632.040 ;
        RECT 4.400 628.640 695.600 630.040 ;
        RECT 4.000 626.640 696.130 628.640 ;
        RECT 4.400 625.240 695.600 626.640 ;
        RECT 4.000 622.560 696.130 625.240 ;
        RECT 4.400 621.160 695.600 622.560 ;
        RECT 4.000 619.160 696.130 621.160 ;
        RECT 4.400 617.760 695.600 619.160 ;
        RECT 4.000 615.760 696.130 617.760 ;
        RECT 4.400 614.360 695.600 615.760 ;
        RECT 4.000 612.360 696.130 614.360 ;
        RECT 4.400 610.960 695.600 612.360 ;
        RECT 4.000 608.280 696.130 610.960 ;
        RECT 4.400 606.880 695.600 608.280 ;
        RECT 4.000 604.880 696.130 606.880 ;
        RECT 4.400 603.480 695.600 604.880 ;
        RECT 4.000 601.480 696.130 603.480 ;
        RECT 4.400 600.080 695.600 601.480 ;
        RECT 4.000 597.400 696.130 600.080 ;
        RECT 4.400 596.000 695.600 597.400 ;
        RECT 4.000 594.000 696.130 596.000 ;
        RECT 4.400 592.600 695.600 594.000 ;
        RECT 4.000 590.600 696.130 592.600 ;
        RECT 4.400 589.200 695.600 590.600 ;
        RECT 4.000 587.200 696.130 589.200 ;
        RECT 4.400 585.800 695.600 587.200 ;
        RECT 4.000 583.120 696.130 585.800 ;
        RECT 4.400 581.720 695.600 583.120 ;
        RECT 4.000 579.720 696.130 581.720 ;
        RECT 4.400 578.320 695.600 579.720 ;
        RECT 4.000 576.320 696.130 578.320 ;
        RECT 4.400 574.920 695.600 576.320 ;
        RECT 4.000 572.920 696.130 574.920 ;
        RECT 4.400 571.520 695.600 572.920 ;
        RECT 4.000 568.840 696.130 571.520 ;
        RECT 4.400 567.440 695.600 568.840 ;
        RECT 4.000 565.440 696.130 567.440 ;
        RECT 4.400 564.040 695.600 565.440 ;
        RECT 4.000 562.040 696.130 564.040 ;
        RECT 4.400 560.640 695.600 562.040 ;
        RECT 4.000 557.960 696.130 560.640 ;
        RECT 4.400 556.560 695.600 557.960 ;
        RECT 4.000 554.560 696.130 556.560 ;
        RECT 4.400 553.160 695.600 554.560 ;
        RECT 4.000 551.160 696.130 553.160 ;
        RECT 4.400 549.760 695.600 551.160 ;
        RECT 4.000 547.760 696.130 549.760 ;
        RECT 4.400 546.360 695.600 547.760 ;
        RECT 4.000 543.680 696.130 546.360 ;
        RECT 4.400 542.280 695.600 543.680 ;
        RECT 4.000 540.280 696.130 542.280 ;
        RECT 4.400 538.880 695.600 540.280 ;
        RECT 4.000 536.880 696.130 538.880 ;
        RECT 4.400 535.480 695.600 536.880 ;
        RECT 4.000 532.800 696.130 535.480 ;
        RECT 4.400 531.400 695.600 532.800 ;
        RECT 4.000 529.400 696.130 531.400 ;
        RECT 4.400 528.000 695.600 529.400 ;
        RECT 4.000 526.000 696.130 528.000 ;
        RECT 4.400 524.600 695.600 526.000 ;
        RECT 4.000 522.600 696.130 524.600 ;
        RECT 4.400 521.200 695.600 522.600 ;
        RECT 4.000 518.520 696.130 521.200 ;
        RECT 4.400 517.120 695.600 518.520 ;
        RECT 4.000 515.120 696.130 517.120 ;
        RECT 4.400 513.720 695.600 515.120 ;
        RECT 4.000 511.720 696.130 513.720 ;
        RECT 4.400 510.320 695.600 511.720 ;
        RECT 4.000 508.320 696.130 510.320 ;
        RECT 4.400 506.920 695.600 508.320 ;
        RECT 4.000 504.240 696.130 506.920 ;
        RECT 4.400 502.840 695.600 504.240 ;
        RECT 4.000 500.840 696.130 502.840 ;
        RECT 4.400 499.440 695.600 500.840 ;
        RECT 4.000 497.440 696.130 499.440 ;
        RECT 4.400 496.040 695.600 497.440 ;
        RECT 4.000 493.360 696.130 496.040 ;
        RECT 4.400 491.960 695.600 493.360 ;
        RECT 4.000 489.960 696.130 491.960 ;
        RECT 4.400 488.560 695.600 489.960 ;
        RECT 4.000 486.560 696.130 488.560 ;
        RECT 4.400 485.160 695.600 486.560 ;
        RECT 4.000 483.160 696.130 485.160 ;
        RECT 4.400 481.760 695.600 483.160 ;
        RECT 4.000 479.080 696.130 481.760 ;
        RECT 4.400 477.680 695.600 479.080 ;
        RECT 4.000 475.680 696.130 477.680 ;
        RECT 4.400 474.280 695.600 475.680 ;
        RECT 4.000 472.280 696.130 474.280 ;
        RECT 4.400 470.880 695.600 472.280 ;
        RECT 4.000 468.880 696.130 470.880 ;
        RECT 4.400 467.480 695.600 468.880 ;
        RECT 4.000 464.800 696.130 467.480 ;
        RECT 4.400 463.400 695.600 464.800 ;
        RECT 4.000 461.400 696.130 463.400 ;
        RECT 4.400 460.000 695.600 461.400 ;
        RECT 4.000 458.000 696.130 460.000 ;
        RECT 4.400 456.600 695.600 458.000 ;
        RECT 4.000 453.920 696.130 456.600 ;
        RECT 4.400 452.520 695.600 453.920 ;
        RECT 4.000 450.520 696.130 452.520 ;
        RECT 4.400 449.120 695.600 450.520 ;
        RECT 4.000 447.120 696.130 449.120 ;
        RECT 4.400 445.720 695.600 447.120 ;
        RECT 4.000 443.720 696.130 445.720 ;
        RECT 4.400 442.320 695.600 443.720 ;
        RECT 4.000 439.640 696.130 442.320 ;
        RECT 4.400 438.240 695.600 439.640 ;
        RECT 4.000 436.240 696.130 438.240 ;
        RECT 4.400 434.840 695.600 436.240 ;
        RECT 4.000 432.840 696.130 434.840 ;
        RECT 4.400 431.440 695.600 432.840 ;
        RECT 4.000 428.760 696.130 431.440 ;
        RECT 4.400 427.360 695.600 428.760 ;
        RECT 4.000 425.360 696.130 427.360 ;
        RECT 4.400 423.960 695.600 425.360 ;
        RECT 4.000 421.960 696.130 423.960 ;
        RECT 4.400 420.560 695.600 421.960 ;
        RECT 4.000 418.560 696.130 420.560 ;
        RECT 4.400 417.160 695.600 418.560 ;
        RECT 4.000 414.480 696.130 417.160 ;
        RECT 4.400 413.080 695.600 414.480 ;
        RECT 4.000 411.080 696.130 413.080 ;
        RECT 4.400 409.680 695.600 411.080 ;
        RECT 4.000 407.680 696.130 409.680 ;
        RECT 4.400 406.280 695.600 407.680 ;
        RECT 4.000 404.280 696.130 406.280 ;
        RECT 4.400 402.880 695.600 404.280 ;
        RECT 4.000 400.200 696.130 402.880 ;
        RECT 4.400 398.800 695.600 400.200 ;
        RECT 4.000 396.800 696.130 398.800 ;
        RECT 4.400 395.400 695.600 396.800 ;
        RECT 4.000 393.400 696.130 395.400 ;
        RECT 4.400 392.000 695.600 393.400 ;
        RECT 4.000 389.320 696.130 392.000 ;
        RECT 4.400 387.920 695.600 389.320 ;
        RECT 4.000 385.920 696.130 387.920 ;
        RECT 4.400 384.520 695.600 385.920 ;
        RECT 4.000 382.520 696.130 384.520 ;
        RECT 4.400 381.120 695.600 382.520 ;
        RECT 4.000 379.120 696.130 381.120 ;
        RECT 4.400 377.720 695.600 379.120 ;
        RECT 4.000 375.040 696.130 377.720 ;
        RECT 4.400 373.640 695.600 375.040 ;
        RECT 4.000 371.640 696.130 373.640 ;
        RECT 4.400 370.240 695.600 371.640 ;
        RECT 4.000 368.240 696.130 370.240 ;
        RECT 4.400 366.840 695.600 368.240 ;
        RECT 4.000 364.160 696.130 366.840 ;
        RECT 4.400 362.760 695.600 364.160 ;
        RECT 4.000 360.760 696.130 362.760 ;
        RECT 4.400 359.360 695.600 360.760 ;
        RECT 4.000 357.360 696.130 359.360 ;
        RECT 4.400 355.960 695.600 357.360 ;
        RECT 4.000 353.960 696.130 355.960 ;
        RECT 4.400 352.560 695.600 353.960 ;
        RECT 4.000 349.880 696.130 352.560 ;
        RECT 4.400 348.480 695.600 349.880 ;
        RECT 4.000 346.480 696.130 348.480 ;
        RECT 4.400 345.080 695.600 346.480 ;
        RECT 4.000 343.080 696.130 345.080 ;
        RECT 4.400 341.680 695.600 343.080 ;
        RECT 4.000 339.680 696.130 341.680 ;
        RECT 4.400 338.280 695.600 339.680 ;
        RECT 4.000 335.600 696.130 338.280 ;
        RECT 4.400 334.200 695.600 335.600 ;
        RECT 4.000 332.200 696.130 334.200 ;
        RECT 4.400 330.800 695.600 332.200 ;
        RECT 4.000 328.800 696.130 330.800 ;
        RECT 4.400 327.400 695.600 328.800 ;
        RECT 4.000 324.720 696.130 327.400 ;
        RECT 4.400 323.320 695.600 324.720 ;
        RECT 4.000 321.320 696.130 323.320 ;
        RECT 4.400 319.920 695.600 321.320 ;
        RECT 4.000 317.920 696.130 319.920 ;
        RECT 4.400 316.520 695.600 317.920 ;
        RECT 4.000 314.520 696.130 316.520 ;
        RECT 4.400 313.120 695.600 314.520 ;
        RECT 4.000 310.440 696.130 313.120 ;
        RECT 4.400 309.040 695.600 310.440 ;
        RECT 4.000 307.040 696.130 309.040 ;
        RECT 4.400 305.640 695.600 307.040 ;
        RECT 4.000 303.640 696.130 305.640 ;
        RECT 4.400 302.240 695.600 303.640 ;
        RECT 4.000 299.560 696.130 302.240 ;
        RECT 4.400 298.160 695.600 299.560 ;
        RECT 4.000 296.160 696.130 298.160 ;
        RECT 4.400 294.760 695.600 296.160 ;
        RECT 4.000 292.760 696.130 294.760 ;
        RECT 4.400 291.360 695.600 292.760 ;
        RECT 4.000 289.360 696.130 291.360 ;
        RECT 4.400 287.960 695.600 289.360 ;
        RECT 4.000 285.280 696.130 287.960 ;
        RECT 4.400 283.880 695.600 285.280 ;
        RECT 4.000 281.880 696.130 283.880 ;
        RECT 4.400 280.480 695.600 281.880 ;
        RECT 4.000 278.480 696.130 280.480 ;
        RECT 4.400 277.080 695.600 278.480 ;
        RECT 4.000 275.080 696.130 277.080 ;
        RECT 4.400 273.680 695.600 275.080 ;
        RECT 4.000 271.000 696.130 273.680 ;
        RECT 4.400 269.600 695.600 271.000 ;
        RECT 4.000 267.600 696.130 269.600 ;
        RECT 4.400 266.200 695.600 267.600 ;
        RECT 4.000 264.200 696.130 266.200 ;
        RECT 4.400 262.800 695.600 264.200 ;
        RECT 4.000 260.120 696.130 262.800 ;
        RECT 4.400 258.720 695.600 260.120 ;
        RECT 4.000 256.720 696.130 258.720 ;
        RECT 4.400 255.320 695.600 256.720 ;
        RECT 4.000 253.320 696.130 255.320 ;
        RECT 4.400 251.920 695.600 253.320 ;
        RECT 4.000 249.920 696.130 251.920 ;
        RECT 4.400 248.520 695.600 249.920 ;
        RECT 4.000 245.840 696.130 248.520 ;
        RECT 4.400 244.440 695.600 245.840 ;
        RECT 4.000 242.440 696.130 244.440 ;
        RECT 4.400 241.040 695.600 242.440 ;
        RECT 4.000 239.040 696.130 241.040 ;
        RECT 4.400 237.640 695.600 239.040 ;
        RECT 4.000 235.640 696.130 237.640 ;
        RECT 4.400 234.240 695.600 235.640 ;
        RECT 4.000 231.560 696.130 234.240 ;
        RECT 4.400 230.160 695.600 231.560 ;
        RECT 4.000 228.160 696.130 230.160 ;
        RECT 4.400 226.760 695.600 228.160 ;
        RECT 4.000 224.760 696.130 226.760 ;
        RECT 4.400 223.360 695.600 224.760 ;
        RECT 4.000 220.680 696.130 223.360 ;
        RECT 4.400 219.280 695.600 220.680 ;
        RECT 4.000 217.280 696.130 219.280 ;
        RECT 4.400 215.880 695.600 217.280 ;
        RECT 4.000 213.880 696.130 215.880 ;
        RECT 4.400 212.480 695.600 213.880 ;
        RECT 4.000 210.480 696.130 212.480 ;
        RECT 4.400 209.080 695.600 210.480 ;
        RECT 4.000 206.400 696.130 209.080 ;
        RECT 4.400 205.000 695.600 206.400 ;
        RECT 4.000 203.000 696.130 205.000 ;
        RECT 4.400 201.600 695.600 203.000 ;
        RECT 4.000 199.600 696.130 201.600 ;
        RECT 4.400 198.200 695.600 199.600 ;
        RECT 4.000 195.520 696.130 198.200 ;
        RECT 4.400 194.120 695.600 195.520 ;
        RECT 4.000 192.120 696.130 194.120 ;
        RECT 4.400 190.720 695.600 192.120 ;
        RECT 4.000 188.720 696.130 190.720 ;
        RECT 4.400 187.320 695.600 188.720 ;
        RECT 4.000 185.320 696.130 187.320 ;
        RECT 4.400 183.920 695.600 185.320 ;
        RECT 4.000 181.240 696.130 183.920 ;
        RECT 4.400 179.840 695.600 181.240 ;
        RECT 4.000 177.840 696.130 179.840 ;
        RECT 4.400 176.440 695.600 177.840 ;
        RECT 4.000 174.440 696.130 176.440 ;
        RECT 4.400 173.040 695.600 174.440 ;
        RECT 4.000 171.040 696.130 173.040 ;
        RECT 4.400 169.640 695.600 171.040 ;
        RECT 4.000 166.960 696.130 169.640 ;
        RECT 4.400 165.560 695.600 166.960 ;
        RECT 4.000 163.560 696.130 165.560 ;
        RECT 4.400 162.160 695.600 163.560 ;
        RECT 4.000 160.160 696.130 162.160 ;
        RECT 4.400 158.760 695.600 160.160 ;
        RECT 4.000 156.080 696.130 158.760 ;
        RECT 4.400 154.680 695.600 156.080 ;
        RECT 4.000 152.680 696.130 154.680 ;
        RECT 4.400 151.280 695.600 152.680 ;
        RECT 4.000 149.280 696.130 151.280 ;
        RECT 4.400 147.880 695.600 149.280 ;
        RECT 4.000 145.880 696.130 147.880 ;
        RECT 4.400 144.480 695.600 145.880 ;
        RECT 4.000 141.800 696.130 144.480 ;
        RECT 4.400 140.400 695.600 141.800 ;
        RECT 4.000 138.400 696.130 140.400 ;
        RECT 4.400 137.000 695.600 138.400 ;
        RECT 4.000 135.000 696.130 137.000 ;
        RECT 4.400 133.600 695.600 135.000 ;
        RECT 4.000 130.920 696.130 133.600 ;
        RECT 4.400 129.520 695.600 130.920 ;
        RECT 4.000 127.520 696.130 129.520 ;
        RECT 4.400 126.120 695.600 127.520 ;
        RECT 4.000 124.120 696.130 126.120 ;
        RECT 4.400 122.720 695.600 124.120 ;
        RECT 4.000 120.720 696.130 122.720 ;
        RECT 4.400 119.320 695.600 120.720 ;
        RECT 4.000 116.640 696.130 119.320 ;
        RECT 4.400 115.240 695.600 116.640 ;
        RECT 4.000 113.240 696.130 115.240 ;
        RECT 4.400 111.840 695.600 113.240 ;
        RECT 4.000 109.840 696.130 111.840 ;
        RECT 4.400 108.440 695.600 109.840 ;
        RECT 4.000 106.440 696.130 108.440 ;
        RECT 4.400 105.040 695.600 106.440 ;
        RECT 4.000 102.360 696.130 105.040 ;
        RECT 4.400 100.960 695.600 102.360 ;
        RECT 4.000 98.960 696.130 100.960 ;
        RECT 4.400 97.560 695.600 98.960 ;
        RECT 4.000 95.560 696.130 97.560 ;
        RECT 4.400 94.160 695.600 95.560 ;
        RECT 4.000 91.480 696.130 94.160 ;
        RECT 4.400 90.080 695.600 91.480 ;
        RECT 4.000 88.080 696.130 90.080 ;
        RECT 4.400 86.680 695.600 88.080 ;
        RECT 4.000 84.680 696.130 86.680 ;
        RECT 4.400 83.280 695.600 84.680 ;
        RECT 4.000 81.280 696.130 83.280 ;
        RECT 4.400 79.880 695.600 81.280 ;
        RECT 4.000 77.200 696.130 79.880 ;
        RECT 4.400 75.800 695.600 77.200 ;
        RECT 4.000 73.800 696.130 75.800 ;
        RECT 4.400 72.400 695.600 73.800 ;
        RECT 4.000 70.400 696.130 72.400 ;
        RECT 4.400 69.000 695.600 70.400 ;
        RECT 4.000 66.320 696.130 69.000 ;
        RECT 4.400 64.920 695.600 66.320 ;
        RECT 4.000 62.920 696.130 64.920 ;
        RECT 4.400 61.520 695.600 62.920 ;
        RECT 4.000 59.520 696.130 61.520 ;
        RECT 4.400 58.120 695.600 59.520 ;
        RECT 4.000 56.120 696.130 58.120 ;
        RECT 4.400 54.720 695.600 56.120 ;
        RECT 4.000 52.040 696.130 54.720 ;
        RECT 4.400 50.640 695.600 52.040 ;
        RECT 4.000 48.640 696.130 50.640 ;
        RECT 4.400 47.240 695.600 48.640 ;
        RECT 4.000 45.240 696.130 47.240 ;
        RECT 4.400 43.840 695.600 45.240 ;
        RECT 4.000 41.840 696.130 43.840 ;
        RECT 4.400 40.440 695.600 41.840 ;
        RECT 4.000 37.760 696.130 40.440 ;
        RECT 4.400 36.360 695.600 37.760 ;
        RECT 4.000 34.360 696.130 36.360 ;
        RECT 4.400 32.960 695.600 34.360 ;
        RECT 4.000 30.960 696.130 32.960 ;
        RECT 4.400 29.560 695.600 30.960 ;
        RECT 4.000 26.880 696.130 29.560 ;
        RECT 4.400 25.480 695.600 26.880 ;
        RECT 4.000 23.480 696.130 25.480 ;
        RECT 4.400 22.080 695.600 23.480 ;
        RECT 4.000 20.080 696.130 22.080 ;
        RECT 4.400 18.680 695.600 20.080 ;
        RECT 4.000 16.680 696.130 18.680 ;
        RECT 4.400 15.280 695.600 16.680 ;
        RECT 4.000 12.600 696.130 15.280 ;
        RECT 4.400 11.200 695.600 12.600 ;
        RECT 4.000 9.200 696.130 11.200 ;
        RECT 4.400 7.800 695.600 9.200 ;
        RECT 4.000 5.800 696.130 7.800 ;
        RECT 4.400 4.400 695.600 5.800 ;
        RECT 4.000 2.400 696.130 4.400 ;
        RECT 4.400 1.535 695.600 2.400 ;
      LAYER met4 ;
        RECT 16.855 688.800 681.425 697.505 ;
        RECT 16.855 10.640 20.640 688.800 ;
        RECT 23.040 10.640 97.440 688.800 ;
        RECT 99.840 10.640 681.425 688.800 ;
  END
END baked_disjoint_switch_box
END LIBRARY

