VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2860.860 BY 3400.460 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 70.990 2855.580 71.590 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 212.430 2855.580 213.030 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 353.870 2855.580 354.470 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 495.990 2855.580 496.590 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 637.430 2855.580 638.030 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 778.870 2855.580 779.470 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 920.990 2855.580 921.590 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1062.430 2855.580 1063.030 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1203.870 2855.580 1204.470 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1345.990 2855.580 1346.590 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 43.850 3396.230 44.130 3400.230 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 120.670 3396.230 120.950 3400.230 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 197.490 3396.230 197.770 3400.230 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 274.770 3396.230 275.050 3400.230 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 351.590 3396.230 351.870 3400.230 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 428.870 3396.230 429.150 3400.230 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 505.690 3396.230 505.970 3400.230 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 582.970 3396.230 583.250 3400.230 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 659.790 3396.230 660.070 3400.230 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 737.070 3396.230 737.350 3400.230 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 30.970 0.230 31.250 4.230 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.570 0.230 81.850 4.230 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 132.630 0.230 132.910 4.230 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 183.230 0.230 183.510 4.230 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 234.290 0.230 234.570 4.230 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 285.350 0.230 285.630 4.230 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 335.950 0.230 336.230 4.230 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 387.010 0.230 387.290 4.230 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 62.830 9.580 63.430 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 188.630 9.580 189.230 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 314.430 9.580 315.030 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 440.230 9.580 440.830 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 566.030 9.580 566.630 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 691.830 9.580 692.430 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 818.310 9.580 818.910 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 944.110 9.580 944.710 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1069.910 9.580 1070.510 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1195.710 9.580 1196.310 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2066.470 0.230 2066.750 4.230 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.530 0.230 2117.810 4.230 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2168.590 0.230 2168.870 4.230 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2219.190 0.230 2219.470 4.230 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.910 3396.230 1199.190 3400.230 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.190 3396.230 1276.470 3400.230 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1353.010 3396.230 1353.290 3400.230 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1447.990 9.580 1448.590 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1573.790 9.580 1574.390 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1430.290 3396.230 1430.570 3400.230 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2371.910 0.230 2372.190 4.230 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2422.970 0.230 2423.250 4.230 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1628.870 2855.580 1629.470 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1770.990 2855.580 1771.590 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2270.250 0.230 2270.530 4.230 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1507.110 3396.230 1507.390 3400.230 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1584.390 3396.230 1584.670 3400.230 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.210 3396.230 1661.490 3400.230 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1699.590 9.580 1700.190 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1912.430 2855.580 1913.030 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.490 3396.230 1738.770 3400.230 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1815.310 3396.230 1815.590 3400.230 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1892.590 3396.230 1892.870 3400.230 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1825.390 9.580 1825.990 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1969.410 3396.230 1969.690 3400.230 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.890 3396.230 814.170 3400.230 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2053.870 2855.580 2054.470 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1951.190 9.580 1951.790 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2320.850 0.230 2321.130 4.230 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.170 3396.230 891.450 3400.230 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 1321.510 9.580 1322.110 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.990 3396.230 968.270 3400.230 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.810 3396.230 1045.090 3400.230 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 1487.430 2855.580 1488.030 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.090 3396.230 1122.370 3400.230 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2195.990 2855.580 2196.590 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2337.430 2855.580 2338.030 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2329.270 9.580 2329.870 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2354.430 3396.230 2354.710 3400.230 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2620.990 2855.580 2621.590 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2431.710 3396.230 2431.990 3400.230 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2455.070 9.580 2455.670 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2508.530 3396.230 2508.810 3400.230 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2575.690 0.230 2575.970 4.230 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2626.290 0.230 2626.570 4.230 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2677.350 0.230 2677.630 4.230 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2762.430 2855.580 2763.030 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2076.990 9.580 2077.590 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2903.870 2855.580 2904.470 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2580.870 9.580 2581.470 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2706.670 9.580 2707.270 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2728.410 0.230 2728.690 4.230 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 3045.990 2855.580 3046.590 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2585.810 3396.230 2586.090 3400.230 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2779.010 0.230 2779.290 4.230 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2662.630 3396.230 2662.910 3400.230 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2739.910 3396.230 2740.190 3400.230 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2830.070 0.230 2830.350 4.230 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2046.230 3396.230 2046.510 3400.230 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2833.150 9.580 2833.750 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2816.730 3396.230 2817.010 3400.230 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.570 0.230 2473.850 4.230 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2203.470 9.580 2204.070 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2123.510 3396.230 2123.790 3400.230 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2200.330 3396.230 2200.610 3400.230 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2524.630 0.230 2524.910 4.230 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 2478.870 2855.580 2479.470 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2277.610 3396.230 2277.890 3400.230 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.070 0.230 438.350 4.230 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 946.830 0.230 947.110 4.230 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.890 0.230 998.170 4.230 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1048.490 0.230 1048.770 4.230 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1099.550 0.230 1099.830 4.230 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1150.610 0.230 1150.890 4.230 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.210 0.230 1201.490 4.230 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1252.270 0.230 1252.550 4.230 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.330 0.230 1303.610 4.230 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.930 0.230 1354.210 4.230 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1404.990 0.230 1405.270 4.230 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.670 0.230 488.950 4.230 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.050 0.230 1456.330 4.230 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1506.650 0.230 1506.930 4.230 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1557.710 0.230 1557.990 4.230 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1608.310 0.230 1608.590 4.230 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1659.370 0.230 1659.650 4.230 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1710.430 0.230 1710.710 4.230 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1761.030 0.230 1761.310 4.230 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1812.090 0.230 1812.370 4.230 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1863.150 0.230 1863.430 4.230 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1913.750 0.230 1914.030 4.230 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.730 0.230 540.010 4.230 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1964.810 0.230 1965.090 4.230 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2015.870 0.230 2016.150 4.230 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 590.790 0.230 591.070 4.230 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 641.390 0.230 641.670 4.230 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.450 0.230 692.730 4.230 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 743.510 0.230 743.790 4.230 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.110 0.230 794.390 4.230 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.170 0.230 845.450 4.230 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 895.770 0.230 896.050 4.230 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 2958.950 9.580 2959.550 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 3084.750 9.580 3085.350 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 3210.550 9.580 3211.150 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 3187.430 2855.580 3188.030 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.580 3336.350 9.580 3336.950 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2851.580 3328.870 2855.580 3329.470 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 4.600 4.610 2856.260 7.610 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.010 2860.860 3.010 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 11.100 11.025 2849.760 3389.435 ;
      LAYER met1 ;
        RECT 11.100 10.870 2849.760 3389.590 ;
      LAYER met2 ;
        RECT 19.930 3395.950 43.570 3396.230 ;
        RECT 44.410 3395.950 120.390 3396.230 ;
        RECT 121.230 3395.950 197.210 3396.230 ;
        RECT 198.050 3395.950 274.490 3396.230 ;
        RECT 275.330 3395.950 351.310 3396.230 ;
        RECT 352.150 3395.950 428.590 3396.230 ;
        RECT 429.430 3395.950 505.410 3396.230 ;
        RECT 506.250 3395.950 582.690 3396.230 ;
        RECT 583.530 3395.950 659.510 3396.230 ;
        RECT 660.350 3395.950 736.790 3396.230 ;
        RECT 737.630 3395.950 813.610 3396.230 ;
        RECT 814.450 3395.950 890.890 3396.230 ;
        RECT 891.730 3395.950 967.710 3396.230 ;
        RECT 968.550 3395.950 1044.530 3396.230 ;
        RECT 1045.370 3395.950 1121.810 3396.230 ;
        RECT 1122.650 3395.950 1198.630 3396.230 ;
        RECT 1199.470 3395.950 1275.910 3396.230 ;
        RECT 1276.750 3395.950 1352.730 3396.230 ;
        RECT 1353.570 3395.950 1430.010 3396.230 ;
        RECT 1430.850 3395.950 1506.830 3396.230 ;
        RECT 1507.670 3395.950 1584.110 3396.230 ;
        RECT 1584.950 3395.950 1660.930 3396.230 ;
        RECT 1661.770 3395.950 1738.210 3396.230 ;
        RECT 1739.050 3395.950 1815.030 3396.230 ;
        RECT 1815.870 3395.950 1892.310 3396.230 ;
        RECT 1893.150 3395.950 1969.130 3396.230 ;
        RECT 1969.970 3395.950 2045.950 3396.230 ;
        RECT 2046.790 3395.950 2123.230 3396.230 ;
        RECT 2124.070 3395.950 2200.050 3396.230 ;
        RECT 2200.890 3395.950 2277.330 3396.230 ;
        RECT 2278.170 3395.950 2354.150 3396.230 ;
        RECT 2354.990 3395.950 2431.430 3396.230 ;
        RECT 2432.270 3395.950 2508.250 3396.230 ;
        RECT 2509.090 3395.950 2585.530 3396.230 ;
        RECT 2586.370 3395.950 2662.350 3396.230 ;
        RECT 2663.190 3395.950 2739.630 3396.230 ;
        RECT 2740.470 3395.950 2816.450 3396.230 ;
        RECT 2817.290 3395.950 2844.160 3396.230 ;
        RECT 19.930 4.510 2844.160 3395.950 ;
        RECT 19.930 4.230 30.690 4.510 ;
        RECT 31.530 4.230 81.290 4.510 ;
        RECT 82.130 4.230 132.350 4.510 ;
        RECT 133.190 4.230 182.950 4.510 ;
        RECT 183.790 4.230 234.010 4.510 ;
        RECT 234.850 4.230 285.070 4.510 ;
        RECT 285.910 4.230 335.670 4.510 ;
        RECT 336.510 4.230 386.730 4.510 ;
        RECT 387.570 4.230 437.790 4.510 ;
        RECT 438.630 4.230 488.390 4.510 ;
        RECT 489.230 4.230 539.450 4.510 ;
        RECT 540.290 4.230 590.510 4.510 ;
        RECT 591.350 4.230 641.110 4.510 ;
        RECT 641.950 4.230 692.170 4.510 ;
        RECT 693.010 4.230 743.230 4.510 ;
        RECT 744.070 4.230 793.830 4.510 ;
        RECT 794.670 4.230 844.890 4.510 ;
        RECT 845.730 4.230 895.490 4.510 ;
        RECT 896.330 4.230 946.550 4.510 ;
        RECT 947.390 4.230 997.610 4.510 ;
        RECT 998.450 4.230 1048.210 4.510 ;
        RECT 1049.050 4.230 1099.270 4.510 ;
        RECT 1100.110 4.230 1150.330 4.510 ;
        RECT 1151.170 4.230 1200.930 4.510 ;
        RECT 1201.770 4.230 1251.990 4.510 ;
        RECT 1252.830 4.230 1303.050 4.510 ;
        RECT 1303.890 4.230 1353.650 4.510 ;
        RECT 1354.490 4.230 1404.710 4.510 ;
        RECT 1405.550 4.230 1455.770 4.510 ;
        RECT 1456.610 4.230 1506.370 4.510 ;
        RECT 1507.210 4.230 1557.430 4.510 ;
        RECT 1558.270 4.230 1608.030 4.510 ;
        RECT 1608.870 4.230 1659.090 4.510 ;
        RECT 1659.930 4.230 1710.150 4.510 ;
        RECT 1710.990 4.230 1760.750 4.510 ;
        RECT 1761.590 4.230 1811.810 4.510 ;
        RECT 1812.650 4.230 1862.870 4.510 ;
        RECT 1863.710 4.230 1913.470 4.510 ;
        RECT 1914.310 4.230 1964.530 4.510 ;
        RECT 1965.370 4.230 2015.590 4.510 ;
        RECT 2016.430 4.230 2066.190 4.510 ;
        RECT 2067.030 4.230 2117.250 4.510 ;
        RECT 2118.090 4.230 2168.310 4.510 ;
        RECT 2169.150 4.230 2218.910 4.510 ;
        RECT 2219.750 4.230 2269.970 4.510 ;
        RECT 2270.810 4.230 2320.570 4.510 ;
        RECT 2321.410 4.230 2371.630 4.510 ;
        RECT 2372.470 4.230 2422.690 4.510 ;
        RECT 2423.530 4.230 2473.290 4.510 ;
        RECT 2474.130 4.230 2524.350 4.510 ;
        RECT 2525.190 4.230 2575.410 4.510 ;
        RECT 2576.250 4.230 2626.010 4.510 ;
        RECT 2626.850 4.230 2677.070 4.510 ;
        RECT 2677.910 4.230 2728.130 4.510 ;
        RECT 2728.970 4.230 2778.730 4.510 ;
        RECT 2779.570 4.230 2829.790 4.510 ;
        RECT 2830.630 4.230 2844.160 4.510 ;
      LAYER met3 ;
        RECT 9.580 3337.350 2851.580 3389.515 ;
        RECT 9.980 3335.950 2851.580 3337.350 ;
        RECT 9.580 3329.870 2851.580 3335.950 ;
        RECT 9.580 3328.470 2851.180 3329.870 ;
        RECT 9.580 3211.550 2851.580 3328.470 ;
        RECT 9.980 3210.150 2851.580 3211.550 ;
        RECT 9.580 3188.430 2851.580 3210.150 ;
        RECT 9.580 3187.030 2851.180 3188.430 ;
        RECT 9.580 3085.750 2851.580 3187.030 ;
        RECT 9.980 3084.350 2851.580 3085.750 ;
        RECT 9.580 3046.990 2851.580 3084.350 ;
        RECT 9.580 3045.590 2851.180 3046.990 ;
        RECT 9.580 2959.950 2851.580 3045.590 ;
        RECT 9.980 2958.550 2851.580 2959.950 ;
        RECT 9.580 2904.870 2851.580 2958.550 ;
        RECT 9.580 2903.470 2851.180 2904.870 ;
        RECT 9.580 2834.150 2851.580 2903.470 ;
        RECT 9.980 2832.750 2851.580 2834.150 ;
        RECT 9.580 2763.430 2851.580 2832.750 ;
        RECT 9.580 2762.030 2851.180 2763.430 ;
        RECT 9.580 2707.670 2851.580 2762.030 ;
        RECT 9.980 2706.270 2851.580 2707.670 ;
        RECT 9.580 2621.990 2851.580 2706.270 ;
        RECT 9.580 2620.590 2851.180 2621.990 ;
        RECT 9.580 2581.870 2851.580 2620.590 ;
        RECT 9.980 2580.470 2851.580 2581.870 ;
        RECT 9.580 2479.870 2851.580 2580.470 ;
        RECT 9.580 2478.470 2851.180 2479.870 ;
        RECT 9.580 2456.070 2851.580 2478.470 ;
        RECT 9.980 2454.670 2851.580 2456.070 ;
        RECT 9.580 2338.430 2851.580 2454.670 ;
        RECT 9.580 2337.030 2851.180 2338.430 ;
        RECT 9.580 2330.270 2851.580 2337.030 ;
        RECT 9.980 2328.870 2851.580 2330.270 ;
        RECT 9.580 2204.470 2851.580 2328.870 ;
        RECT 9.980 2203.070 2851.580 2204.470 ;
        RECT 9.580 2196.990 2851.580 2203.070 ;
        RECT 9.580 2195.590 2851.180 2196.990 ;
        RECT 9.580 2077.990 2851.580 2195.590 ;
        RECT 9.980 2076.590 2851.580 2077.990 ;
        RECT 9.580 2054.870 2851.580 2076.590 ;
        RECT 9.580 2053.470 2851.180 2054.870 ;
        RECT 9.580 1952.190 2851.580 2053.470 ;
        RECT 9.980 1950.790 2851.580 1952.190 ;
        RECT 9.580 1913.430 2851.580 1950.790 ;
        RECT 9.580 1912.030 2851.180 1913.430 ;
        RECT 9.580 1826.390 2851.580 1912.030 ;
        RECT 9.980 1824.990 2851.580 1826.390 ;
        RECT 9.580 1771.990 2851.580 1824.990 ;
        RECT 9.580 1770.590 2851.180 1771.990 ;
        RECT 9.580 1700.590 2851.580 1770.590 ;
        RECT 9.980 1699.190 2851.580 1700.590 ;
        RECT 9.580 1629.870 2851.580 1699.190 ;
        RECT 9.580 1628.470 2851.180 1629.870 ;
        RECT 9.580 1574.790 2851.580 1628.470 ;
        RECT 9.980 1573.390 2851.580 1574.790 ;
        RECT 9.580 1488.430 2851.580 1573.390 ;
        RECT 9.580 1487.030 2851.180 1488.430 ;
        RECT 9.580 1448.990 2851.580 1487.030 ;
        RECT 9.980 1447.590 2851.580 1448.990 ;
        RECT 9.580 1346.990 2851.580 1447.590 ;
        RECT 9.580 1345.590 2851.180 1346.990 ;
        RECT 9.580 1322.510 2851.580 1345.590 ;
        RECT 9.980 1321.110 2851.580 1322.510 ;
        RECT 9.580 1204.870 2851.580 1321.110 ;
        RECT 9.580 1203.470 2851.180 1204.870 ;
        RECT 9.580 1196.710 2851.580 1203.470 ;
        RECT 9.980 1195.310 2851.580 1196.710 ;
        RECT 9.580 1070.910 2851.580 1195.310 ;
        RECT 9.980 1069.510 2851.580 1070.910 ;
        RECT 9.580 1063.430 2851.580 1069.510 ;
        RECT 9.580 1062.030 2851.180 1063.430 ;
        RECT 9.580 945.110 2851.580 1062.030 ;
        RECT 9.980 943.710 2851.580 945.110 ;
        RECT 9.580 921.990 2851.580 943.710 ;
        RECT 9.580 920.590 2851.180 921.990 ;
        RECT 9.580 819.310 2851.580 920.590 ;
        RECT 9.980 817.910 2851.580 819.310 ;
        RECT 9.580 779.870 2851.580 817.910 ;
        RECT 9.580 778.470 2851.180 779.870 ;
        RECT 9.580 692.830 2851.580 778.470 ;
        RECT 9.980 691.430 2851.580 692.830 ;
        RECT 9.580 638.430 2851.580 691.430 ;
        RECT 9.580 637.030 2851.180 638.430 ;
        RECT 9.580 567.030 2851.580 637.030 ;
        RECT 9.980 565.630 2851.580 567.030 ;
        RECT 9.580 496.990 2851.580 565.630 ;
        RECT 9.580 495.590 2851.180 496.990 ;
        RECT 9.580 441.230 2851.580 495.590 ;
        RECT 9.980 439.830 2851.580 441.230 ;
        RECT 9.580 354.870 2851.580 439.830 ;
        RECT 9.580 353.470 2851.180 354.870 ;
        RECT 9.580 315.430 2851.580 353.470 ;
        RECT 9.980 314.030 2851.580 315.430 ;
        RECT 9.580 213.430 2851.580 314.030 ;
        RECT 9.580 212.030 2851.180 213.430 ;
        RECT 9.580 189.630 2851.580 212.030 ;
        RECT 9.980 188.230 2851.580 189.630 ;
        RECT 9.580 71.990 2851.580 188.230 ;
        RECT 9.580 70.590 2851.180 71.990 ;
        RECT 9.580 63.830 2851.580 70.590 ;
        RECT 9.980 62.430 2851.580 63.830 ;
        RECT 9.580 10.945 2851.580 62.430 ;
      LAYER met4 ;
        RECT 0.000 0.010 2860.860 3400.450 ;
      LAYER met5 ;
        RECT 0.000 9.210 2860.860 3400.460 ;
        RECT 0.000 4.610 3.000 9.210 ;
        RECT 2857.860 4.610 2860.860 9.210 ;
  END
END fpga
END LIBRARY

