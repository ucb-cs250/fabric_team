magic
tech sky130A
magscale 1 2
timestamp 1623572100
<< locali >>
rect 9505 10999 9539 11101
rect 4537 9979 4571 10217
rect 121 3859 155 4097
rect 673 1819 707 4233
rect 765 2635 799 4165
rect 857 3655 891 9469
rect 6285 9367 6319 9469
rect 2697 7803 2731 8041
rect 2881 6103 2915 6409
rect 949 1411 983 5729
rect 2881 5559 2915 5865
rect 6469 5151 6503 5321
rect 6411 5117 6503 5151
rect 8493 5015 8527 5117
rect 12449 4811 12483 7361
rect 8585 3587 8619 3689
rect 4721 2839 4755 3145
rect 6285 2839 6319 3145
rect 7389 2839 7423 2941
<< viali >>
rect 6193 12937 6227 12971
rect 7757 12937 7791 12971
rect 7941 12937 7975 12971
rect 8401 12937 8435 12971
rect 8861 12937 8895 12971
rect 9873 12937 9907 12971
rect 11345 12937 11379 12971
rect 2973 12869 3007 12903
rect 6561 12869 6595 12903
rect 8585 12869 8619 12903
rect 10333 12869 10367 12903
rect 3341 12801 3375 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 11069 12801 11103 12835
rect 1961 12733 1995 12767
rect 2513 12733 2547 12767
rect 2789 12733 2823 12767
rect 3074 12733 3108 12767
rect 3525 12733 3559 12767
rect 4353 12733 4387 12767
rect 4629 12733 4663 12767
rect 4997 12733 5031 12767
rect 5549 12733 5583 12767
rect 5641 12733 5675 12767
rect 6101 12733 6135 12767
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 7205 12733 7239 12767
rect 8125 12733 8159 12767
rect 8585 12733 8619 12767
rect 8769 12733 8803 12767
rect 9045 12733 9079 12767
rect 9229 12733 9263 12767
rect 10057 12733 10091 12767
rect 10517 12733 10551 12767
rect 10885 12733 10919 12767
rect 11713 12733 11747 12767
rect 7665 12665 7699 12699
rect 8309 12665 8343 12699
rect 9781 12665 9815 12699
rect 11253 12665 11287 12699
rect 1869 12597 1903 12631
rect 2145 12597 2179 12631
rect 2421 12597 2455 12631
rect 2697 12597 2731 12631
rect 4169 12597 4203 12631
rect 4905 12597 4939 12631
rect 5365 12597 5399 12631
rect 9321 12597 9355 12631
rect 11529 12597 11563 12631
rect 5273 12393 5307 12427
rect 8493 12393 8527 12427
rect 9137 12393 9171 12427
rect 3709 12325 3743 12359
rect 4160 12325 4194 12359
rect 9965 12325 9999 12359
rect 10394 12325 10428 12359
rect 1676 12257 1710 12291
rect 2881 12257 2915 12291
rect 3525 12257 3559 12291
rect 5365 12257 5399 12291
rect 5632 12257 5666 12291
rect 6837 12257 6871 12291
rect 7093 12257 7127 12291
rect 8585 12257 8619 12291
rect 8769 12257 8803 12291
rect 9321 12257 9355 12291
rect 9879 12257 9913 12291
rect 10057 12257 10091 12291
rect 11621 12257 11655 12291
rect 1409 12189 1443 12223
rect 3893 12189 3927 12223
rect 9597 12189 9631 12223
rect 10156 12189 10190 12223
rect 6745 12121 6779 12155
rect 8309 12121 8343 12155
rect 2789 12053 2823 12087
rect 8217 12053 8251 12087
rect 9505 12053 9539 12087
rect 11529 12053 11563 12087
rect 4537 11849 4571 11883
rect 5089 11849 5123 11883
rect 6561 11849 6595 11883
rect 6653 11849 6687 11883
rect 7481 11849 7515 11883
rect 9137 11849 9171 11883
rect 9413 11849 9447 11883
rect 10241 11849 10275 11883
rect 11253 11849 11287 11883
rect 1685 11781 1719 11815
rect 2145 11713 2179 11747
rect 2329 11713 2363 11747
rect 2513 11713 2547 11747
rect 4997 11713 5031 11747
rect 5181 11713 5215 11747
rect 6745 11713 6779 11747
rect 10333 11713 10367 11747
rect 1409 11645 1443 11679
rect 4169 11645 4203 11679
rect 4445 11645 4479 11679
rect 4905 11645 4939 11679
rect 5273 11645 5307 11679
rect 5733 11645 5767 11679
rect 6009 11645 6043 11679
rect 6285 11645 6319 11679
rect 6469 11645 6503 11679
rect 6837 11645 6871 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 8024 11645 8058 11679
rect 9321 11645 9355 11679
rect 9689 11645 9723 11679
rect 9873 11645 9907 11679
rect 10058 11645 10092 11679
rect 10149 11645 10183 11679
rect 10425 11645 10459 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 11161 11645 11195 11679
rect 11437 11645 11471 11679
rect 2780 11577 2814 11611
rect 5365 11577 5399 11611
rect 6929 11577 6963 11611
rect 10517 11577 10551 11611
rect 1501 11509 1535 11543
rect 2053 11509 2087 11543
rect 3893 11509 3927 11543
rect 3985 11509 4019 11543
rect 5549 11509 5583 11543
rect 5825 11509 5859 11543
rect 6101 11509 6135 11543
rect 7205 11509 7239 11543
rect 10977 11509 11011 11543
rect 1685 11305 1719 11339
rect 2789 11305 2823 11339
rect 3065 11305 3099 11339
rect 5273 11305 5307 11339
rect 5457 11305 5491 11339
rect 7481 11305 7515 11339
rect 10149 11305 10183 11339
rect 11161 11305 11195 11339
rect 1869 11237 1903 11271
rect 4169 11237 4203 11271
rect 6368 11237 6402 11271
rect 7849 11237 7883 11271
rect 8493 11237 8527 11271
rect 8709 11237 8743 11271
rect 9965 11237 9999 11271
rect 1409 11169 1443 11203
rect 1777 11169 1811 11203
rect 2145 11169 2179 11203
rect 2329 11169 2363 11203
rect 2513 11169 2547 11203
rect 2881 11169 2915 11203
rect 3341 11169 3375 11203
rect 3525 11169 3559 11203
rect 3893 11169 3927 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 5089 11169 5123 11203
rect 5181 11169 5215 11203
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6101 11169 6135 11203
rect 8125 11169 8159 11203
rect 9137 11169 9171 11203
rect 9689 11169 9723 11203
rect 10589 11169 10623 11203
rect 10682 11169 10716 11203
rect 10798 11169 10832 11203
rect 10977 11169 11011 11203
rect 11075 11169 11109 11203
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 1685 11101 1719 11135
rect 2237 11101 2271 11135
rect 2789 11101 2823 11135
rect 3433 11101 3467 11135
rect 4169 11101 4203 11135
rect 9505 11101 9539 11135
rect 9772 11101 9806 11135
rect 9873 11101 9907 11135
rect 10149 11101 10183 11135
rect 3985 11033 4019 11067
rect 4261 11033 4295 11067
rect 8033 11033 8067 11067
rect 8217 11033 8251 11067
rect 9321 11033 9355 11067
rect 1501 10965 1535 10999
rect 2605 10965 2639 10999
rect 4537 10965 4571 10999
rect 4905 10965 4939 10999
rect 5917 10965 5951 10999
rect 8677 10965 8711 10999
rect 8861 10965 8895 10999
rect 9505 10965 9539 10999
rect 10333 10965 10367 10999
rect 11345 10965 11379 10999
rect 1409 10761 1443 10795
rect 5549 10761 5583 10795
rect 6101 10761 6135 10795
rect 6193 10761 6227 10795
rect 6561 10761 6595 10795
rect 8861 10761 8895 10795
rect 9505 10761 9539 10795
rect 11529 10761 11563 10795
rect 2605 10693 2639 10727
rect 6745 10693 6779 10727
rect 2053 10625 2087 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 5825 10625 5859 10659
rect 6285 10625 6319 10659
rect 7297 10625 7331 10659
rect 9781 10625 9815 10659
rect 9965 10625 9999 10659
rect 1777 10557 1811 10591
rect 1869 10557 1903 10591
rect 2329 10557 2363 10591
rect 2513 10557 2547 10591
rect 2789 10557 2823 10591
rect 3065 10557 3099 10591
rect 3617 10557 3651 10591
rect 4252 10557 4286 10591
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 5917 10557 5951 10591
rect 6009 10557 6043 10591
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 6929 10557 6963 10591
rect 7021 10557 7055 10591
rect 7564 10557 7598 10591
rect 9045 10557 9079 10591
rect 9321 10557 9355 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 10149 10557 10183 10591
rect 10405 10557 10439 10591
rect 11897 10557 11931 10591
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 3157 10421 3191 10455
rect 3525 10421 3559 10455
rect 5365 10421 5399 10455
rect 7205 10421 7239 10455
rect 8677 10421 8711 10455
rect 9229 10421 9263 10455
rect 11713 10421 11747 10455
rect 4537 10217 4571 10251
rect 4905 10217 4939 10251
rect 5181 10217 5215 10251
rect 9505 10217 9539 10251
rect 9965 10217 9999 10251
rect 10425 10217 10459 10251
rect 1685 10149 1719 10183
rect 2022 10149 2056 10183
rect 3617 10149 3651 10183
rect 1409 10081 1443 10115
rect 1501 10081 1535 10115
rect 3433 10081 3467 10115
rect 3525 10081 3559 10115
rect 4077 10081 4111 10115
rect 4353 10081 4387 10115
rect 1685 10013 1719 10047
rect 1777 10013 1811 10047
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 5816 10081 5850 10115
rect 7113 10081 7147 10115
rect 7481 10081 7515 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 8033 10081 8067 10115
rect 8493 10081 8527 10115
rect 8769 10081 8803 10115
rect 8953 10081 8987 10115
rect 9137 10081 9171 10115
rect 9781 10081 9815 10115
rect 10241 10081 10275 10115
rect 10425 10081 10459 10115
rect 10876 10081 10910 10115
rect 5549 10013 5583 10047
rect 7389 10013 7423 10047
rect 7849 10013 7883 10047
rect 10609 10013 10643 10047
rect 3157 9945 3191 9979
rect 4537 9945 4571 9979
rect 4721 9945 4755 9979
rect 3249 9877 3283 9911
rect 3893 9877 3927 9911
rect 4169 9877 4203 9911
rect 6929 9877 6963 9911
rect 7205 9877 7239 9911
rect 7297 9877 7331 9911
rect 8769 9877 8803 9911
rect 9505 9877 9539 9911
rect 9689 9877 9723 9911
rect 11989 9877 12023 9911
rect 2881 9673 2915 9707
rect 5733 9673 5767 9707
rect 6929 9673 6963 9707
rect 8769 9673 8803 9707
rect 10609 9673 10643 9707
rect 10793 9673 10827 9707
rect 1961 9605 1995 9639
rect 3341 9605 3375 9639
rect 4261 9605 4295 9639
rect 8493 9605 8527 9639
rect 2513 9537 2547 9571
rect 3985 9537 4019 9571
rect 4445 9537 4479 9571
rect 4813 9537 4847 9571
rect 5365 9537 5399 9571
rect 7113 9537 7147 9571
rect 11897 9537 11931 9571
rect 857 9469 891 9503
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 3065 9469 3099 9503
rect 3801 9469 3835 9503
rect 4169 9469 4203 9503
rect 4721 9469 4755 9503
rect 4905 9469 4939 9503
rect 5181 9469 5215 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 5825 9469 5859 9503
rect 6009 9469 6043 9503
rect 6193 9469 6227 9503
rect 6285 9469 6319 9503
rect 6469 9469 6503 9503
rect 6837 9469 6871 9503
rect 7380 9469 7414 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 9689 9469 9723 9503
rect 10149 9469 10183 9503
rect 10885 9469 10919 9503
rect 11529 9469 11563 9503
rect 673 4233 707 4267
rect 121 4097 155 4131
rect 121 3825 155 3859
rect 765 4165 799 4199
rect 3709 9401 3743 9435
rect 6101 9401 6135 9435
rect 9965 9401 9999 9435
rect 10333 9401 10367 9435
rect 10425 9401 10459 9435
rect 10641 9401 10675 9435
rect 1409 9333 1443 9367
rect 1685 9333 1719 9367
rect 2421 9333 2455 9367
rect 3157 9333 3191 9367
rect 4445 9333 4479 9367
rect 4997 9333 5031 9367
rect 6285 9333 6319 9367
rect 2789 9129 2823 9163
rect 5273 9129 5307 9163
rect 5825 9129 5859 9163
rect 6561 9129 6595 9163
rect 6653 9129 6687 9163
rect 8401 9129 8435 9163
rect 9137 9129 9171 9163
rect 9597 9129 9631 9163
rect 3525 9061 3559 9095
rect 3709 9061 3743 9095
rect 4160 9061 4194 9095
rect 9965 9061 9999 9095
rect 10333 9061 10367 9095
rect 10425 9061 10459 9095
rect 10641 9061 10675 9095
rect 10977 9061 11011 9095
rect 1409 8993 1443 9027
rect 1676 8993 1710 9027
rect 3065 8993 3099 9027
rect 3341 8993 3375 9027
rect 5733 8993 5767 9027
rect 7021 8993 7055 9027
rect 7205 8993 7239 9027
rect 7297 8993 7331 9027
rect 7573 8993 7607 9027
rect 8033 8993 8067 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 8677 8993 8711 9027
rect 9505 8993 9539 9027
rect 10149 8993 10183 9027
rect 10885 8993 10919 9027
rect 11069 8993 11103 9027
rect 3893 8925 3927 8959
rect 6009 8925 6043 8959
rect 6745 8925 6779 8959
rect 8861 8925 8895 8959
rect 9689 8925 9723 8959
rect 2881 8857 2915 8891
rect 5365 8857 5399 8891
rect 3157 8789 3191 8823
rect 6193 8789 6227 8823
rect 7113 8789 7147 8823
rect 10609 8789 10643 8823
rect 10793 8789 10827 8823
rect 11345 8789 11379 8823
rect 11621 8789 11655 8823
rect 11897 8789 11931 8823
rect 1409 8585 1443 8619
rect 1869 8585 1903 8619
rect 2053 8585 2087 8619
rect 4261 8585 4295 8619
rect 8401 8585 8435 8619
rect 8953 8585 8987 8619
rect 9413 8585 9447 8619
rect 11253 8585 11287 8619
rect 1777 8517 1811 8551
rect 6101 8517 6135 8551
rect 1961 8449 1995 8483
rect 2421 8449 2455 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5641 8449 5675 8483
rect 6929 8449 6963 8483
rect 10149 8449 10183 8483
rect 1593 8381 1627 8415
rect 1685 8381 1719 8415
rect 2237 8381 2271 8415
rect 2329 8381 2363 8415
rect 2513 8381 2547 8415
rect 2614 8381 2648 8415
rect 2881 8381 2915 8415
rect 4905 8381 4939 8415
rect 5365 8381 5399 8415
rect 5457 8381 5491 8415
rect 6653 8381 6687 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 8493 8381 8527 8415
rect 8861 8381 8895 8415
rect 9229 8381 9263 8415
rect 9781 8381 9815 8415
rect 9873 8381 9907 8415
rect 11897 8381 11931 8415
rect 3126 8313 3160 8347
rect 5917 8313 5951 8347
rect 6929 8313 6963 8347
rect 7266 8313 7300 8347
rect 4537 8245 4571 8279
rect 5641 8245 5675 8279
rect 2513 8041 2547 8075
rect 2697 8041 2731 8075
rect 3065 8041 3099 8075
rect 4537 8041 4571 8075
rect 6377 8041 6411 8075
rect 8401 8041 8435 8075
rect 2053 7973 2087 8007
rect 1961 7905 1995 7939
rect 2421 7905 2455 7939
rect 2237 7837 2271 7871
rect 3985 7973 4019 8007
rect 4988 7973 5022 8007
rect 10600 7973 10634 8007
rect 2789 7905 2823 7939
rect 2881 7905 2915 7939
rect 3249 7905 3283 7939
rect 3433 7905 3467 7939
rect 3525 7905 3559 7939
rect 4445 7905 4479 7939
rect 4721 7905 4755 7939
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 7021 7905 7055 7939
rect 7941 7905 7975 7939
rect 9137 7905 9171 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 6653 7837 6687 7871
rect 7205 7837 7239 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10333 7837 10367 7871
rect 1593 7769 1627 7803
rect 2697 7769 2731 7803
rect 4169 7769 4203 7803
rect 9229 7769 9263 7803
rect 6101 7701 6135 7735
rect 7113 7701 7147 7735
rect 7665 7701 7699 7735
rect 8033 7701 8067 7735
rect 9321 7701 9355 7735
rect 9965 7701 9999 7735
rect 10241 7701 10275 7735
rect 11713 7701 11747 7735
rect 11989 7701 12023 7735
rect 2697 7497 2731 7531
rect 3985 7497 4019 7531
rect 5181 7497 5215 7531
rect 6193 7497 6227 7531
rect 8401 7497 8435 7531
rect 10057 7497 10091 7531
rect 10425 7497 10459 7531
rect 3065 7429 3099 7463
rect 3525 7429 3559 7463
rect 10333 7429 10367 7463
rect 3709 7361 3743 7395
rect 5365 7361 5399 7395
rect 5825 7361 5859 7395
rect 8217 7361 8251 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 11345 7361 11379 7395
rect 12449 7361 12483 7395
rect 1501 7293 1535 7327
rect 1777 7293 1811 7327
rect 2237 7293 2271 7327
rect 2513 7293 2547 7327
rect 2605 7293 2639 7327
rect 3249 7293 3283 7327
rect 3433 7293 3467 7327
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 4813 7293 4847 7327
rect 5089 7293 5123 7327
rect 5457 7293 5491 7327
rect 5733 7293 5767 7327
rect 5917 7293 5951 7327
rect 8309 7293 8343 7327
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 8944 7293 8978 7327
rect 10241 7293 10275 7327
rect 10609 7293 10643 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 11897 7293 11931 7327
rect 3893 7225 3927 7259
rect 6101 7225 6135 7259
rect 6469 7225 6503 7259
rect 10701 7225 10735 7259
rect 2053 7157 2087 7191
rect 2329 7157 2363 7191
rect 3709 7157 3743 7191
rect 5365 7157 5399 7191
rect 2881 6953 2915 6987
rect 6745 6953 6779 6987
rect 9781 6953 9815 6987
rect 9873 6953 9907 6987
rect 10609 6953 10643 6987
rect 10701 6953 10735 6987
rect 3249 6885 3283 6919
rect 7104 6885 7138 6919
rect 8493 6885 8527 6919
rect 8677 6885 8711 6919
rect 1676 6817 1710 6851
rect 4149 6817 4183 6851
rect 5365 6817 5399 6851
rect 5632 6817 5666 6851
rect 6837 6817 6871 6851
rect 8769 6817 8803 6851
rect 8861 6817 8895 6851
rect 9137 6817 9171 6851
rect 11069 6817 11103 6851
rect 1409 6749 1443 6783
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 3893 6749 3927 6783
rect 9965 6749 9999 6783
rect 10793 6749 10827 6783
rect 11529 6749 11563 6783
rect 2789 6681 2823 6715
rect 8217 6681 8251 6715
rect 9229 6681 9263 6715
rect 9413 6681 9447 6715
rect 5273 6613 5307 6647
rect 10241 6613 10275 6647
rect 11161 6613 11195 6647
rect 11805 6613 11839 6647
rect 1501 6409 1535 6443
rect 1593 6409 1627 6443
rect 2697 6409 2731 6443
rect 2881 6409 2915 6443
rect 3709 6409 3743 6443
rect 3985 6409 4019 6443
rect 5917 6409 5951 6443
rect 6561 6409 6595 6443
rect 7113 6409 7147 6443
rect 1685 6273 1719 6307
rect 2421 6273 2455 6307
rect 1409 6205 1443 6239
rect 2237 6205 2271 6239
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 2145 6137 2179 6171
rect 8309 6341 8343 6375
rect 5549 6273 5583 6307
rect 6745 6273 6779 6307
rect 7757 6273 7791 6307
rect 8493 6273 8527 6307
rect 10149 6273 10183 6307
rect 3065 6205 3099 6239
rect 3341 6205 3375 6239
rect 3617 6205 3651 6239
rect 3893 6205 3927 6239
rect 4077 6205 4111 6239
rect 4169 6205 4203 6239
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 5825 6205 5859 6239
rect 6285 6205 6319 6239
rect 6469 6205 6503 6239
rect 6837 6205 6871 6239
rect 7481 6205 7515 6239
rect 7941 6205 7975 6239
rect 8217 6205 8251 6239
rect 8401 6205 8435 6239
rect 11713 6205 11747 6239
rect 11897 6205 11931 6239
rect 5365 6137 5399 6171
rect 5457 6137 5491 6171
rect 6929 6137 6963 6171
rect 8760 6137 8794 6171
rect 10416 6137 10450 6171
rect 1777 6069 1811 6103
rect 2881 6069 2915 6103
rect 4997 6069 5031 6103
rect 6745 6069 6779 6103
rect 7573 6069 7607 6103
rect 8125 6069 8159 6103
rect 9873 6069 9907 6103
rect 11529 6069 11563 6103
rect 11805 6069 11839 6103
rect 1777 5865 1811 5899
rect 2421 5865 2455 5899
rect 2881 5865 2915 5899
rect 3893 5865 3927 5899
rect 5181 5865 5215 5899
rect 5733 5865 5767 5899
rect 7941 5865 7975 5899
rect 9781 5865 9815 5899
rect 10701 5865 10735 5899
rect 857 3621 891 3655
rect 949 5729 983 5763
rect 1593 5729 1627 5763
rect 1685 5729 1719 5763
rect 765 2601 799 2635
rect 673 1785 707 1819
rect 2513 5661 2547 5695
rect 2605 5661 2639 5695
rect 1409 5593 1443 5627
rect 4261 5797 4295 5831
rect 6193 5797 6227 5831
rect 6806 5797 6840 5831
rect 8953 5797 8987 5831
rect 11069 5797 11103 5831
rect 2973 5729 3007 5763
rect 3525 5729 3559 5763
rect 4721 5729 4755 5763
rect 5089 5729 5123 5763
rect 5365 5729 5399 5763
rect 6101 5729 6135 5763
rect 6561 5729 6595 5763
rect 8401 5729 8435 5763
rect 8585 5729 8619 5763
rect 8677 5729 8711 5763
rect 9145 5729 9179 5763
rect 9597 5729 9631 5763
rect 9781 5729 9815 5763
rect 9873 5729 9907 5763
rect 10425 5729 10459 5763
rect 10885 5729 10919 5763
rect 11897 5729 11931 5763
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 4353 5661 4387 5695
rect 4537 5661 4571 5695
rect 6285 5661 6319 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 10149 5661 10183 5695
rect 10701 5661 10735 5695
rect 9965 5593 9999 5627
rect 10517 5593 10551 5627
rect 11345 5593 11379 5627
rect 2053 5525 2087 5559
rect 2881 5525 2915 5559
rect 3157 5525 3191 5559
rect 8309 5525 8343 5559
rect 8769 5525 8803 5559
rect 10057 5525 10091 5559
rect 11621 5525 11655 5559
rect 2789 5321 2823 5355
rect 2973 5321 3007 5355
rect 4537 5321 4571 5355
rect 6285 5321 6319 5355
rect 6469 5321 6503 5355
rect 8677 5321 8711 5355
rect 9597 5321 9631 5355
rect 11529 5321 11563 5355
rect 5273 5253 5307 5287
rect 7113 5185 7147 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 9137 5185 9171 5219
rect 9229 5185 9263 5219
rect 10149 5185 10183 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 3157 5117 3191 5151
rect 3413 5117 3447 5151
rect 4629 5117 4663 5151
rect 5641 5117 5675 5151
rect 5825 5117 5859 5151
rect 6377 5117 6411 5151
rect 6929 5117 6963 5151
rect 7389 5117 7423 5151
rect 7481 5117 7515 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 8401 5117 8435 5151
rect 8493 5117 8527 5151
rect 9045 5117 9079 5151
rect 9505 5117 9539 5151
rect 10405 5117 10439 5151
rect 11805 5117 11839 5151
rect 1676 5049 1710 5083
rect 5089 5049 5123 5083
rect 5457 5049 5491 5083
rect 7021 5049 7055 5083
rect 9873 5049 9907 5083
rect 11989 5049 12023 5083
rect 4813 4981 4847 5015
rect 5917 4981 5951 5015
rect 6561 4981 6595 5015
rect 7665 4981 7699 5015
rect 8125 4981 8159 5015
rect 8493 4981 8527 5015
rect 9965 4981 9999 5015
rect 2421 4777 2455 4811
rect 4353 4777 4387 4811
rect 8677 4777 8711 4811
rect 9137 4777 9171 4811
rect 9505 4777 9539 4811
rect 10425 4777 10459 4811
rect 10793 4777 10827 4811
rect 12449 4777 12483 4811
rect 2605 4709 2639 4743
rect 4905 4709 4939 4743
rect 6745 4709 6779 4743
rect 7564 4709 7598 4743
rect 9597 4709 9631 4743
rect 10885 4709 10919 4743
rect 11437 4709 11471 4743
rect 1501 4641 1535 4675
rect 1869 4641 1903 4675
rect 2145 4641 2179 4675
rect 2513 4641 2547 4675
rect 2789 4641 2823 4675
rect 2973 4641 3007 4675
rect 3249 4641 3283 4675
rect 3525 4641 3559 4675
rect 3985 4641 4019 4675
rect 4169 4641 4203 4675
rect 4261 4641 4295 4675
rect 4445 4641 4479 4675
rect 4721 4641 4755 4675
rect 5448 4641 5482 4675
rect 7021 4641 7055 4675
rect 8769 4641 8803 4675
rect 10057 4641 10091 4675
rect 11805 4641 11839 4675
rect 2421 4573 2455 4607
rect 2881 4573 2915 4607
rect 5181 4573 5215 4607
rect 7297 4573 7331 4607
rect 9689 4573 9723 4607
rect 10977 4573 11011 4607
rect 2237 4505 2271 4539
rect 7113 4505 7147 4539
rect 11989 4505 12023 4539
rect 1593 4437 1627 4471
rect 4077 4437 4111 4471
rect 4997 4437 5031 4471
rect 6561 4437 6595 4471
rect 6837 4437 6871 4471
rect 8861 4437 8895 4471
rect 10149 4437 10183 4471
rect 11529 4437 11563 4471
rect 2237 4233 2271 4267
rect 3433 4233 3467 4267
rect 5457 4233 5491 4267
rect 6009 4233 6043 4267
rect 6561 4233 6595 4267
rect 7573 4233 7607 4267
rect 8401 4233 8435 4267
rect 9045 4165 9079 4199
rect 2789 4097 2823 4131
rect 3617 4097 3651 4131
rect 6756 4097 6790 4131
rect 6929 4097 6963 4131
rect 7389 4097 7423 4131
rect 9229 4097 9263 4131
rect 11161 4097 11195 4131
rect 1685 4029 1719 4063
rect 2605 4029 2639 4063
rect 2697 4029 2731 4063
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 3341 4029 3375 4063
rect 3709 4029 3743 4063
rect 5733 4029 5767 4063
rect 6285 4029 6319 4063
rect 6469 4029 6503 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7481 4029 7515 4063
rect 7941 4029 7975 4063
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 8953 4029 8987 4063
rect 9321 4029 9355 4063
rect 10977 4029 11011 4063
rect 11805 4029 11839 4063
rect 1501 3961 1535 3995
rect 1869 3961 1903 3995
rect 3617 3961 3651 3995
rect 3954 3961 3988 3995
rect 8309 3961 8343 3995
rect 9229 3961 9263 3995
rect 9566 3961 9600 3995
rect 11345 3961 11379 3995
rect 11529 3961 11563 3995
rect 1961 3893 1995 3927
rect 3157 3893 3191 3927
rect 5089 3893 5123 3927
rect 6745 3893 6779 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 10701 3893 10735 3927
rect 11897 3893 11931 3927
rect 2789 3689 2823 3723
rect 3985 3689 4019 3723
rect 7389 3689 7423 3723
rect 7757 3689 7791 3723
rect 8493 3689 8527 3723
rect 8585 3689 8619 3723
rect 9689 3689 9723 3723
rect 10425 3689 10459 3723
rect 3157 3621 3191 3655
rect 5273 3621 5307 3655
rect 6745 3621 6779 3655
rect 9229 3621 9263 3655
rect 9965 3621 9999 3655
rect 10701 3621 10735 3655
rect 10885 3621 10919 3655
rect 11437 3621 11471 3655
rect 11805 3621 11839 3655
rect 1409 3553 1443 3587
rect 1676 3553 1710 3587
rect 2881 3553 2915 3587
rect 3249 3553 3283 3587
rect 3525 3553 3559 3587
rect 3893 3553 3927 3587
rect 4169 3553 4203 3587
rect 4353 3553 4387 3587
rect 4813 3553 4847 3587
rect 5181 3553 5215 3587
rect 5457 3553 5491 3587
rect 5641 3553 5675 3587
rect 5917 3553 5951 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 8217 3553 8251 3587
rect 8585 3553 8619 3587
rect 8769 3553 8803 3587
rect 8953 3553 8987 3587
rect 9597 3553 9631 3587
rect 10333 3553 10367 3587
rect 11069 3553 11103 3587
rect 3157 3485 3191 3519
rect 4905 3485 4939 3519
rect 5089 3485 5123 3519
rect 5549 3485 5583 3519
rect 6561 3485 6595 3519
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 8493 3485 8527 3519
rect 9413 3485 9447 3519
rect 11253 3485 11287 3519
rect 3617 3417 3651 3451
rect 6469 3417 6503 3451
rect 7297 3417 7331 3451
rect 10149 3417 10183 3451
rect 11989 3417 12023 3451
rect 2973 3349 3007 3383
rect 3341 3349 3375 3383
rect 4261 3349 4295 3383
rect 4721 3349 4755 3383
rect 4997 3349 5031 3383
rect 6193 3349 6227 3383
rect 6377 3349 6411 3383
rect 8309 3349 8343 3383
rect 11529 3349 11563 3383
rect 2697 3145 2731 3179
rect 3893 3145 3927 3179
rect 4721 3145 4755 3179
rect 6193 3145 6227 3179
rect 6285 3145 6319 3179
rect 6469 3145 6503 3179
rect 8861 3145 8895 3179
rect 11897 3145 11931 3179
rect 3617 3077 3651 3111
rect 2053 3009 2087 3043
rect 3341 3009 3375 3043
rect 3801 3009 3835 3043
rect 4537 3009 4571 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 2145 2941 2179 2975
rect 3065 2941 3099 2975
rect 3525 2941 3559 2975
rect 3157 2873 3191 2907
rect 4261 2873 4295 2907
rect 4813 3009 4847 3043
rect 5080 2941 5114 2975
rect 3801 2805 3835 2839
rect 4353 2805 4387 2839
rect 4721 2805 4755 2839
rect 10609 3077 10643 3111
rect 6929 3009 6963 3043
rect 7021 3009 7055 3043
rect 9321 3009 9355 3043
rect 7389 2941 7423 2975
rect 7481 2941 7515 2975
rect 10057 2941 10091 2975
rect 10793 2941 10827 2975
rect 10977 2941 11011 2975
rect 11805 2941 11839 2975
rect 7748 2873 7782 2907
rect 9137 2873 9171 2907
rect 9505 2873 9539 2907
rect 10241 2873 10275 2907
rect 10425 2873 10459 2907
rect 11161 2873 11195 2907
rect 6285 2805 6319 2839
rect 6837 2805 6871 2839
rect 7389 2805 7423 2839
rect 9597 2805 9631 2839
rect 11253 2805 11287 2839
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 5365 2601 5399 2635
rect 5733 2601 5767 2635
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 8953 2601 8987 2635
rect 10057 2601 10091 2635
rect 2789 2533 2823 2567
rect 4160 2533 4194 2567
rect 6828 2533 6862 2567
rect 8401 2533 8435 2567
rect 9321 2533 9355 2567
rect 9689 2533 9723 2567
rect 11069 2533 11103 2567
rect 11437 2533 11471 2567
rect 1593 2465 1627 2499
rect 1961 2465 1995 2499
rect 2145 2465 2179 2499
rect 2697 2465 2731 2499
rect 3893 2465 3927 2499
rect 5825 2465 5859 2499
rect 6193 2465 6227 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 8493 2465 8527 2499
rect 8861 2465 8895 2499
rect 9965 2465 9999 2499
rect 10149 2465 10183 2499
rect 10333 2465 10367 2499
rect 10701 2465 10735 2499
rect 3433 2397 3467 2431
rect 3525 2397 3559 2431
rect 5917 2397 5951 2431
rect 8585 2397 8619 2431
rect 5273 2329 5307 2363
rect 8033 2329 8067 2363
rect 9873 2329 9907 2363
rect 10517 2329 10551 2363
rect 9413 2261 9447 2295
rect 10793 2261 10827 2295
rect 11161 2261 11195 2295
rect 11529 2261 11563 2295
rect 949 1377 983 1411
<< metal1 >>
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 10042 13512 10048 13524
rect 2740 13484 10048 13512
rect 2740 13472 2746 13484
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 658 13404 664 13456
rect 716 13444 722 13456
rect 9030 13444 9036 13456
rect 716 13416 9036 13444
rect 716 13404 722 13416
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 474 13336 480 13388
rect 532 13376 538 13388
rect 8110 13376 8116 13388
rect 532 13348 8116 13376
rect 532 13336 538 13348
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 7926 13240 7932 13252
rect 2372 13212 7932 13240
rect 2372 13200 2378 13212
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 382 13132 388 13184
rect 440 13172 446 13184
rect 6178 13172 6184 13184
rect 440 13144 6184 13172
rect 440 13132 446 13144
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 1104 13082 12328 13104
rect 1104 13030 2852 13082
rect 2904 13030 2916 13082
rect 2968 13030 2980 13082
rect 3032 13030 3044 13082
rect 3096 13030 6594 13082
rect 6646 13030 6658 13082
rect 6710 13030 6722 13082
rect 6774 13030 6786 13082
rect 6838 13030 10335 13082
rect 10387 13030 10399 13082
rect 10451 13030 10463 13082
rect 10515 13030 10527 13082
rect 10579 13030 12328 13082
rect 1104 13008 12328 13030
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5224 12940 6193 12968
rect 5224 12928 5230 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 6972 12940 7757 12968
rect 6972 12928 6978 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7745 12931 7803 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8849 12971 8907 12977
rect 8849 12968 8861 12971
rect 8496 12940 8861 12968
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 3418 12900 3424 12912
rect 3007 12872 3424 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 3418 12860 3424 12872
rect 3476 12860 3482 12912
rect 4338 12860 4344 12912
rect 4396 12900 4402 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 4396 12872 6561 12900
rect 4396 12860 4402 12872
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 6549 12863 6607 12869
rect 290 12792 296 12844
rect 348 12832 354 12844
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 348 12804 2820 12832
rect 348 12792 354 12804
rect 1854 12724 1860 12776
rect 1912 12764 1918 12776
rect 1949 12767 2007 12773
rect 1949 12764 1961 12767
rect 1912 12736 1961 12764
rect 1912 12724 1918 12736
rect 1949 12733 1961 12736
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 2792 12773 2820 12804
rect 2976 12804 3341 12832
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 2464 12736 2513 12764
rect 2464 12724 2470 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 2976 12764 3004 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4580 12804 4721 12832
rect 4580 12792 4586 12804
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 5258 12832 5264 12844
rect 4939 12804 5264 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 8496 12832 8524 12940
rect 8849 12937 8861 12940
rect 8895 12937 8907 12971
rect 8849 12931 8907 12937
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9732 12940 9873 12968
rect 9732 12928 9738 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11296 12940 11345 12968
rect 11296 12928 11302 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 10321 12903 10379 12909
rect 8628 12872 8673 12900
rect 8628 12860 8634 12872
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 11146 12900 11152 12912
rect 10367 12872 11152 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 8846 12832 8852 12844
rect 5500 12804 8524 12832
rect 8588 12804 8852 12832
rect 5500 12792 5506 12804
rect 2823 12736 3004 12764
rect 3062 12767 3120 12773
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3062 12733 3074 12767
rect 3108 12764 3120 12767
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3108 12736 3525 12764
rect 3108 12733 3120 12736
rect 3062 12727 3120 12733
rect 3513 12733 3525 12736
rect 3559 12733 3571 12767
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 3513 12727 3571 12733
rect 4172 12736 4353 12764
rect 934 12656 940 12708
rect 992 12696 998 12708
rect 3068 12696 3096 12727
rect 992 12668 3096 12696
rect 992 12656 998 12668
rect 4172 12640 4200 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4614 12764 4620 12776
rect 4575 12736 4620 12764
rect 4341 12727 4399 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5166 12764 5172 12776
rect 5031 12736 5172 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5534 12764 5540 12776
rect 5495 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5684 12736 6101 12764
rect 5684 12724 5690 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 6733 12767 6791 12773
rect 6733 12764 6745 12767
rect 6236 12736 6745 12764
rect 6236 12724 6242 12736
rect 6733 12733 6745 12736
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 6825 12727 6883 12733
rect 6840 12696 6868 12727
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8588 12773 8616 12804
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 11057 12835 11115 12841
rect 9180 12804 10916 12832
rect 9180 12792 9186 12804
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 8754 12764 8760 12776
rect 8715 12736 8760 12764
rect 8573 12727 8631 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9214 12764 9220 12776
rect 9175 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10888 12773 10916 12804
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 12618 12832 12624 12844
rect 11103 12804 12624 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 10873 12727 10931 12733
rect 10980 12736 11713 12764
rect 7098 12696 7104 12708
rect 6840 12668 7104 12696
rect 7098 12656 7104 12668
rect 7156 12696 7162 12708
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 7156 12668 7665 12696
rect 7156 12656 7162 12668
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 8297 12699 8355 12705
rect 8297 12696 8309 12699
rect 8260 12668 8309 12696
rect 8260 12656 8266 12668
rect 8297 12665 8309 12668
rect 8343 12665 8355 12699
rect 9769 12699 9827 12705
rect 9769 12696 9781 12699
rect 8297 12659 8355 12665
rect 8404 12668 9781 12696
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 2096 12600 2145 12628
rect 2096 12588 2102 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2406 12628 2412 12640
rect 2367 12600 2412 12628
rect 2133 12591 2191 12597
rect 2406 12588 2412 12600
rect 2464 12588 2470 12640
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2648 12600 2697 12628
rect 2648 12588 2654 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 2685 12591 2743 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4304 12600 4905 12628
rect 4304 12588 4310 12600
rect 4893 12597 4905 12600
rect 4939 12597 4951 12631
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 4893 12591 4951 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8404 12628 8432 12668
rect 9769 12665 9781 12668
rect 9815 12665 9827 12699
rect 9769 12659 9827 12665
rect 10520 12696 10548 12727
rect 10980 12696 11008 12736
rect 11701 12733 11713 12736
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 10520 12668 11008 12696
rect 11241 12699 11299 12705
rect 9306 12628 9312 12640
rect 8076 12600 8432 12628
rect 9267 12600 9312 12628
rect 8076 12588 8082 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 10520 12628 10548 12668
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 11606 12696 11612 12708
rect 11287 12668 11612 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11514 12628 11520 12640
rect 9548 12600 10548 12628
rect 11475 12600 11520 12628
rect 9548 12588 9554 12600
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 1104 12538 12328 12560
rect 1104 12486 4723 12538
rect 4775 12486 4787 12538
rect 4839 12486 4851 12538
rect 4903 12486 4915 12538
rect 4967 12486 8464 12538
rect 8516 12486 8528 12538
rect 8580 12486 8592 12538
rect 8644 12486 8656 12538
rect 8708 12486 12328 12538
rect 1104 12464 12328 12486
rect 2406 12384 2412 12436
rect 2464 12424 2470 12436
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 2464 12396 2912 12424
rect 2464 12384 2470 12396
rect 1670 12297 1676 12300
rect 1664 12251 1676 12297
rect 1728 12288 1734 12300
rect 2884 12297 2912 12396
rect 5184 12396 5273 12424
rect 5184 12368 5212 12396
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 6362 12424 6368 12436
rect 5684 12396 6368 12424
rect 5684 12384 5690 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 8481 12427 8539 12433
rect 6472 12396 7411 12424
rect 3694 12356 3700 12368
rect 3655 12328 3700 12356
rect 3694 12316 3700 12328
rect 3752 12316 3758 12368
rect 4148 12359 4206 12365
rect 4148 12325 4160 12359
rect 4194 12356 4206 12359
rect 4246 12356 4252 12368
rect 4194 12328 4252 12356
rect 4194 12325 4206 12328
rect 4148 12319 4206 12325
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 5166 12356 5172 12368
rect 4448 12328 5172 12356
rect 4448 12300 4476 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 6472 12356 6500 12396
rect 7282 12356 7288 12368
rect 5368 12328 6500 12356
rect 6840 12328 7288 12356
rect 2869 12291 2927 12297
rect 1728 12260 1764 12288
rect 1670 12248 1676 12251
rect 1728 12248 1734 12260
rect 2869 12257 2881 12291
rect 2915 12257 2927 12291
rect 2869 12251 2927 12257
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12288 3571 12291
rect 4430 12288 4436 12300
rect 3559 12260 4436 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5368 12297 5396 12328
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5620 12291 5678 12297
rect 5620 12257 5632 12291
rect 5666 12288 5678 12291
rect 5902 12288 5908 12300
rect 5666 12260 5908 12288
rect 5666 12257 5678 12260
rect 5620 12251 5678 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 1412 12084 1440 12183
rect 1762 12084 1768 12096
rect 1412 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2777 12087 2835 12093
rect 2777 12084 2789 12087
rect 2188 12056 2789 12084
rect 2188 12044 2194 12056
rect 2777 12053 2789 12056
rect 2823 12053 2835 12087
rect 2777 12047 2835 12053
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 3896 12084 3924 12183
rect 5368 12152 5396 12251
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6840 12297 6868 12328
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 7383 12356 7411 12396
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 8754 12424 8760 12436
rect 8527 12396 8760 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8904 12396 9137 12424
rect 8904 12384 8910 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 11606 12424 11612 12436
rect 9640 12396 11612 12424
rect 9640 12384 9646 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 9766 12356 9772 12368
rect 7383 12328 9772 12356
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9953 12359 10011 12365
rect 9953 12325 9965 12359
rect 9999 12356 10011 12359
rect 10382 12359 10440 12365
rect 10382 12356 10394 12359
rect 9999 12328 10394 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 10382 12325 10394 12328
rect 10428 12325 10440 12359
rect 10382 12319 10440 12325
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7081 12291 7139 12297
rect 7081 12288 7093 12291
rect 6972 12260 7093 12288
rect 6972 12248 6978 12260
rect 7081 12257 7093 12260
rect 7127 12257 7139 12291
rect 7081 12251 7139 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 8938 12288 8944 12300
rect 8803 12260 8944 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 8588 12220 8616 12251
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9306 12288 9312 12300
rect 9267 12260 9312 12288
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9858 12248 9864 12300
rect 9916 12297 9922 12300
rect 9916 12288 9925 12297
rect 9916 12260 9961 12288
rect 9916 12251 9925 12260
rect 9916 12248 9922 12251
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 11606 12288 11612 12300
rect 10100 12260 10145 12288
rect 11567 12260 11612 12288
rect 10100 12248 10106 12260
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 9398 12220 9404 12232
rect 8588 12192 9404 12220
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 9950 12220 9956 12232
rect 9631 12192 9956 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10144 12223 10202 12229
rect 10144 12189 10156 12223
rect 10190 12189 10202 12223
rect 10144 12183 10202 12189
rect 4816 12124 5396 12152
rect 4816 12084 4844 12124
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 6733 12155 6791 12161
rect 6733 12152 6745 12155
rect 6420 12124 6745 12152
rect 6420 12112 6426 12124
rect 6733 12121 6745 12124
rect 6779 12121 6791 12155
rect 6733 12115 6791 12121
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8297 12155 8355 12161
rect 8297 12152 8309 12155
rect 8168 12124 8309 12152
rect 8168 12112 8174 12124
rect 8297 12121 8309 12124
rect 8343 12121 8355 12155
rect 8297 12115 8355 12121
rect 3844 12056 4844 12084
rect 3844 12044 3850 12056
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 7006 12084 7012 12096
rect 5040 12056 7012 12084
rect 5040 12044 5046 12056
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 8202 12084 8208 12096
rect 7248 12056 8208 12084
rect 7248 12044 7254 12056
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9493 12087 9551 12093
rect 9493 12084 9505 12087
rect 8996 12056 9505 12084
rect 8996 12044 9002 12056
rect 9493 12053 9505 12056
rect 9539 12053 9551 12087
rect 9493 12047 9551 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10152 12084 10180 12183
rect 9824 12056 10180 12084
rect 9824 12044 9830 12056
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 10836 12056 11529 12084
rect 10836 12044 10842 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11517 12047 11575 12053
rect 1104 11994 12328 12016
rect 1104 11942 2852 11994
rect 2904 11942 2916 11994
rect 2968 11942 2980 11994
rect 3032 11942 3044 11994
rect 3096 11942 6594 11994
rect 6646 11942 6658 11994
rect 6710 11942 6722 11994
rect 6774 11942 6786 11994
rect 6838 11942 10335 11994
rect 10387 11942 10399 11994
rect 10451 11942 10463 11994
rect 10515 11942 10527 11994
rect 10579 11942 12328 11994
rect 1104 11920 12328 11942
rect 1118 11840 1124 11892
rect 1176 11880 1182 11892
rect 4525 11883 4583 11889
rect 1176 11852 4200 11880
rect 1176 11840 1182 11852
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11781 1731 11815
rect 1673 11775 1731 11781
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1688 11676 1716 11775
rect 1762 11772 1768 11824
rect 1820 11812 1826 11824
rect 1820 11784 2544 11812
rect 1820 11772 1826 11784
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2516 11753 2544 11784
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 1443 11648 1716 11676
rect 2332 11676 2360 11707
rect 2406 11676 2412 11688
rect 2332 11648 2412 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 2516 11676 2544 11707
rect 3786 11676 3792 11688
rect 2516 11648 3792 11676
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 4172 11685 4200 11852
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 4614 11880 4620 11892
rect 4571 11852 4620 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5074 11880 5080 11892
rect 5035 11852 5080 11880
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5810 11880 5816 11892
rect 5224 11852 5816 11880
rect 5224 11840 5230 11852
rect 5810 11840 5816 11852
rect 5868 11880 5874 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 5868 11852 6561 11880
rect 5868 11840 5874 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 6914 11880 6920 11892
rect 6687 11852 6920 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7469 11883 7527 11889
rect 7469 11880 7481 11883
rect 7064 11852 7481 11880
rect 7064 11840 7070 11852
rect 7469 11849 7481 11852
rect 7515 11849 7527 11883
rect 7469 11843 7527 11849
rect 9125 11883 9183 11889
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 9214 11880 9220 11892
rect 9171 11852 9220 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 9916 11852 10241 11880
rect 9916 11840 9922 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 11238 11880 11244 11892
rect 11199 11852 11244 11880
rect 10229 11843 10287 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 5350 11812 5356 11824
rect 4255 11784 5356 11812
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 2774 11617 2780 11620
rect 2768 11571 2780 11617
rect 2832 11608 2838 11620
rect 4255 11608 4283 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 7742 11812 7748 11824
rect 6104 11784 7748 11812
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4580 11716 4997 11744
rect 4580 11704 4586 11716
rect 4985 11713 4997 11716
rect 5031 11744 5043 11747
rect 5074 11744 5080 11756
rect 5031 11716 5080 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5534 11744 5540 11756
rect 5215 11716 5540 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 4430 11676 4436 11688
rect 4391 11648 4436 11676
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11676 5319 11679
rect 5718 11676 5724 11688
rect 5307 11648 5488 11676
rect 5679 11648 5724 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 2832 11580 2868 11608
rect 3252 11580 4283 11608
rect 4908 11608 4936 11639
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 4908 11580 5365 11608
rect 2774 11568 2780 11571
rect 2832 11568 2838 11580
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 1946 11540 1952 11552
rect 1535 11512 1952 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 3252 11540 3280 11580
rect 5353 11577 5365 11580
rect 5399 11577 5411 11611
rect 5460 11608 5488 11648
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 5994 11676 6000 11688
rect 5955 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 5626 11608 5632 11620
rect 5460 11580 5632 11608
rect 5353 11571 5411 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6104 11608 6132 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 9784 11784 10640 11812
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6420 11716 6745 11744
rect 6420 11704 6426 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 9784 11744 9812 11784
rect 10321 11747 10379 11753
rect 6733 11707 6791 11713
rect 9692 11716 9812 11744
rect 9876 11716 10272 11744
rect 9692 11688 9720 11716
rect 9876 11688 9904 11716
rect 6270 11676 6276 11688
rect 6231 11648 6276 11676
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 6457 11679 6515 11685
rect 6457 11645 6469 11679
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7190 11676 7196 11688
rect 6871 11648 7196 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 5736 11580 6132 11608
rect 6472 11608 6500 11639
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7650 11676 7656 11688
rect 7611 11648 7656 11676
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8012 11679 8070 11685
rect 8012 11645 8024 11679
rect 8058 11676 8070 11679
rect 8294 11676 8300 11688
rect 8058 11648 8300 11676
rect 8058 11645 8070 11648
rect 8012 11639 8070 11645
rect 6917 11611 6975 11617
rect 6917 11608 6929 11611
rect 6472 11580 6929 11608
rect 2087 11512 3280 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 3326 11500 3332 11552
rect 3384 11540 3390 11552
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3384 11512 3893 11540
rect 3384 11500 3390 11512
rect 3881 11509 3893 11512
rect 3927 11509 3939 11543
rect 3881 11503 3939 11509
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5537 11543 5595 11549
rect 4028 11512 4073 11540
rect 4028 11500 4034 11512
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 5736 11540 5764 11580
rect 6917 11577 6929 11580
rect 6963 11577 6975 11611
rect 6917 11571 6975 11577
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 7760 11608 7788 11639
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9272 11648 9321 11676
rect 9272 11636 9278 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9674 11676 9680 11688
rect 9587 11648 9680 11676
rect 9309 11639 9367 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9858 11676 9864 11688
rect 9771 11648 9864 11676
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10046 11679 10104 11685
rect 10046 11676 10058 11679
rect 10008 11648 10058 11676
rect 10008 11636 10014 11648
rect 10046 11645 10058 11648
rect 10092 11645 10104 11679
rect 10046 11639 10104 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11645 10195 11679
rect 10244 11676 10272 11716
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10502 11744 10508 11756
rect 10367 11716 10508 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10612 11744 10640 11784
rect 10778 11744 10784 11756
rect 10612 11716 10784 11744
rect 10410 11676 10416 11688
rect 10244 11648 10416 11676
rect 10137 11639 10195 11645
rect 9766 11608 9772 11620
rect 7340 11580 9772 11608
rect 7340 11568 7346 11580
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 9876 11580 9996 11608
rect 5583 11512 5764 11540
rect 5813 11543 5871 11549
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 5902 11540 5908 11552
rect 5859 11512 5908 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6086 11540 6092 11552
rect 6047 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 7193 11543 7251 11549
rect 7193 11509 7205 11543
rect 7239 11540 7251 11543
rect 7558 11540 7564 11552
rect 7239 11512 7564 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9876 11540 9904 11580
rect 8996 11512 9904 11540
rect 9968 11540 9996 11580
rect 10152 11540 10180 11639
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10612 11685 10640 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11645 10747 11679
rect 11146 11676 11152 11688
rect 11107 11648 11152 11676
rect 10689 11639 10747 11645
rect 10226 11568 10232 11620
rect 10284 11608 10290 11620
rect 10505 11611 10563 11617
rect 10505 11608 10517 11611
rect 10284 11580 10517 11608
rect 10284 11568 10290 11580
rect 10505 11577 10517 11580
rect 10551 11577 10563 11611
rect 10505 11571 10563 11577
rect 9968 11512 10180 11540
rect 8996 11500 9002 11512
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10704 11540 10732 11639
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 11514 11676 11520 11688
rect 11471 11648 11520 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 10962 11540 10968 11552
rect 10376 11512 10732 11540
rect 10923 11512 10968 11540
rect 10376 11500 10382 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 1104 11450 12328 11472
rect 1104 11398 4723 11450
rect 4775 11398 4787 11450
rect 4839 11398 4851 11450
rect 4903 11398 4915 11450
rect 4967 11398 8464 11450
rect 8516 11398 8528 11450
rect 8580 11398 8592 11450
rect 8644 11398 8656 11450
rect 8708 11398 12328 11450
rect 1104 11376 12328 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2280 11308 2636 11336
rect 2280 11296 2286 11308
rect 1857 11271 1915 11277
rect 1857 11268 1869 11271
rect 1412 11240 1869 11268
rect 1412 11209 1440 11240
rect 1857 11237 1869 11240
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 2608 11268 2636 11308
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3053 11339 3111 11345
rect 2832 11308 2877 11336
rect 2832 11296 2838 11308
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 5074 11336 5080 11348
rect 3099 11308 5080 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 5626 11336 5632 11348
rect 5491 11308 5632 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 7098 11336 7104 11348
rect 5828 11308 7104 11336
rect 4157 11271 4215 11277
rect 2004 11240 2544 11268
rect 2608 11240 2774 11268
rect 2004 11228 2010 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1397 11163 1455 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2130 11200 2136 11212
rect 2091 11172 2136 11200
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2516 11209 2544 11240
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11169 2375 11203
rect 2317 11163 2375 11169
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11169 2559 11203
rect 2746 11200 2774 11240
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 4246 11268 4252 11280
rect 4203 11240 4252 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2746 11172 2881 11200
rect 2501 11163 2559 11169
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 3326 11200 3332 11212
rect 3287 11172 3332 11200
rect 2869 11163 2927 11169
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1719 11104 2237 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2332 11064 2360 11163
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11169 3571 11203
rect 3513 11163 3571 11169
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 3421 11135 3479 11141
rect 3421 11132 3433 11135
rect 2823 11104 3433 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 3421 11101 3433 11104
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 2498 11064 2504 11076
rect 2332 11036 2504 11064
rect 2498 11024 2504 11036
rect 2556 11064 2562 11076
rect 3528 11064 3556 11163
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3660 11172 3893 11200
rect 3660 11160 3666 11172
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 4120 11172 4283 11200
rect 4120 11160 4126 11172
rect 4154 11132 4160 11144
rect 4115 11104 4160 11132
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4255 11132 4283 11172
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4396 11172 4445 11200
rect 4396 11160 4402 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4580 11172 4721 11200
rect 4580 11160 4586 11172
rect 4709 11169 4721 11172
rect 4755 11169 4767 11203
rect 5074 11200 5080 11212
rect 5035 11172 5080 11200
rect 4709 11163 4767 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5442 11200 5448 11212
rect 5399 11172 5448 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5184 11132 5212 11163
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5828 11209 5856 11308
rect 7098 11296 7104 11308
rect 7156 11336 7162 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7156 11308 7481 11336
rect 7156 11296 7162 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 10100 11308 10149 11336
rect 10100 11296 10106 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 10594 11296 10600 11348
rect 10652 11296 10658 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10704 11308 11161 11336
rect 6356 11271 6414 11277
rect 6356 11237 6368 11271
rect 6402 11268 6414 11271
rect 6546 11268 6552 11280
rect 6402 11240 6552 11268
rect 6402 11237 6414 11240
rect 6356 11231 6414 11237
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 7837 11271 7895 11277
rect 7837 11237 7849 11271
rect 7883 11268 7895 11271
rect 8294 11268 8300 11280
rect 7883 11240 8300 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 8478 11268 8484 11280
rect 8439 11240 8484 11268
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8697 11271 8755 11277
rect 8697 11237 8709 11271
rect 8743 11268 8755 11271
rect 8938 11268 8944 11280
rect 8743 11240 8944 11268
rect 8743 11237 8755 11240
rect 8697 11231 8755 11237
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9232 11240 9803 11268
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 7282 11200 7288 11212
rect 6135 11172 7288 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 8110 11200 8116 11212
rect 8071 11172 8116 11200
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 9088 11172 9137 11200
rect 9088 11160 9094 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 5994 11132 6000 11144
rect 4255 11104 5212 11132
rect 5736 11104 6000 11132
rect 2556 11036 3556 11064
rect 3973 11067 4031 11073
rect 2556 11024 2562 11036
rect 3973 11033 3985 11067
rect 4019 11033 4031 11067
rect 3973 11027 4031 11033
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 5626 11064 5632 11076
rect 4295 11036 5632 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10996 1550 11008
rect 2593 10999 2651 11005
rect 2593 10996 2605 10999
rect 1544 10968 2605 10996
rect 1544 10956 1550 10968
rect 2593 10965 2605 10968
rect 2639 10996 2651 10999
rect 3878 10996 3884 11008
rect 2639 10968 3884 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 3878 10956 3884 10968
rect 3936 10996 3942 11008
rect 3988 10996 4016 11027
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 5736 11008 5764 11104
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 7926 11064 7932 11076
rect 5868 11036 6132 11064
rect 5868 11024 5874 11036
rect 3936 10968 4016 10996
rect 4525 10999 4583 11005
rect 3936 10956 3942 10968
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 4798 10996 4804 11008
rect 4571 10968 4804 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 4948 10968 4993 10996
rect 4948 10956 4954 10968
rect 5718 10956 5724 11008
rect 5776 10956 5782 11008
rect 5905 10999 5963 11005
rect 5905 10965 5917 10999
rect 5951 10996 5963 10999
rect 5994 10996 6000 11008
rect 5951 10968 6000 10996
rect 5951 10965 5963 10968
rect 5905 10959 5963 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6104 10996 6132 11036
rect 7024 11036 7932 11064
rect 7024 10996 7052 11036
rect 7926 11024 7932 11036
rect 7984 11064 7990 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 7984 11036 8033 11064
rect 7984 11024 7990 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 9232 11064 9260 11240
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9775 11200 9803 11240
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10008 11240 10053 11268
rect 10008 11228 10014 11240
rect 10410 11200 10416 11212
rect 9775 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10612 11209 10640 11296
rect 10704 11209 10732 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 10928 11240 11008 11268
rect 10928 11228 10934 11240
rect 10980 11209 11008 11240
rect 10577 11203 10640 11209
rect 10577 11169 10589 11203
rect 10623 11172 10640 11203
rect 10670 11203 10732 11209
rect 10623 11169 10635 11172
rect 10577 11163 10635 11169
rect 10670 11169 10682 11203
rect 10716 11172 10732 11203
rect 10786 11203 10844 11209
rect 10716 11169 10728 11172
rect 10670 11163 10728 11169
rect 10786 11169 10798 11203
rect 10832 11169 10844 11203
rect 10786 11163 10844 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11063 11203 11121 11209
rect 11063 11169 11075 11203
rect 11109 11169 11121 11203
rect 11238 11200 11244 11212
rect 11199 11172 11244 11200
rect 11063 11163 11121 11169
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9760 11135 9818 11141
rect 9760 11132 9772 11135
rect 9539 11104 9772 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9760 11101 9772 11104
rect 9806 11101 9818 11135
rect 9760 11095 9818 11101
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 9861 11095 9919 11101
rect 8251 11036 9260 11064
rect 9309 11067 9367 11073
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8680 11005 8708 11036
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9876 11064 9904 11095
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10428 11132 10456 11160
rect 10796 11132 10824 11163
rect 10428 11104 10824 11132
rect 9355 11036 10436 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9784 11008 9812 11036
rect 6104 10968 7052 10996
rect 8665 10999 8723 11005
rect 8665 10965 8677 10999
rect 8711 10965 8723 10999
rect 8846 10996 8852 11008
rect 8807 10968 8852 10996
rect 8665 10959 8723 10965
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 9493 10999 9551 11005
rect 9493 10996 9505 10999
rect 9272 10968 9505 10996
rect 9272 10956 9278 10968
rect 9493 10965 9505 10968
rect 9539 10965 9551 10999
rect 9493 10959 9551 10965
rect 9766 10956 9772 11008
rect 9824 10956 9830 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 10284 10968 10333 10996
rect 10284 10956 10290 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10408 10996 10436 11036
rect 11072 10996 11100 11163
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11514 11200 11520 11212
rect 11475 11172 11520 11200
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 11330 10996 11336 11008
rect 10408 10968 11100 10996
rect 11291 10968 11336 10996
rect 10321 10959 10379 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 1104 10906 12328 10928
rect 1104 10854 2852 10906
rect 2904 10854 2916 10906
rect 2968 10854 2980 10906
rect 3032 10854 3044 10906
rect 3096 10854 6594 10906
rect 6646 10854 6658 10906
rect 6710 10854 6722 10906
rect 6774 10854 6786 10906
rect 6838 10854 10335 10906
rect 10387 10854 10399 10906
rect 10451 10854 10463 10906
rect 10515 10854 10527 10906
rect 10579 10854 12328 10906
rect 1104 10832 12328 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 1762 10792 1768 10804
rect 1443 10764 1768 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 4614 10792 4620 10804
rect 1872 10764 4620 10792
rect 1872 10656 1900 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6089 10795 6147 10801
rect 6089 10792 6101 10795
rect 5868 10764 6101 10792
rect 5868 10752 5874 10764
rect 6089 10761 6101 10764
rect 6135 10761 6147 10795
rect 6089 10755 6147 10761
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6236 10764 6281 10792
rect 6236 10752 6242 10764
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6420 10764 6561 10792
rect 6420 10752 6426 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 6840 10764 8248 10792
rect 6840 10736 6868 10764
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 2774 10724 2780 10736
rect 2639 10696 2780 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 5316 10696 6745 10724
rect 5316 10684 5322 10696
rect 6733 10693 6745 10696
rect 6779 10693 6791 10727
rect 6733 10687 6791 10693
rect 6822 10684 6828 10736
rect 6880 10684 6886 10736
rect 8220 10724 8248 10764
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8536 10764 8861 10792
rect 8536 10752 8542 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 10870 10792 10876 10804
rect 9539 10764 10876 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11296 10764 11529 10792
rect 11296 10752 11302 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 9674 10724 9680 10736
rect 8220 10696 9680 10724
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 9858 10684 9864 10736
rect 9916 10684 9922 10736
rect 1780 10628 1900 10656
rect 2041 10659 2099 10665
rect 1780 10597 1808 10628
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2130 10656 2136 10668
rect 2087 10628 2136 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2130 10616 2136 10628
rect 2188 10656 2194 10668
rect 2406 10656 2412 10668
rect 2188 10628 2412 10656
rect 2188 10616 2194 10628
rect 2406 10616 2412 10628
rect 2464 10656 2470 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 2464 10628 3709 10656
rect 2464 10616 2470 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3844 10628 3985 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5813 10659 5871 10665
rect 5408 10628 5764 10656
rect 5408 10616 5414 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2317 10591 2375 10597
rect 2317 10588 2329 10591
rect 1903 10560 2329 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2317 10557 2329 10560
rect 2363 10557 2375 10591
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2317 10551 2375 10557
rect 106 10480 112 10532
rect 164 10520 170 10532
rect 2222 10520 2228 10532
rect 164 10492 2228 10520
rect 164 10480 170 10492
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 2332 10520 2360 10551
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 2866 10588 2872 10600
rect 2823 10560 2872 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3234 10588 3240 10600
rect 3099 10560 3240 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 4246 10597 4252 10600
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 3384 10560 3617 10588
rect 3384 10548 3390 10560
rect 3605 10557 3617 10560
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 4240 10551 4252 10597
rect 4304 10588 4310 10600
rect 4304 10560 4340 10588
rect 4246 10548 4252 10551
rect 4304 10548 4310 10560
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 4764 10560 5457 10588
rect 4764 10548 4770 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5736 10597 5764 10628
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5859 10628 6285 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 6273 10619 6331 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 9766 10656 9772 10668
rect 9048 10628 9772 10656
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5592 10560 5641 10588
rect 5592 10548 5598 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 2958 10520 2964 10532
rect 2332 10492 2964 10520
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 3694 10480 3700 10532
rect 3752 10520 3758 10532
rect 3752 10492 4108 10520
rect 3752 10480 3758 10492
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2866 10452 2872 10464
rect 2827 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3970 10452 3976 10464
rect 3559 10424 3976 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4080 10452 4108 10492
rect 4430 10480 4436 10532
rect 4488 10520 4494 10532
rect 5644 10520 5672 10551
rect 5920 10520 5948 10551
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6457 10591 6515 10597
rect 6052 10560 6097 10588
rect 6052 10548 6058 10560
rect 6457 10557 6469 10591
rect 6503 10588 6515 10591
rect 6546 10588 6552 10600
rect 6503 10560 6552 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10557 6699 10591
rect 6914 10588 6920 10600
rect 6875 10560 6920 10588
rect 6641 10551 6699 10557
rect 6656 10520 6684 10551
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7552 10591 7610 10597
rect 7552 10557 7564 10591
rect 7598 10588 7610 10591
rect 8846 10588 8852 10600
rect 7598 10560 8852 10588
rect 7598 10557 7610 10560
rect 7552 10551 7610 10557
rect 7024 10520 7052 10551
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9048 10597 9076 10628
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 9876 10656 9904 10684
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9876 10628 9965 10656
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 9272 10560 9321 10588
rect 9272 10548 9278 10560
rect 9309 10557 9321 10560
rect 9355 10588 9367 10591
rect 9674 10588 9680 10600
rect 9355 10560 9680 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9784 10560 9873 10588
rect 8294 10520 8300 10532
rect 4488 10492 5488 10520
rect 5644 10492 6960 10520
rect 7024 10492 8300 10520
rect 4488 10480 4494 10492
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 4080 10424 5365 10452
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5460 10452 5488 10492
rect 6822 10452 6828 10464
rect 5460 10424 6828 10452
rect 5353 10415 5411 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6932 10452 6960 10492
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 9784 10464 9812 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 10100 10560 10149 10588
rect 10100 10548 10106 10560
rect 10137 10557 10149 10560
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10393 10591 10451 10597
rect 10393 10588 10405 10591
rect 10284 10560 10405 10588
rect 10284 10548 10290 10560
rect 10393 10557 10405 10560
rect 10439 10557 10451 10591
rect 10393 10551 10451 10557
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11204 10560 11897 10588
rect 11204 10548 11210 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6932 10424 7205 10452
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7193 10415 7251 10421
rect 8665 10455 8723 10461
rect 8665 10421 8677 10455
rect 8711 10452 8723 10455
rect 9030 10452 9036 10464
rect 8711 10424 9036 10452
rect 8711 10421 8723 10424
rect 8665 10415 8723 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9217 10455 9275 10461
rect 9217 10421 9229 10455
rect 9263 10452 9275 10455
rect 9766 10452 9772 10464
rect 9263 10424 9772 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 9766 10412 9772 10424
rect 9824 10452 9830 10464
rect 10134 10452 10140 10464
rect 9824 10424 10140 10452
rect 9824 10412 9830 10424
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 10284 10424 11713 10452
rect 10284 10412 10290 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 1104 10362 12328 10384
rect 1104 10310 4723 10362
rect 4775 10310 4787 10362
rect 4839 10310 4851 10362
rect 4903 10310 4915 10362
rect 4967 10310 8464 10362
rect 8516 10310 8528 10362
rect 8580 10310 8592 10362
rect 8644 10310 8656 10362
rect 8708 10310 12328 10362
rect 1104 10288 12328 10310
rect 1854 10208 1860 10260
rect 1912 10248 1918 10260
rect 2590 10248 2596 10260
rect 1912 10220 2596 10248
rect 1912 10208 1918 10220
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 2740 10220 4108 10248
rect 2740 10208 2746 10220
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 2010 10183 2068 10189
rect 2010 10180 2022 10183
rect 1719 10152 2022 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 2010 10149 2022 10152
rect 2056 10149 2068 10183
rect 2010 10143 2068 10149
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 3200 10152 3556 10180
rect 3200 10140 3206 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 2406 10112 2412 10124
rect 1544 10084 1589 10112
rect 1688 10084 2412 10112
rect 1544 10072 1550 10084
rect 1688 10053 1716 10084
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 3234 10112 3240 10124
rect 2924 10084 3240 10112
rect 2924 10072 2930 10084
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 3528 10121 3556 10152
rect 3602 10140 3608 10192
rect 3660 10180 3666 10192
rect 3660 10152 3705 10180
rect 3660 10140 3666 10152
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 3384 10084 3433 10112
rect 3384 10072 3390 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4080 10121 4108 10220
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4212 10220 4537 10248
rect 4212 10208 4218 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4525 10211 4583 10217
rect 4724 10220 4905 10248
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 4724 10180 4752 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 7374 10248 7380 10260
rect 5215 10220 7380 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 8846 10248 8852 10260
rect 7484 10220 8852 10248
rect 5534 10180 5540 10192
rect 4488 10152 4752 10180
rect 4816 10152 5540 10180
rect 4488 10140 4494 10152
rect 4065 10115 4123 10121
rect 3752 10084 4016 10112
rect 3752 10072 3758 10084
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 1820 10016 1865 10044
rect 1820 10004 1826 10016
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3145 9979 3203 9985
rect 3145 9976 3157 9979
rect 3016 9948 3157 9976
rect 3016 9936 3022 9948
rect 3145 9945 3157 9948
rect 3191 9945 3203 9979
rect 3988 9976 4016 10084
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4341 10115 4399 10121
rect 4341 10112 4353 10115
rect 4212 10084 4353 10112
rect 4212 10072 4218 10084
rect 4341 10081 4353 10084
rect 4387 10081 4399 10115
rect 4614 10112 4620 10124
rect 4341 10075 4399 10081
rect 4448 10084 4620 10112
rect 4448 9976 4476 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4816 10121 4844 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5994 10180 6000 10192
rect 5736 10152 6000 10180
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 5077 10115 5135 10121
rect 5077 10112 5089 10115
rect 4948 10084 5089 10112
rect 4948 10072 4954 10084
rect 5077 10081 5089 10084
rect 5123 10081 5135 10115
rect 5077 10075 5135 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5736 10112 5764 10152
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 5399 10084 5764 10112
rect 5804 10115 5862 10121
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5804 10081 5816 10115
rect 5850 10112 5862 10115
rect 6178 10112 6184 10124
rect 5850 10084 6184 10112
rect 5850 10081 5862 10084
rect 5804 10075 5862 10081
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 7484 10121 7512 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9674 10248 9680 10260
rect 9539 10220 9680 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9674 10208 9680 10220
rect 9732 10248 9738 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9732 10220 9965 10248
rect 9732 10208 9738 10220
rect 9953 10217 9965 10220
rect 9999 10248 10011 10251
rect 10413 10251 10471 10257
rect 9999 10220 10272 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 8386 10180 8392 10192
rect 7760 10152 8392 10180
rect 7760 10121 7788 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 9858 10180 9864 10192
rect 8772 10152 9168 10180
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 7064 10084 7113 10112
rect 7064 10072 7070 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8202 10112 8208 10124
rect 8067 10084 8208 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7423 10016 7849 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 3988 9948 4476 9976
rect 4525 9979 4583 9985
rect 3145 9939 3203 9945
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 4709 9979 4767 9985
rect 4709 9976 4721 9979
rect 4571 9948 4721 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 4709 9945 4721 9948
rect 4755 9945 4767 9979
rect 4709 9939 4767 9945
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5552 9976 5580 10007
rect 7944 9976 7972 10075
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8662 10112 8668 10124
rect 8527 10084 8668 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 8772 10121 8800 10152
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10081 8815 10115
rect 8938 10112 8944 10124
rect 8899 10084 8944 10112
rect 8757 10075 8815 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9140 10121 9168 10152
rect 9508 10152 9864 10180
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9398 10112 9404 10124
rect 9171 10084 9404 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9214 9976 9220 9988
rect 5040 9948 5580 9976
rect 6472 9948 7972 9976
rect 8036 9948 9220 9976
rect 5040 9936 5046 9948
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3602 9908 3608 9920
rect 3283 9880 3608 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 4062 9908 4068 9920
rect 3927 9880 4068 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9908 4215 9911
rect 4430 9908 4436 9920
rect 4203 9880 4436 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6472 9908 6500 9948
rect 6914 9908 6920 9920
rect 5592 9880 6500 9908
rect 6875 9880 6920 9908
rect 5592 9868 5598 9880
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7190 9908 7196 9920
rect 7151 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7374 9908 7380 9920
rect 7331 9880 7380 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8036 9908 8064 9948
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 7984 9880 8064 9908
rect 8757 9911 8815 9917
rect 7984 9868 7990 9880
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9122 9908 9128 9920
rect 8803 9880 9128 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9508 9917 9536 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10244 10121 10272 10220
rect 10413 10217 10425 10251
rect 10459 10248 10471 10251
rect 10686 10248 10692 10260
rect 10459 10220 10692 10248
rect 10459 10217 10471 10220
rect 10413 10211 10471 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11330 10180 11336 10192
rect 10612 10152 11336 10180
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9877 9551 9911
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9784 9908 9812 10075
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10428 10044 10456 10075
rect 10612 10053 10640 10152
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 10870 10121 10876 10124
rect 10864 10075 10876 10121
rect 10928 10112 10934 10124
rect 10928 10084 10964 10112
rect 10870 10072 10876 10075
rect 10928 10072 10934 10084
rect 9916 10016 10456 10044
rect 10597 10047 10655 10053
rect 9916 10004 9922 10016
rect 10597 10013 10609 10047
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10612 9976 10640 10007
rect 10100 9948 10640 9976
rect 10100 9936 10106 9948
rect 9950 9908 9956 9920
rect 9784 9880 9956 9908
rect 9950 9868 9956 9880
rect 10008 9908 10014 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 10008 9880 11989 9908
rect 10008 9868 10014 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 1104 9818 12328 9840
rect 1104 9766 2852 9818
rect 2904 9766 2916 9818
rect 2968 9766 2980 9818
rect 3032 9766 3044 9818
rect 3096 9766 6594 9818
rect 6646 9766 6658 9818
rect 6710 9766 6722 9818
rect 6774 9766 6786 9818
rect 6838 9766 10335 9818
rect 10387 9766 10399 9818
rect 10451 9766 10463 9818
rect 10515 9766 10527 9818
rect 10579 9766 12328 9818
rect 1104 9744 12328 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2869 9707 2927 9713
rect 2869 9704 2881 9707
rect 1452 9676 2881 9704
rect 1452 9664 1458 9676
rect 2869 9673 2881 9676
rect 2915 9673 2927 9707
rect 2869 9667 2927 9673
rect 3252 9676 3648 9704
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9636 2007 9639
rect 2590 9636 2596 9648
rect 1995 9608 2596 9636
rect 1995 9605 2007 9608
rect 1949 9599 2007 9605
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 1084 9540 1716 9568
rect 1084 9528 1090 9540
rect 845 9503 903 9509
rect 845 9469 857 9503
rect 891 9500 903 9503
rect 1581 9503 1639 9509
rect 1581 9500 1593 9503
rect 891 9472 1593 9500
rect 891 9469 903 9472
rect 845 9463 903 9469
rect 1581 9469 1593 9472
rect 1627 9469 1639 9503
rect 1688 9500 1716 9540
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2188 9540 2513 9568
rect 2188 9528 2194 9540
rect 2501 9537 2513 9540
rect 2547 9568 2559 9571
rect 3252 9568 3280 9676
rect 3329 9639 3387 9645
rect 3329 9605 3341 9639
rect 3375 9605 3387 9639
rect 3329 9599 3387 9605
rect 2547 9540 3280 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1688 9472 1869 9500
rect 1581 9463 1639 9469
rect 1857 9469 1869 9472
rect 1903 9469 1915 9503
rect 2314 9500 2320 9512
rect 2275 9472 2320 9500
rect 1857 9463 1915 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 2648 9472 2789 9500
rect 2648 9460 2654 9472
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3344 9500 3372 9599
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3620 9568 3648 9676
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 4798 9704 4804 9716
rect 3752 9676 4804 9704
rect 3752 9664 3758 9676
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 5721 9707 5779 9713
rect 5721 9673 5733 9707
rect 5767 9704 5779 9707
rect 6178 9704 6184 9716
rect 5767 9676 6184 9704
rect 5767 9673 5779 9676
rect 5721 9667 5779 9673
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9704 6975 9707
rect 7006 9704 7012 9716
rect 6963 9676 7012 9704
rect 6963 9673 6975 9676
rect 6917 9667 6975 9673
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 7282 9704 7288 9716
rect 7116 9676 7288 9704
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 4249 9639 4307 9645
rect 4249 9636 4261 9639
rect 3936 9608 4261 9636
rect 3936 9596 3942 9608
rect 4249 9605 4261 9608
rect 4295 9605 4307 9639
rect 4614 9636 4620 9648
rect 4249 9599 4307 9605
rect 4356 9608 4620 9636
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3568 9540 3985 9568
rect 3568 9528 3574 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 4356 9568 4384 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 4948 9608 5212 9636
rect 4948 9596 4954 9608
rect 3973 9531 4031 9537
rect 4080 9540 4384 9568
rect 4433 9571 4491 9577
rect 3099 9472 3372 9500
rect 3789 9503 3847 9509
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4080 9500 4108 9540
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4479 9540 4813 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 3835 9472 4108 9500
rect 4157 9503 4215 9509
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4157 9469 4169 9503
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 3697 9435 3755 9441
rect 3697 9432 3709 9435
rect 1688 9404 3709 9432
rect 1394 9364 1400 9376
rect 1355 9336 1400 9364
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 1688 9373 1716 9404
rect 3697 9401 3709 9404
rect 3743 9401 3755 9435
rect 3697 9395 3755 9401
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9333 1731 9367
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 1673 9327 1731 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 4172 9364 4200 9463
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5184 9509 5212 9608
rect 5276 9608 6960 9636
rect 5276 9509 5304 9608
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 6730 9568 6736 9580
rect 5399 9540 5856 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 4672 9472 4721 9500
rect 4672 9460 4678 9472
rect 4709 9469 4721 9472
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9469 5319 9503
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 5261 9463 5319 9469
rect 4908 9432 4936 9463
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5828 9509 5856 9540
rect 6012 9540 6736 9568
rect 6012 9509 6040 9540
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 6178 9500 6184 9512
rect 6139 9472 6184 9500
rect 5997 9463 6055 9469
rect 5534 9432 5540 9444
rect 4908 9404 5540 9432
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 5644 9432 5672 9463
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9500 6331 9503
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 6319 9472 6469 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6457 9463 6515 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 6089 9435 6147 9441
rect 6089 9432 6101 9435
rect 5644 9404 6101 9432
rect 6089 9401 6101 9404
rect 6135 9401 6147 9435
rect 6932 9432 6960 9608
rect 7116 9577 7144 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 8938 9704 8944 9716
rect 8803 9676 8944 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 10226 9704 10232 9716
rect 9272 9676 10232 9704
rect 9272 9664 9278 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10597 9707 10655 9713
rect 10597 9673 10609 9707
rect 10643 9704 10655 9707
rect 10781 9707 10839 9713
rect 10643 9676 10677 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10781 9673 10793 9707
rect 10827 9704 10839 9707
rect 10870 9704 10876 9716
rect 10827 9676 10876 9704
rect 10827 9673 10839 9676
rect 10781 9667 10839 9673
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8444 9608 8493 9636
rect 8444 9596 8450 9608
rect 8481 9605 8493 9608
rect 8527 9636 8539 9639
rect 9582 9636 9588 9648
rect 8527 9608 9588 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 10612 9636 10640 9667
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 10560 9608 10640 9636
rect 10560 9596 10566 9608
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 9950 9568 9956 9580
rect 7101 9531 7159 9537
rect 8864 9540 9956 9568
rect 7374 9509 7380 9512
rect 7368 9500 7380 9509
rect 7335 9472 7380 9500
rect 7368 9463 7380 9472
rect 7374 9460 7380 9463
rect 7432 9460 7438 9512
rect 8864 9509 8892 9540
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10612 9568 10640 9608
rect 10778 9568 10784 9580
rect 10612 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11204 9540 11897 9568
rect 11204 9528 11210 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 8849 9463 8907 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 10134 9500 10140 9512
rect 9723 9472 10140 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10284 9472 10885 9500
rect 10284 9460 10290 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 11514 9500 11520 9512
rect 11475 9472 11520 9500
rect 10873 9463 10931 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 7650 9432 7656 9444
rect 6932 9404 7656 9432
rect 6089 9395 6147 9401
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10686 9441 10692 9444
rect 10321 9435 10379 9441
rect 10008 9404 10053 9432
rect 10008 9392 10014 9404
rect 10321 9401 10333 9435
rect 10367 9432 10379 9435
rect 10413 9435 10471 9441
rect 10413 9432 10425 9435
rect 10367 9404 10425 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 10413 9401 10425 9404
rect 10459 9401 10471 9435
rect 10413 9395 10471 9401
rect 10629 9435 10692 9441
rect 10629 9401 10641 9435
rect 10675 9401 10692 9435
rect 10629 9395 10692 9401
rect 10686 9392 10692 9395
rect 10744 9392 10750 9444
rect 4430 9364 4436 9376
rect 3191 9336 4200 9364
rect 4391 9336 4436 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5626 9364 5632 9376
rect 5031 9336 5632 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6273 9367 6331 9373
rect 6273 9364 6285 9367
rect 6052 9336 6285 9364
rect 6052 9324 6058 9336
rect 6273 9333 6285 9336
rect 6319 9333 6331 9367
rect 6273 9327 6331 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 10870 9364 10876 9376
rect 6420 9336 10876 9364
rect 6420 9324 6426 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 1104 9274 12328 9296
rect 1104 9222 4723 9274
rect 4775 9222 4787 9274
rect 4839 9222 4851 9274
rect 4903 9222 4915 9274
rect 4967 9222 8464 9274
rect 8516 9222 8528 9274
rect 8580 9222 8592 9274
rect 8644 9222 8656 9274
rect 8708 9222 12328 9274
rect 1104 9200 12328 9222
rect 1762 9160 1768 9172
rect 1412 9132 1768 9160
rect 1412 9033 1440 9132
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2464 9132 2789 9160
rect 2464 9120 2470 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 4246 9160 4252 9172
rect 2777 9123 2835 9129
rect 3528 9132 4252 9160
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 3528 9101 3556 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5442 9160 5448 9172
rect 5307 9132 5448 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5442 9120 5448 9132
rect 5500 9160 5506 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5500 9132 5825 9160
rect 5500 9120 5506 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 6144 9132 6561 9160
rect 6144 9120 6150 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 6730 9160 6736 9172
rect 6687 9132 6736 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 8352 9132 8401 9160
rect 8352 9120 8358 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 9585 9163 9643 9169
rect 9585 9129 9597 9163
rect 9631 9160 9643 9163
rect 9674 9160 9680 9172
rect 9631 9132 9680 9160
rect 9631 9129 9643 9132
rect 9585 9123 9643 9129
rect 3513 9095 3571 9101
rect 1636 9064 3372 9092
rect 1636 9052 1642 9064
rect 1670 9033 1676 9036
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1664 8987 1676 9033
rect 1728 9024 1734 9036
rect 1728 8996 1764 9024
rect 1670 8984 1676 8987
rect 1728 8984 1734 8996
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 3344 9033 3372 9064
rect 3513 9061 3525 9095
rect 3559 9061 3571 9095
rect 3513 9055 3571 9061
rect 3697 9095 3755 9101
rect 3697 9061 3709 9095
rect 3743 9092 3755 9095
rect 3878 9092 3884 9104
rect 3743 9064 3884 9092
rect 3743 9061 3755 9064
rect 3697 9055 3755 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4148 9095 4206 9101
rect 4148 9061 4160 9095
rect 4194 9092 4206 9095
rect 4430 9092 4436 9104
rect 4194 9064 4436 9092
rect 4194 9061 4206 9064
rect 4148 9055 4206 9061
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 7650 9092 7656 9104
rect 5684 9064 7656 9092
rect 5684 9052 5690 9064
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 9140 9092 9168 9123
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 9140 9064 9965 9092
rect 9953 9061 9965 9064
rect 9999 9092 10011 9095
rect 10321 9095 10379 9101
rect 9999 9064 10272 9092
rect 9999 9061 10011 9064
rect 9953 9055 10011 9061
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2280 8996 3065 9024
rect 2280 8984 2286 8996
rect 3053 8993 3065 8996
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 8993 3387 9027
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 3329 8987 3387 8993
rect 4908 8996 5733 9024
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3878 8956 3884 8968
rect 3476 8928 3884 8956
rect 3476 8916 3482 8928
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 2869 8891 2927 8897
rect 2869 8888 2881 8891
rect 2648 8860 2881 8888
rect 2648 8848 2654 8860
rect 2869 8857 2881 8860
rect 2915 8857 2927 8891
rect 2869 8851 2927 8857
rect 2976 8860 3648 8888
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 2976 8820 3004 8860
rect 1452 8792 3004 8820
rect 3145 8823 3203 8829
rect 1452 8780 1458 8792
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3510 8820 3516 8832
rect 3191 8792 3516 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3620 8820 3648 8860
rect 4908 8820 4936 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 7006 9024 7012 9036
rect 5721 8987 5779 8993
rect 5828 8996 7012 9024
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5828 8956 5856 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 5040 8928 5856 8956
rect 5997 8959 6055 8965
rect 5040 8916 5046 8928
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6086 8956 6092 8968
rect 6043 8928 6092 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6086 8916 6092 8928
rect 6144 8956 6150 8968
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 6144 8928 6745 8956
rect 6144 8916 6150 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 6822 8888 6828 8900
rect 5399 8860 6828 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7300 8888 7328 8987
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7432 8996 7573 9024
rect 7432 8984 7438 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 7561 8987 7619 8993
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8662 9024 8668 9036
rect 8623 8996 8668 9024
rect 8481 8987 8539 8993
rect 8496 8956 8524 8987
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 8938 8984 8944 9036
rect 8996 9024 9002 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8996 8996 9505 9024
rect 8996 8984 9002 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 10134 9024 10140 9036
rect 9493 8987 9551 8993
rect 9600 8996 10140 9024
rect 8849 8959 8907 8965
rect 8849 8956 8861 8959
rect 8496 8928 8861 8956
rect 8849 8925 8861 8928
rect 8895 8956 8907 8959
rect 9214 8956 9220 8968
rect 8895 8928 9220 8956
rect 8895 8925 8907 8928
rect 8849 8919 8907 8925
rect 9214 8916 9220 8928
rect 9272 8956 9278 8968
rect 9600 8956 9628 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10244 9024 10272 9064
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 10413 9095 10471 9101
rect 10413 9092 10425 9095
rect 10367 9064 10425 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 10413 9061 10425 9064
rect 10459 9061 10471 9095
rect 10413 9055 10471 9061
rect 10629 9095 10687 9101
rect 10629 9061 10641 9095
rect 10675 9092 10687 9095
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 10675 9064 10977 9092
rect 10675 9061 10687 9064
rect 10629 9055 10687 9061
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 10965 9055 11023 9061
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10244 8996 10885 9024
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 9272 8928 9628 8956
rect 9677 8959 9735 8965
rect 9272 8916 9278 8928
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 7064 8860 7328 8888
rect 7064 8848 7070 8860
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9306 8888 9312 8900
rect 8720 8860 9312 8888
rect 8720 8848 8726 8860
rect 9306 8848 9312 8860
rect 9364 8888 9370 8900
rect 9692 8888 9720 8919
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 11072 8956 11100 8987
rect 9824 8928 11100 8956
rect 9824 8916 9830 8928
rect 9364 8860 9720 8888
rect 9364 8848 9370 8860
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10560 8860 10640 8888
rect 10560 8848 10566 8860
rect 3620 8792 4936 8820
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 6270 8820 6276 8832
rect 6227 8792 6276 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 10612 8829 10640 8860
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 6972 8792 7113 8820
rect 6972 8780 6978 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 7101 8783 7159 8789
rect 10597 8823 10655 8829
rect 10597 8789 10609 8823
rect 10643 8789 10655 8823
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 10597 8783 10655 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11330 8820 11336 8832
rect 11291 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11480 8792 11621 8820
rect 11480 8780 11486 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 12066 8820 12072 8832
rect 11931 8792 12072 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 1104 8730 12328 8752
rect 1104 8678 2852 8730
rect 2904 8678 2916 8730
rect 2968 8678 2980 8730
rect 3032 8678 3044 8730
rect 3096 8678 6594 8730
rect 6646 8678 6658 8730
rect 6710 8678 6722 8730
rect 6774 8678 6786 8730
rect 6838 8678 10335 8730
rect 10387 8678 10399 8730
rect 10451 8678 10463 8730
rect 10515 8678 10527 8730
rect 10579 8678 12328 8730
rect 1104 8656 12328 8678
rect 1394 8616 1400 8628
rect 1355 8588 1400 8616
rect 1394 8576 1400 8588
rect 1452 8576 1458 8628
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1857 8619 1915 8625
rect 1857 8616 1869 8619
rect 1728 8588 1869 8616
rect 1728 8576 1734 8588
rect 1857 8585 1869 8588
rect 1903 8585 1915 8619
rect 1857 8579 1915 8585
rect 2041 8619 2099 8625
rect 2041 8585 2053 8619
rect 2087 8616 2099 8619
rect 2406 8616 2412 8628
rect 2087 8588 2412 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 3292 8588 4261 8616
rect 3292 8576 3298 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5592 8588 6776 8616
rect 5592 8576 5598 8588
rect 6748 8560 6776 8588
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 7248 8588 8401 8616
rect 7248 8576 7254 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8938 8616 8944 8628
rect 8899 8588 8944 8616
rect 8389 8579 8447 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9766 8616 9772 8628
rect 9447 8588 9772 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 9876 8588 11253 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 2866 8548 2872 8560
rect 1811 8520 2872 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1780 8480 1808 8511
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6178 8548 6184 8560
rect 6135 8520 6184 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 6178 8508 6184 8520
rect 6236 8508 6242 8560
rect 6730 8508 6736 8560
rect 6788 8508 6794 8560
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9876 8548 9904 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11241 8579 11299 8585
rect 9364 8520 9904 8548
rect 9364 8508 9370 8520
rect 1452 8452 1808 8480
rect 1949 8483 2007 8489
rect 1452 8440 1458 8452
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 1995 8452 2421 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2409 8449 2421 8452
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2608 8452 2728 8480
rect 842 8372 848 8424
rect 900 8412 906 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 900 8384 1593 8412
rect 900 8372 906 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 1728 8384 1773 8412
rect 1728 8372 1734 8384
rect 2130 8372 2136 8424
rect 2188 8412 2194 8424
rect 2608 8421 2636 8452
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2188 8384 2237 8412
rect 2188 8372 2194 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 2317 8375 2375 8381
rect 2424 8384 2513 8412
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 2332 8344 2360 8375
rect 1544 8316 2360 8344
rect 1544 8304 1550 8316
rect 2424 8294 2452 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2602 8415 2660 8421
rect 2602 8381 2614 8415
rect 2648 8381 2660 8415
rect 2602 8375 2660 8381
rect 2700 8344 2728 8452
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 4982 8480 4988 8492
rect 2832 8452 2912 8480
rect 4943 8452 4988 8480
rect 2832 8440 2838 8452
rect 2884 8421 2912 8452
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5629 8483 5687 8489
rect 5132 8452 5177 8480
rect 5132 8440 5138 8452
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 6454 8480 6460 8492
rect 5675 8452 6460 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 10137 8483 10195 8489
rect 8352 8452 8892 8480
rect 8352 8440 8358 8452
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 5166 8412 5172 8424
rect 4939 8384 5172 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5350 8412 5356 8424
rect 5311 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5534 8412 5540 8424
rect 5491 8384 5540 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 6638 8412 6644 8424
rect 5592 8384 6500 8412
rect 6599 8384 6644 8412
rect 5592 8372 5598 8384
rect 2958 8344 2964 8356
rect 2700 8316 2964 8344
rect 2498 8294 2504 8306
rect 2424 8266 2504 8294
rect 2498 8254 2504 8266
rect 2556 8276 2562 8306
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3050 8304 3056 8356
rect 3108 8353 3114 8356
rect 3108 8347 3172 8353
rect 3108 8313 3126 8347
rect 3160 8313 3172 8347
rect 3108 8307 3172 8313
rect 3108 8304 3114 8307
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 4304 8316 5917 8344
rect 4304 8304 4310 8316
rect 5184 8288 5212 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 6472 8344 6500 8384
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7098 8412 7104 8424
rect 7055 8384 7104 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 6748 8344 6776 8375
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 8864 8421 8892 8452
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10778 8480 10784 8492
rect 10183 8452 10784 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 9214 8412 9220 8424
rect 9175 8384 9220 8412
rect 8849 8375 8907 8381
rect 6822 8344 6828 8356
rect 6472 8316 6828 8344
rect 5905 8307 5963 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 6917 8347 6975 8353
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 7254 8347 7312 8353
rect 7254 8344 7266 8347
rect 6963 8316 7266 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 7254 8313 7266 8316
rect 7300 8313 7312 8347
rect 8496 8344 8524 8375
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9766 8412 9772 8424
rect 9727 8384 9772 8412
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11882 8412 11888 8424
rect 9916 8384 9961 8412
rect 11843 8384 11888 8412
rect 9916 8372 9922 8384
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 8938 8344 8944 8356
rect 8496 8316 8944 8344
rect 7254 8307 7312 8313
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 3418 8276 3424 8288
rect 2556 8254 3424 8276
rect 2516 8248 3424 8254
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 4488 8248 4537 8276
rect 4488 8236 4494 8248
rect 4525 8245 4537 8248
rect 4571 8245 4583 8279
rect 4525 8239 4583 8245
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 5626 8276 5632 8288
rect 5587 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 1104 8186 12328 8208
rect 1104 8134 4723 8186
rect 4775 8134 4787 8186
rect 4839 8134 4851 8186
rect 4903 8134 4915 8186
rect 4967 8134 8464 8186
rect 8516 8134 8528 8186
rect 8580 8134 8592 8186
rect 8644 8134 8656 8186
rect 8708 8134 12328 8186
rect 1104 8112 12328 8134
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 1964 8044 2513 8072
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 1964 8004 1992 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2501 8035 2559 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3050 8072 3056 8084
rect 3011 8044 3056 8072
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 4525 8075 4583 8081
rect 3936 8044 4384 8072
rect 3936 8032 3942 8044
rect 1728 7976 1992 8004
rect 2041 8007 2099 8013
rect 1728 7964 1734 7976
rect 2041 7973 2053 8007
rect 2087 8004 2099 8007
rect 3973 8007 4031 8013
rect 2087 7976 3280 8004
rect 2087 7973 2099 7976
rect 2041 7967 2099 7973
rect 3252 7948 3280 7976
rect 3973 7973 3985 8007
rect 4019 8004 4031 8007
rect 4246 8004 4252 8016
rect 4019 7976 4252 8004
rect 4019 7973 4031 7976
rect 3973 7967 4031 7973
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 4356 8004 4384 8044
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5350 8072 5356 8084
rect 4571 8044 5356 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6638 8072 6644 8084
rect 6411 8044 6644 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 7800 8044 8401 8072
rect 7800 8032 7806 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 9950 8072 9956 8084
rect 8389 8035 8447 8041
rect 9416 8044 9956 8072
rect 4976 8007 5034 8013
rect 4356 7976 4752 8004
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 1949 7899 2007 7905
rect 2409 7939 2467 7945
rect 2409 7905 2421 7939
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 1964 7868 1992 7899
rect 2038 7868 2044 7880
rect 1964 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2314 7868 2320 7880
rect 2271 7840 2320 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2424 7800 2452 7899
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2740 7908 2789 7936
rect 2740 7896 2746 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3234 7936 3240 7948
rect 2924 7908 2969 7936
rect 3195 7908 3240 7936
rect 2924 7896 2930 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3418 7936 3424 7948
rect 3379 7908 3424 7936
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7905 3571 7939
rect 4430 7936 4436 7948
rect 4391 7908 4436 7936
rect 3513 7899 3571 7905
rect 2685 7803 2743 7809
rect 2685 7800 2697 7803
rect 1627 7772 2452 7800
rect 2516 7772 2697 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2038 7692 2044 7744
rect 2096 7732 2102 7744
rect 2516 7732 2544 7772
rect 2685 7769 2697 7772
rect 2731 7769 2743 7803
rect 2884 7800 2912 7896
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3099 7840 3341 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3528 7868 3556 7899
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4724 7945 4752 7976
rect 4976 7973 4988 8007
rect 5022 8004 5034 8007
rect 5626 8004 5632 8016
rect 5022 7976 5632 8004
rect 5022 7973 5034 7976
rect 4976 7967 5034 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 6236 7976 6776 8004
rect 6236 7964 6242 7976
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5810 7936 5816 7948
rect 4856 7908 5816 7936
rect 4856 7896 4862 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6748 7945 6776 7976
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 9416 8004 9444 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10042 8004 10048 8016
rect 6880 7976 7052 8004
rect 6880 7964 6886 7976
rect 7024 7945 7052 7976
rect 7944 7976 9444 8004
rect 9508 7976 10048 8004
rect 7944 7945 7972 7976
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6380 7908 6561 7936
rect 3528 7840 4476 7868
rect 3329 7831 3387 7837
rect 4448 7812 4476 7840
rect 3234 7800 3240 7812
rect 2884 7772 3240 7800
rect 2685 7763 2743 7769
rect 3234 7760 3240 7772
rect 3292 7800 3298 7812
rect 4157 7803 4215 7809
rect 4157 7800 4169 7803
rect 3292 7772 4169 7800
rect 3292 7760 3298 7772
rect 4157 7769 4169 7772
rect 4203 7769 4215 7803
rect 4157 7763 4215 7769
rect 4430 7760 4436 7812
rect 4488 7760 4494 7812
rect 6380 7800 6408 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 9122 7936 9128 7948
rect 9083 7908 9128 7936
rect 7929 7899 7987 7905
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6512 7840 6653 7868
rect 6512 7828 6518 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6104 7772 6408 7800
rect 6932 7800 6960 7899
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9508 7945 9536 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10588 8007 10646 8013
rect 10588 7973 10600 8007
rect 10634 8004 10646 8007
rect 10686 8004 10692 8016
rect 10634 7976 10692 8004
rect 10634 7973 10646 7976
rect 10588 7967 10646 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 11054 7936 11060 7948
rect 9723 7908 11060 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 8352 7840 8493 7868
rect 8352 7828 8358 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 9306 7868 9312 7880
rect 8711 7840 9312 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9447 7840 9597 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9916 7840 10333 7868
rect 9916 7828 9922 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 8846 7800 8852 7812
rect 6932 7772 8852 7800
rect 6104 7744 6132 7772
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 9217 7803 9275 7809
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 9674 7800 9680 7812
rect 9263 7772 9680 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 2096 7704 2544 7732
rect 2096 7692 2102 7704
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 5442 7732 5448 7744
rect 2648 7704 5448 7732
rect 2648 7692 2654 7704
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7156 7704 7201 7732
rect 7156 7692 7162 7704
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 7653 7735 7711 7741
rect 7653 7732 7665 7735
rect 7616 7704 7665 7732
rect 7616 7692 7622 7704
rect 7653 7701 7665 7704
rect 7699 7701 7711 7735
rect 7653 7695 7711 7701
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 9030 7732 9036 7744
rect 8067 7704 9036 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9950 7732 9956 7744
rect 9364 7704 9409 7732
rect 9911 7704 9956 7732
rect 9364 7692 9370 7704
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 10192 7704 10241 7732
rect 10192 7692 10198 7704
rect 10229 7701 10241 7704
rect 10275 7701 10287 7735
rect 10229 7695 10287 7701
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11020 7704 11713 7732
rect 11020 7692 11026 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11974 7732 11980 7744
rect 11935 7704 11980 7732
rect 11701 7695 11759 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 1104 7642 12328 7664
rect 1104 7590 2852 7642
rect 2904 7590 2916 7642
rect 2968 7590 2980 7642
rect 3032 7590 3044 7642
rect 3096 7590 6594 7642
rect 6646 7590 6658 7642
rect 6710 7590 6722 7642
rect 6774 7590 6786 7642
rect 6838 7590 10335 7642
rect 10387 7590 10399 7642
rect 10451 7590 10463 7642
rect 10515 7590 10527 7642
rect 10579 7590 12328 7642
rect 1104 7568 12328 7590
rect 2682 7528 2688 7540
rect 2643 7500 2688 7528
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3476 7500 3985 7528
rect 3476 7488 3482 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 4798 7528 4804 7540
rect 3973 7491 4031 7497
rect 4080 7500 4804 7528
rect 2958 7460 2964 7472
rect 2516 7432 2964 7460
rect 1486 7324 1492 7336
rect 1447 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7284 1550 7336
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2314 7324 2320 7336
rect 2271 7296 2320 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2516 7333 2544 7432
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3050 7420 3056 7472
rect 3108 7460 3114 7472
rect 3108 7432 3153 7460
rect 3108 7420 3114 7432
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 3513 7463 3571 7469
rect 3513 7460 3525 7463
rect 3292 7432 3525 7460
rect 3292 7420 3298 7432
rect 3513 7429 3525 7432
rect 3559 7429 3571 7463
rect 3513 7423 3571 7429
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 3697 7395 3755 7401
rect 2740 7364 3004 7392
rect 2740 7352 2746 7364
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 2866 7324 2872 7336
rect 2639 7296 2872 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 2976 7324 3004 7364
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3970 7392 3976 7404
rect 3743 7364 3976 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 3237 7327 3295 7333
rect 3237 7324 3249 7327
rect 2976 7296 3249 7324
rect 3237 7293 3249 7296
rect 3283 7293 3295 7327
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3237 7287 3295 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 4080 7324 4108 7500
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5534 7528 5540 7540
rect 5215 7500 5540 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5534 7488 5540 7500
rect 5592 7528 5598 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 5592 7500 6193 7528
rect 5592 7488 5598 7500
rect 6181 7497 6193 7500
rect 6227 7528 6239 7531
rect 6362 7528 6368 7540
rect 6227 7500 6368 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 7248 7500 8401 7528
rect 7248 7488 7254 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 9582 7528 9588 7540
rect 8389 7491 8447 7497
rect 8588 7500 9588 7528
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4614 7460 4620 7472
rect 4304 7432 4620 7460
rect 4304 7420 4310 7432
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 7282 7460 7288 7472
rect 4816 7432 7288 7460
rect 4264 7364 4660 7392
rect 4264 7333 4292 7364
rect 4632 7336 4660 7364
rect 3804 7296 4108 7324
rect 4249 7327 4307 7333
rect 3804 7256 3832 7296
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7293 4583 7327
rect 4525 7287 4583 7293
rect 2056 7228 3832 7256
rect 3881 7259 3939 7265
rect 2056 7197 2084 7228
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 4430 7256 4436 7268
rect 3927 7228 4436 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 4540 7256 4568 7287
rect 4614 7284 4620 7336
rect 4672 7284 4678 7336
rect 4816 7333 4844 7432
rect 7282 7420 7288 7432
rect 7340 7420 7346 7472
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5399 7364 5825 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8588 7392 8616 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10413 7531 10471 7537
rect 10413 7497 10425 7531
rect 10459 7528 10471 7531
rect 10686 7528 10692 7540
rect 10459 7500 10692 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10318 7460 10324 7472
rect 10279 7432 10324 7460
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 8251 7364 8616 7392
rect 10505 7395 10563 7401
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 10551 7364 10977 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 11379 7364 12449 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12437 7361 12449 7364
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5534 7324 5540 7336
rect 5491 7296 5540 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5000 7256 5028 7284
rect 4540 7228 5028 7256
rect 5092 7256 5120 7287
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5718 7324 5724 7336
rect 5679 7296 5724 7324
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6178 7324 6184 7336
rect 5951 7296 6184 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 8294 7324 8300 7336
rect 8255 7296 8300 7324
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8932 7327 8990 7333
rect 8932 7293 8944 7327
rect 8978 7324 8990 7327
rect 9306 7324 9312 7336
rect 8978 7296 9312 7324
rect 8978 7293 8990 7296
rect 8932 7287 8990 7293
rect 5810 7256 5816 7268
rect 5092 7228 5816 7256
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7225 6147 7259
rect 6454 7256 6460 7268
rect 6415 7228 6460 7256
rect 6089 7219 6147 7225
rect 2041 7191 2099 7197
rect 2041 7157 2053 7191
rect 2087 7157 2099 7191
rect 2041 7151 2099 7157
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2590 7188 2596 7200
rect 2363 7160 2596 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 3694 7188 3700 7200
rect 3655 7160 3700 7188
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5626 7188 5632 7200
rect 5399 7160 5632 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6104 7188 6132 7219
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 6914 7188 6920 7200
rect 6104 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7188 6978 7200
rect 7190 7188 7196 7200
rect 6972 7160 7196 7188
rect 6972 7148 6978 7160
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8496 7188 8524 7287
rect 8680 7256 8708 7287
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10594 7324 10600 7336
rect 10275 7296 10456 7324
rect 10555 7296 10600 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 9858 7256 9864 7268
rect 8680 7228 9864 7256
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10428 7256 10456 7296
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 10870 7324 10876 7336
rect 10831 7296 10876 7324
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11054 7324 11060 7336
rect 10967 7296 11060 7324
rect 11054 7284 11060 7296
rect 11112 7324 11118 7336
rect 11238 7324 11244 7336
rect 11112 7296 11244 7324
rect 11112 7284 11118 7296
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11756 7296 11897 7324
rect 11756 7284 11762 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 10689 7259 10747 7265
rect 10689 7256 10701 7259
rect 10428 7228 10701 7256
rect 10689 7225 10701 7228
rect 10735 7225 10747 7259
rect 10689 7219 10747 7225
rect 9306 7188 9312 7200
rect 8496 7160 9312 7188
rect 9306 7148 9312 7160
rect 9364 7188 9370 7200
rect 11072 7188 11100 7284
rect 9364 7160 11100 7188
rect 9364 7148 9370 7160
rect 1104 7098 12328 7120
rect 1104 7046 4723 7098
rect 4775 7046 4787 7098
rect 4839 7046 4851 7098
rect 4903 7046 4915 7098
rect 4967 7046 8464 7098
rect 8516 7046 8528 7098
rect 8580 7046 8592 7098
rect 8644 7046 8656 7098
rect 8708 7046 12328 7098
rect 1104 7024 12328 7046
rect 2866 6984 2872 6996
rect 2827 6956 2872 6984
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 3936 6956 5396 6984
rect 3936 6944 3942 6956
rect 1854 6876 1860 6928
rect 1912 6916 1918 6928
rect 3237 6919 3295 6925
rect 3237 6916 3249 6919
rect 1912 6888 3249 6916
rect 1912 6876 1918 6888
rect 3237 6885 3249 6888
rect 3283 6885 3295 6919
rect 4246 6916 4252 6928
rect 3237 6879 3295 6885
rect 3620 6888 4252 6916
rect 1670 6857 1676 6860
rect 1664 6811 1676 6857
rect 1728 6848 1734 6860
rect 1728 6820 1764 6848
rect 1670 6808 1676 6811
rect 1728 6808 1734 6820
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2740 6820 3464 6848
rect 2740 6808 2746 6820
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 3436 6789 3464 6820
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 1268 6752 1409 6780
rect 1268 6740 1274 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 1397 6743 1455 6749
rect 2792 6752 3341 6780
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2792 6721 2820 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2648 6684 2789 6712
rect 2648 6672 2654 6684
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 3620 6644 3648 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5368 6916 5396 6956
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 6178 6984 6184 6996
rect 5776 6956 6184 6984
rect 5776 6944 5782 6956
rect 6178 6944 6184 6956
rect 6236 6984 6242 6996
rect 6733 6987 6791 6993
rect 6733 6984 6745 6987
rect 6236 6956 6745 6984
rect 6236 6944 6242 6956
rect 6733 6953 6745 6956
rect 6779 6953 6791 6987
rect 7742 6984 7748 6996
rect 6733 6947 6791 6953
rect 6840 6956 7748 6984
rect 6840 6916 6868 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 7892 6956 9781 6984
rect 7892 6944 7898 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 10042 6984 10048 6996
rect 9907 6956 10048 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10560 6956 10609 6984
rect 10560 6944 10566 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 10689 6987 10747 6993
rect 10689 6953 10701 6987
rect 10735 6984 10747 6987
rect 10870 6984 10876 6996
rect 10735 6956 10876 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 7098 6925 7104 6928
rect 7092 6916 7104 6925
rect 5368 6888 6868 6916
rect 7059 6888 7104 6916
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 5368 6857 5396 6888
rect 7092 6879 7104 6888
rect 7098 6876 7104 6879
rect 7156 6876 7162 6928
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 7248 6888 8493 6916
rect 7248 6876 7254 6888
rect 8481 6885 8493 6888
rect 8527 6885 8539 6919
rect 8481 6879 8539 6885
rect 8665 6919 8723 6925
rect 8665 6885 8677 6919
rect 8711 6916 8723 6919
rect 9674 6916 9680 6928
rect 8711 6888 9680 6916
rect 8711 6885 8723 6888
rect 8665 6879 8723 6885
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 5626 6857 5632 6860
rect 4137 6851 4195 6857
rect 4137 6848 4149 6851
rect 3752 6820 4149 6848
rect 3752 6808 3758 6820
rect 4137 6817 4149 6820
rect 4183 6817 4195 6851
rect 4137 6811 4195 6817
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6817 5411 6851
rect 5620 6848 5632 6857
rect 5587 6820 5632 6848
rect 5353 6811 5411 6817
rect 5620 6811 5632 6820
rect 5626 6808 5632 6811
rect 5684 6808 5690 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 6914 6848 6920 6860
rect 6871 6820 6920 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 6914 6808 6920 6820
rect 6972 6848 6978 6860
rect 8754 6848 8760 6860
rect 6972 6820 8294 6848
rect 8715 6820 8760 6848
rect 6972 6808 6978 6820
rect 3878 6780 3884 6792
rect 3712 6752 3884 6780
rect 3712 6724 3740 6752
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 8266 6780 8294 6820
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 8904 6820 8949 6848
rect 8904 6808 8910 6820
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 9088 6820 9137 6848
rect 9088 6808 9094 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 11057 6851 11115 6857
rect 9456 6820 10824 6848
rect 9456 6808 9462 6820
rect 8478 6780 8484 6792
rect 8266 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 9968 6789 9996 6820
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 10502 6780 10508 6792
rect 9953 6743 10011 6749
rect 10060 6752 10508 6780
rect 3694 6672 3700 6724
rect 3752 6672 3758 6724
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 8294 6712 8300 6724
rect 8251 6684 8300 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 9180 6684 9229 6712
rect 9180 6672 9186 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 9401 6715 9459 6721
rect 9401 6681 9413 6715
rect 9447 6712 9459 6715
rect 10060 6712 10088 6752
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 10796 6789 10824 6820
rect 11057 6817 11069 6851
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 11072 6712 11100 6811
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11204 6752 11529 6780
rect 11204 6740 11210 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 9447 6684 10088 6712
rect 10796 6684 11100 6712
rect 9447 6681 9459 6684
rect 9401 6675 9459 6681
rect 1636 6616 3648 6644
rect 1636 6604 1642 6616
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 3936 6616 5273 6644
rect 3936 6604 3942 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 9030 6644 9036 6656
rect 8720 6616 9036 6644
rect 8720 6604 8726 6616
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 10796 6644 10824 6684
rect 10275 6616 10824 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 11020 6616 11161 6644
rect 11020 6604 11026 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11664 6616 11805 6644
rect 11664 6604 11670 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 1104 6554 12328 6576
rect 1104 6502 2852 6554
rect 2904 6502 2916 6554
rect 2968 6502 2980 6554
rect 3032 6502 3044 6554
rect 3096 6502 6594 6554
rect 6646 6502 6658 6554
rect 6710 6502 6722 6554
rect 6774 6502 6786 6554
rect 6838 6502 10335 6554
rect 10387 6502 10399 6554
rect 10451 6502 10463 6554
rect 10515 6502 10527 6554
rect 10579 6502 12328 6554
rect 1104 6480 12328 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 1452 6412 1501 6440
rect 1452 6400 1458 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 1489 6403 1547 6409
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 2915 6412 3372 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 2700 6372 2728 6403
rect 1688 6344 2728 6372
rect 1688 6313 1716 6344
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 3234 6372 3240 6384
rect 3108 6344 3240 6372
rect 3108 6332 3114 6344
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3344 6372 3372 6412
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3476 6412 3709 6440
rect 3476 6400 3482 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3697 6403 3755 6409
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4246 6440 4252 6452
rect 4019 6412 4252 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5868 6412 5917 6440
rect 5868 6400 5874 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6420 6412 6561 6440
rect 6420 6400 6426 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 8754 6440 8760 6452
rect 7147 6412 8760 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 5350 6372 5356 6384
rect 3344 6344 5356 6372
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 8297 6375 8355 6381
rect 8297 6372 8309 6375
rect 6748 6344 8309 6372
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2682 6304 2688 6316
rect 2455 6276 2688 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3418 6304 3424 6316
rect 2792 6276 3424 6304
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2271 6208 2544 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6168 2191 6171
rect 2516 6168 2544 6208
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 2792 6245 2820 6276
rect 3418 6264 3424 6276
rect 3476 6304 3482 6316
rect 5074 6304 5080 6316
rect 3476 6276 4108 6304
rect 3476 6264 3482 6276
rect 2777 6239 2835 6245
rect 2648 6208 2693 6236
rect 2648 6196 2654 6208
rect 2777 6205 2789 6239
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 3016 6208 3065 6236
rect 3016 6196 3022 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 3292 6208 3341 6236
rect 3292 6196 3298 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 3602 6236 3608 6248
rect 3563 6208 3608 6236
rect 3329 6199 3387 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4080 6245 4108 6276
rect 4448 6276 5080 6304
rect 4448 6245 4476 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 6748 6313 6776 6344
rect 8297 6341 8309 6344
rect 8343 6341 8355 6375
rect 8297 6335 8355 6341
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5500 6276 5549 6304
rect 5500 6264 5506 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 6972 6276 7757 6304
rect 6972 6264 6978 6276
rect 7745 6273 7757 6276
rect 7791 6304 7803 6307
rect 8110 6304 8116 6316
rect 7791 6276 8116 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 9916 6276 10149 6304
rect 9916 6264 9922 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11296 6276 11928 6304
rect 11296 6264 11302 6276
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 3896 6168 3924 6196
rect 2179 6140 2452 6168
rect 2516 6140 3924 6168
rect 4172 6168 4200 6199
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4672 6208 4721 6236
rect 4672 6196 4678 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 4709 6199 4767 6205
rect 5184 6208 5825 6236
rect 5074 6168 5080 6180
rect 4172 6140 5080 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1765 6103 1823 6109
rect 1765 6100 1777 6103
rect 1728 6072 1777 6100
rect 1728 6060 1734 6072
rect 1765 6069 1777 6072
rect 1811 6069 1823 6103
rect 1765 6063 1823 6069
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2314 6100 2320 6112
rect 2096 6072 2320 6100
rect 2096 6060 2102 6072
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2424 6100 2452 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2424 6072 2881 6100
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 2869 6063 2927 6069
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5184 6100 5212 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 6362 6236 6368 6248
rect 6319 6208 6368 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 5258 6128 5264 6180
rect 5316 6168 5322 6180
rect 5353 6171 5411 6177
rect 5353 6168 5365 6171
rect 5316 6140 5365 6168
rect 5316 6128 5322 6140
rect 5353 6137 5365 6140
rect 5399 6137 5411 6171
rect 5353 6131 5411 6137
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 6086 6168 6092 6180
rect 5491 6140 6092 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 6472 6168 6500 6199
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6696 6208 6837 6236
rect 6696 6196 6702 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 7466 6236 7472 6248
rect 7427 6208 7472 6236
rect 6825 6199 6883 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7892 6208 7941 6236
rect 7892 6196 7898 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 7929 6199 7987 6205
rect 8036 6208 8217 6236
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 6472 6140 6929 6168
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 8036 6168 8064 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 9306 6236 9312 6248
rect 8435 6208 9312 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 6917 6131 6975 6137
rect 7944 6140 8064 6168
rect 7944 6112 7972 6140
rect 6730 6100 6736 6112
rect 5031 6072 5212 6100
rect 6691 6072 6736 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 7926 6100 7932 6112
rect 7607 6072 7932 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8404 6100 8432 6199
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 11900 6245 11928 6276
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11532 6208 11713 6236
rect 8748 6171 8806 6177
rect 8748 6137 8760 6171
rect 8794 6168 8806 6171
rect 8938 6168 8944 6180
rect 8794 6140 8944 6168
rect 8794 6137 8806 6140
rect 8748 6131 8806 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 10404 6171 10462 6177
rect 10404 6137 10416 6171
rect 10450 6168 10462 6171
rect 10686 6168 10692 6180
rect 10450 6140 10692 6168
rect 10450 6137 10462 6140
rect 10404 6131 10462 6137
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 8159 6072 8432 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9861 6103 9919 6109
rect 9861 6100 9873 6103
rect 9548 6072 9873 6100
rect 9548 6060 9554 6072
rect 9861 6069 9873 6072
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 11532 6109 11560 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 10652 6072 11529 6100
rect 10652 6060 10658 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11517 6063 11575 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 1104 6010 12328 6032
rect 1104 5958 4723 6010
rect 4775 5958 4787 6010
rect 4839 5958 4851 6010
rect 4903 5958 4915 6010
rect 4967 5958 8464 6010
rect 8516 5958 8528 6010
rect 8580 5958 8592 6010
rect 8644 5958 8656 6010
rect 8708 5958 12328 6010
rect 1104 5936 12328 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1452 5868 1777 5896
rect 1452 5856 1458 5868
rect 1765 5865 1777 5868
rect 1811 5865 1823 5899
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 1765 5859 1823 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3142 5896 3148 5908
rect 2915 5868 3148 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3660 5868 3893 5896
rect 3660 5856 3666 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 3881 5859 3939 5865
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 6638 5896 6644 5908
rect 5767 5868 6644 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 7374 5896 7380 5908
rect 7156 5868 7380 5896
rect 7156 5856 7162 5868
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7926 5896 7932 5908
rect 7887 5868 7932 5896
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 9306 5896 9312 5908
rect 8168 5868 9312 5896
rect 8168 5856 8174 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9769 5899 9827 5905
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 10686 5896 10692 5908
rect 9815 5868 10180 5896
rect 10647 5868 10692 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 2498 5788 2504 5840
rect 2556 5788 2562 5840
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3844 5800 4261 5828
rect 3844 5788 3850 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 5442 5828 5448 5840
rect 4249 5791 4307 5797
rect 4632 5800 5448 5828
rect 937 5763 995 5769
rect 937 5729 949 5763
rect 983 5760 995 5763
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 983 5732 1593 5760
rect 983 5729 995 5732
rect 937 5723 995 5729
rect 1581 5729 1593 5732
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 2516 5760 2544 5788
rect 2682 5760 2688 5772
rect 1728 5732 1773 5760
rect 2516 5732 2688 5760
rect 1728 5720 1734 5732
rect 2608 5701 2636 5732
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3142 5760 3148 5772
rect 3007 5732 3148 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3559 5732 4476 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 3050 5692 3056 5704
rect 3011 5664 3056 5692
rect 2593 5655 2651 5661
rect 1397 5627 1455 5633
rect 1397 5593 1409 5627
rect 1443 5624 1455 5627
rect 1578 5624 1584 5636
rect 1443 5596 1584 5624
rect 1443 5593 1455 5596
rect 1397 5587 1455 5593
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 2516 5624 2544 5655
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 4154 5692 4160 5704
rect 3283 5664 4160 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 2682 5624 2688 5636
rect 2516 5596 2688 5624
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 4448 5624 4476 5732
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4632 5692 4660 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 6178 5828 6184 5840
rect 6139 5800 6184 5828
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 6730 5788 6736 5840
rect 6788 5837 6794 5840
rect 6788 5831 6852 5837
rect 6788 5797 6806 5831
rect 6840 5797 6852 5831
rect 6788 5791 6852 5797
rect 6788 5788 6794 5791
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 8996 5800 9041 5828
rect 8996 5788 9002 5800
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 9548 5800 9904 5828
rect 9548 5788 9554 5800
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5729 4767 5763
rect 4709 5723 4767 5729
rect 4571 5664 4660 5692
rect 4724 5692 4752 5723
rect 4982 5720 4988 5772
rect 5040 5760 5046 5772
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 5040 5732 5089 5760
rect 5040 5720 5046 5732
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 5350 5760 5356 5772
rect 5311 5732 5356 5760
rect 5077 5723 5135 5729
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5166 5692 5172 5704
rect 4724 5664 5172 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5460 5692 5488 5788
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6089 5763 6147 5769
rect 6089 5760 6101 5763
rect 5960 5732 6101 5760
rect 5960 5720 5966 5732
rect 6089 5729 6101 5732
rect 6135 5729 6147 5763
rect 6546 5760 6552 5772
rect 6507 5732 6552 5760
rect 6089 5723 6147 5729
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7650 5760 7656 5772
rect 6604 5732 7656 5760
rect 6604 5720 6610 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5729 8447 5763
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8389 5723 8447 5729
rect 6178 5692 6184 5704
rect 5460 5664 6184 5692
rect 6178 5652 6184 5664
rect 6236 5692 6242 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6236 5664 6285 5692
rect 6236 5652 6242 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 5626 5624 5632 5636
rect 4448 5596 5632 5624
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 8404 5624 8432 5723
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 8711 5732 9076 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8527 5664 8953 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 9048 5692 9076 5732
rect 9122 5720 9128 5772
rect 9180 5769 9186 5772
rect 9180 5760 9191 5769
rect 9582 5760 9588 5772
rect 9180 5732 9225 5760
rect 9543 5732 9588 5760
rect 9180 5723 9191 5732
rect 9180 5720 9186 5723
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9876 5769 9904 5800
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9048 5664 9229 5692
rect 8941 5655 8999 5661
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9784 5692 9812 5723
rect 10042 5692 10048 5704
rect 9784 5664 10048 5692
rect 9217 5655 9275 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10152 5701 10180 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 10962 5828 10968 5840
rect 10428 5800 10968 5828
rect 10428 5769 10456 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11238 5828 11244 5840
rect 11103 5800 11244 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 10919 5732 11897 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 11885 5729 11897 5732
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 11790 5692 11796 5704
rect 10735 5664 11796 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 9398 5624 9404 5636
rect 8404 5596 9404 5624
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 9674 5624 9680 5636
rect 9646 5584 9680 5624
rect 9732 5624 9738 5636
rect 9953 5627 10011 5633
rect 9953 5624 9965 5627
rect 9732 5596 9965 5624
rect 9732 5584 9738 5596
rect 9953 5593 9965 5596
rect 9999 5624 10011 5627
rect 10505 5627 10563 5633
rect 10505 5624 10517 5627
rect 9999 5596 10517 5624
rect 9999 5593 10011 5596
rect 9953 5587 10011 5593
rect 10505 5593 10517 5596
rect 10551 5593 10563 5627
rect 10505 5587 10563 5593
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11333 5627 11391 5633
rect 11333 5624 11345 5627
rect 10928 5596 11345 5624
rect 10928 5584 10934 5596
rect 11333 5593 11345 5596
rect 11379 5593 11391 5627
rect 11333 5587 11391 5593
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2464 5528 2881 5556
rect 2464 5516 2470 5528
rect 2869 5525 2881 5528
rect 2915 5525 2927 5559
rect 2869 5519 2927 5525
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3234 5556 3240 5568
rect 3191 5528 3240 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 8110 5556 8116 5568
rect 6144 5528 8116 5556
rect 6144 5516 6150 5528
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8294 5556 8300 5568
rect 8255 5528 8300 5556
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 9646 5556 9674 5584
rect 8803 5528 9674 5556
rect 10045 5559 10103 5565
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 10226 5556 10232 5568
rect 10091 5528 10232 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 11020 5528 11621 5556
rect 11020 5516 11026 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 11609 5519 11667 5525
rect 1104 5466 12328 5488
rect 1104 5414 2852 5466
rect 2904 5414 2916 5466
rect 2968 5414 2980 5466
rect 3032 5414 3044 5466
rect 3096 5414 6594 5466
rect 6646 5414 6658 5466
rect 6710 5414 6722 5466
rect 6774 5414 6786 5466
rect 6838 5414 10335 5466
rect 10387 5414 10399 5466
rect 10451 5414 10463 5466
rect 10515 5414 10527 5466
rect 10579 5414 12328 5466
rect 1104 5392 12328 5414
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 2777 5355 2835 5361
rect 2777 5352 2789 5355
rect 2740 5324 2789 5352
rect 2740 5312 2746 5324
rect 2777 5321 2789 5324
rect 2823 5321 2835 5355
rect 2777 5315 2835 5321
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3142 5352 3148 5364
rect 3007 5324 3148 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4396 5324 4537 5352
rect 4396 5312 4402 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 4525 5315 4583 5321
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6273 5355 6331 5361
rect 6273 5352 6285 5355
rect 6144 5324 6285 5352
rect 6144 5312 6150 5324
rect 6273 5321 6285 5324
rect 6319 5321 6331 5355
rect 6273 5315 6331 5321
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 7834 5352 7840 5364
rect 6503 5324 7840 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 9122 5352 9128 5364
rect 8711 5324 9128 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9548 5324 9597 5352
rect 9548 5312 9554 5324
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 9585 5315 9643 5321
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 9732 5324 11529 5352
rect 9732 5312 9738 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 5258 5284 5264 5296
rect 5219 5256 5264 5284
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 6178 5244 6184 5296
rect 6236 5284 6242 5296
rect 6914 5284 6920 5296
rect 6236 5256 6920 5284
rect 6236 5244 6242 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 9306 5244 9312 5296
rect 9364 5244 9370 5296
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 2774 5216 2780 5228
rect 2464 5188 2780 5216
rect 2464 5176 2470 5188
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 6932 5216 6960 5244
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6932 5188 7113 5216
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7699 5188 8309 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8297 5179 8355 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5216 9275 5219
rect 9324 5216 9352 5244
rect 9858 5216 9864 5228
rect 9263 5188 9352 5216
rect 9416 5188 9864 5216
rect 9263 5185 9275 5188
rect 9217 5179 9275 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1443 5120 1532 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1210 4972 1216 5024
rect 1268 5012 1274 5024
rect 1504 5012 1532 5120
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2096 5120 2881 5148
rect 2096 5108 2102 5120
rect 2869 5117 2881 5120
rect 2915 5117 2927 5151
rect 2869 5111 2927 5117
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 1664 5083 1722 5089
rect 1664 5049 1676 5083
rect 1710 5080 1722 5083
rect 2406 5080 2412 5092
rect 1710 5052 2412 5080
rect 1710 5049 1722 5052
rect 1664 5043 1722 5049
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 3160 5080 3188 5111
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3401 5151 3459 5157
rect 3401 5148 3413 5151
rect 3292 5120 3413 5148
rect 3292 5108 3298 5120
rect 3401 5117 3413 5120
rect 3447 5117 3459 5151
rect 4448 5148 4476 5176
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4448 5120 4629 5148
rect 3401 5111 3459 5117
rect 4617 5117 4629 5120
rect 4663 5148 4675 5151
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 4663 5120 5641 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5629 5117 5641 5120
rect 5675 5148 5687 5151
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5675 5120 5825 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5813 5117 5825 5120
rect 5859 5148 5871 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5859 5120 6377 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6512 5120 6929 5148
rect 6512 5108 6518 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 7374 5148 7380 5160
rect 7335 5120 7380 5148
rect 6917 5111 6975 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7524 5120 7569 5148
rect 7524 5108 7530 5120
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7892 5120 7941 5148
rect 7892 5108 7898 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8435 5120 8493 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 8481 5117 8493 5120
rect 8527 5148 8539 5151
rect 8570 5148 8576 5160
rect 8527 5120 8576 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 3878 5080 3884 5092
rect 3160 5052 3884 5080
rect 3160 5012 3188 5052
rect 3878 5040 3884 5052
rect 3936 5040 3942 5092
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 4982 5080 4988 5092
rect 4488 5052 4988 5080
rect 4488 5040 4494 5052
rect 4982 5040 4988 5052
rect 5040 5080 5046 5092
rect 5077 5083 5135 5089
rect 5077 5080 5089 5083
rect 5040 5052 5089 5080
rect 5040 5040 5046 5052
rect 5077 5049 5089 5052
rect 5123 5080 5135 5083
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 5123 5052 5457 5080
rect 5123 5049 5135 5052
rect 5077 5043 5135 5049
rect 5445 5049 5457 5052
rect 5491 5049 5503 5083
rect 5445 5043 5503 5049
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5080 7067 5083
rect 8220 5080 8248 5111
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8996 5120 9045 5148
rect 8996 5108 9002 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 8754 5080 8760 5092
rect 7055 5052 8760 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 9232 5080 9260 5179
rect 9306 5108 9312 5160
rect 9364 5148 9370 5160
rect 9416 5148 9444 5188
rect 9858 5176 9864 5188
rect 9916 5216 9922 5228
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 9916 5188 10149 5216
rect 9916 5176 9922 5188
rect 10137 5185 10149 5188
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 9364 5120 9444 5148
rect 9493 5151 9551 5157
rect 9364 5108 9370 5120
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10042 5148 10048 5160
rect 9539 5120 10048 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10393 5151 10451 5157
rect 10393 5148 10405 5151
rect 10284 5120 10405 5148
rect 10284 5108 10290 5120
rect 10393 5117 10405 5120
rect 10439 5117 10451 5151
rect 10393 5111 10451 5117
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11572 5120 11805 5148
rect 11572 5108 11578 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 9674 5080 9680 5092
rect 9232 5052 9680 5080
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 9861 5083 9919 5089
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 10962 5080 10968 5092
rect 9907 5052 10968 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11977 5083 12035 5089
rect 11977 5049 11989 5083
rect 12023 5080 12035 5083
rect 13262 5080 13268 5092
rect 12023 5052 13268 5080
rect 12023 5049 12035 5052
rect 11977 5043 12035 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 1268 4984 3188 5012
rect 1268 4972 1274 4984
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 3476 4984 4813 5012
rect 3476 4972 3482 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 4801 4975 4859 4981
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5905 5015 5963 5021
rect 5905 5012 5917 5015
rect 5684 4984 5917 5012
rect 5684 4972 5690 4984
rect 5905 4981 5917 4984
rect 5951 4981 5963 5015
rect 5905 4975 5963 4981
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6914 5012 6920 5024
rect 6595 4984 6920 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7650 5012 7656 5024
rect 7611 4984 7656 5012
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7984 4984 8125 5012
rect 7984 4972 7990 4984
rect 8113 4981 8125 4984
rect 8159 5012 8171 5015
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 8159 4984 8493 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 8481 4975 8539 4981
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10226 5012 10232 5024
rect 9999 4984 10232 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 1104 4922 12328 4944
rect 1104 4870 4723 4922
rect 4775 4870 4787 4922
rect 4839 4870 4851 4922
rect 4903 4870 4915 4922
rect 4967 4870 8464 4922
rect 8516 4870 8528 4922
rect 8580 4870 8592 4922
rect 8644 4870 8656 4922
rect 8708 4870 12328 4922
rect 1104 4848 12328 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4212 4780 4353 4808
rect 4212 4768 4218 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 5258 4808 5264 4820
rect 4341 4771 4399 4777
rect 4908 4780 5264 4808
rect 2593 4743 2651 4749
rect 2593 4740 2605 4743
rect 2148 4712 2605 4740
rect 198 4632 204 4684
rect 256 4672 262 4684
rect 1489 4675 1547 4681
rect 1489 4672 1501 4675
rect 256 4644 1501 4672
rect 256 4632 262 4644
rect 1489 4641 1501 4644
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 2148 4681 2176 4712
rect 2593 4709 2605 4712
rect 2639 4709 2651 4743
rect 3418 4740 3424 4752
rect 2593 4703 2651 4709
rect 2976 4712 3424 4740
rect 1857 4675 1915 4681
rect 1857 4672 1869 4675
rect 1728 4644 1869 4672
rect 1728 4632 1734 4644
rect 1857 4641 1869 4644
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4641 2191 4675
rect 2501 4675 2559 4681
rect 2501 4672 2513 4675
rect 2133 4635 2191 4641
rect 2240 4644 2513 4672
rect 2240 4604 2268 4644
rect 2501 4641 2513 4644
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2682 4632 2688 4684
rect 2740 4672 2746 4684
rect 2976 4681 3004 4712
rect 3418 4700 3424 4712
rect 3476 4740 3482 4752
rect 4908 4749 4936 4780
rect 5258 4768 5264 4780
rect 5316 4808 5322 4820
rect 8665 4811 8723 4817
rect 5316 4780 6776 4808
rect 5316 4768 5322 4780
rect 6748 4749 6776 4780
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 8754 4808 8760 4820
rect 8711 4780 8760 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4777 9183 4811
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 9125 4771 9183 4777
rect 4893 4743 4951 4749
rect 3476 4712 4476 4740
rect 3476 4700 3482 4712
rect 2777 4675 2835 4681
rect 2777 4672 2789 4675
rect 2740 4644 2789 4672
rect 2740 4632 2746 4644
rect 2777 4641 2789 4644
rect 2823 4641 2835 4675
rect 2777 4635 2835 4641
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3602 4672 3608 4684
rect 3559 4644 3608 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 2148 4576 2268 4604
rect 2409 4607 2467 4613
rect 2148 4548 2176 4576
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2455 4576 2881 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 3252 4604 3280 4635
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3844 4644 3985 4672
rect 3844 4632 3850 4644
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 4154 4672 4160 4684
rect 4115 4644 4160 4672
rect 3973 4635 4031 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4338 4672 4344 4684
rect 4295 4644 4344 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4448 4681 4476 4712
rect 4893 4709 4905 4743
rect 4939 4709 4951 4743
rect 6733 4743 6791 4749
rect 4893 4703 4951 4709
rect 5000 4712 6684 4740
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5000 4672 5028 4712
rect 5258 4672 5264 4684
rect 4755 4644 5028 4672
rect 5092 4644 5264 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5092 4604 5120 4644
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5436 4675 5494 4681
rect 5436 4641 5448 4675
rect 5482 4672 5494 4675
rect 5482 4644 6224 4672
rect 5482 4641 5494 4644
rect 5436 4635 5494 4641
rect 6196 4616 6224 4644
rect 3252 4576 5120 4604
rect 5169 4607 5227 4613
rect 2869 4567 2927 4573
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 2130 4496 2136 4548
rect 2188 4496 2194 4548
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 3142 4536 3148 4548
rect 2271 4508 3148 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 4338 4536 4344 4548
rect 3936 4508 4344 4536
rect 3936 4496 3942 4508
rect 4338 4496 4344 4508
rect 4396 4536 4402 4548
rect 5184 4536 5212 4567
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6656 4604 6684 4712
rect 6733 4709 6745 4743
rect 6779 4709 6791 4743
rect 6733 4703 6791 4709
rect 7552 4743 7610 4749
rect 7552 4709 7564 4743
rect 7598 4740 7610 4743
rect 7650 4740 7656 4752
rect 7598 4712 7656 4740
rect 7598 4709 7610 4712
rect 7552 4703 7610 4709
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 8386 4740 8392 4752
rect 7892 4712 8392 4740
rect 7892 4700 7898 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6972 4644 7021 4672
rect 6972 4632 6978 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 8757 4675 8815 4681
rect 7009 4635 7067 4641
rect 7208 4644 8708 4672
rect 7208 4604 7236 4644
rect 6656 4576 7236 4604
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 4396 4508 5212 4536
rect 4396 4496 4402 4508
rect 6454 4496 6460 4548
rect 6512 4536 6518 4548
rect 7101 4539 7159 4545
rect 7101 4536 7113 4539
rect 6512 4508 7113 4536
rect 6512 4496 6518 4508
rect 7101 4505 7113 4508
rect 7147 4505 7159 4539
rect 7101 4499 7159 4505
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 2406 4468 2412 4480
rect 1912 4440 2412 4468
rect 1912 4428 1918 4440
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 3602 4428 3608 4480
rect 3660 4468 3666 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 3660 4440 4077 4468
rect 3660 4428 3666 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 4065 4431 4123 4437
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4672 4440 4997 4468
rect 4672 4428 4678 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 6362 4428 6368 4480
rect 6420 4468 6426 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6420 4440 6561 4468
rect 6420 4428 6426 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 6825 4471 6883 4477
rect 6825 4437 6837 4471
rect 6871 4468 6883 4471
rect 6914 4468 6920 4480
rect 6871 4440 6920 4468
rect 6871 4437 6883 4440
rect 6825 4431 6883 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7300 4468 7328 4567
rect 8680 4536 8708 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9140 4672 9168 4771
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 10100 4780 10425 4808
rect 10100 4768 10106 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 10413 4771 10471 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 9398 4700 9404 4752
rect 9456 4740 9462 4752
rect 9585 4743 9643 4749
rect 9585 4740 9597 4743
rect 9456 4712 9597 4740
rect 9456 4700 9462 4712
rect 9585 4709 9597 4712
rect 9631 4709 9643 4743
rect 9585 4703 9643 4709
rect 10686 4700 10692 4752
rect 10744 4740 10750 4752
rect 10873 4743 10931 4749
rect 10873 4740 10885 4743
rect 10744 4712 10885 4740
rect 10744 4700 10750 4712
rect 10873 4709 10885 4712
rect 10919 4709 10931 4743
rect 10873 4703 10931 4709
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11388 4712 11437 4740
rect 11388 4700 11394 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 8803 4644 9168 4672
rect 10045 4675 10103 4681
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10778 4672 10784 4684
rect 10091 4644 10784 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 10888 4644 11805 4672
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10888 4536 10916 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11020 4576 11065 4604
rect 11020 4564 11026 4576
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 12066 4604 12072 4616
rect 11388 4576 12072 4604
rect 11388 4564 11394 4576
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 8680 4508 10916 4536
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12526 4536 12532 4548
rect 12023 4508 12532 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 7558 4468 7564 4480
rect 7300 4440 7564 4468
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8849 4471 8907 4477
rect 8849 4437 8861 4471
rect 8895 4468 8907 4471
rect 8938 4468 8944 4480
rect 8895 4440 8944 4468
rect 8895 4437 8907 4440
rect 8849 4431 8907 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 10008 4440 10149 4468
rect 10008 4428 10014 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 12894 4468 12900 4480
rect 11563 4440 12900 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 1104 4378 12328 4400
rect 1104 4326 2852 4378
rect 2904 4326 2916 4378
rect 2968 4326 2980 4378
rect 3032 4326 3044 4378
rect 3096 4326 6594 4378
rect 6646 4326 6658 4378
rect 6710 4326 6722 4378
rect 6774 4326 6786 4378
rect 6838 4326 10335 4378
rect 10387 4326 10399 4378
rect 10451 4326 10463 4378
rect 10515 4326 10527 4378
rect 10579 4326 12328 4378
rect 1104 4304 12328 4326
rect 661 4267 719 4273
rect 661 4233 673 4267
rect 707 4264 719 4267
rect 1486 4264 1492 4276
rect 707 4236 1492 4264
rect 707 4233 719 4236
rect 661 4227 719 4233
rect 1486 4224 1492 4236
rect 1544 4224 1550 4276
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 2225 4267 2283 4273
rect 2225 4264 2237 4267
rect 2188 4236 2237 4264
rect 2188 4224 2194 4236
rect 2225 4233 2237 4236
rect 2271 4233 2283 4267
rect 2225 4227 2283 4233
rect 2498 4224 2504 4276
rect 2556 4264 2562 4276
rect 3421 4267 3479 4273
rect 2556 4236 2820 4264
rect 2556 4224 2562 4236
rect 753 4199 811 4205
rect 753 4165 765 4199
rect 799 4196 811 4199
rect 1118 4196 1124 4208
rect 799 4168 1124 4196
rect 799 4165 811 4168
rect 753 4159 811 4165
rect 1118 4156 1124 4168
rect 1176 4156 1182 4208
rect 106 4128 112 4140
rect 67 4100 112 4128
rect 106 4088 112 4100
rect 164 4088 170 4140
rect 382 4088 388 4140
rect 440 4128 446 4140
rect 1394 4128 1400 4140
rect 440 4100 1400 4128
rect 440 4088 446 4100
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2498 4128 2504 4140
rect 2004 4100 2504 4128
rect 2004 4088 2010 4100
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2792 4137 2820 4236
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 4614 4264 4620 4276
rect 3467 4236 4620 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 3142 4196 3148 4208
rect 2924 4168 3148 4196
rect 2924 4156 2930 4168
rect 3142 4156 3148 4168
rect 3200 4196 3206 4208
rect 3436 4196 3464 4227
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 5442 4264 5448 4276
rect 5403 4236 5448 4264
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 5997 4267 6055 4273
rect 5997 4264 6009 4267
rect 5960 4236 6009 4264
rect 5960 4224 5966 4236
rect 5997 4233 6009 4236
rect 6043 4233 6055 4267
rect 5997 4227 6055 4233
rect 6178 4224 6184 4276
rect 6236 4224 6242 4276
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6328 4236 6561 4264
rect 6328 4224 6334 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 6914 4224 6920 4276
rect 6972 4224 6978 4276
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7432 4236 7573 4264
rect 7432 4224 7438 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 9122 4264 9128 4276
rect 8435 4236 9128 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 9490 4264 9496 4276
rect 9324 4236 9496 4264
rect 6196 4196 6224 4224
rect 3200 4168 3464 4196
rect 6104 4168 6224 4196
rect 6932 4196 6960 4224
rect 7466 4196 7472 4208
rect 6932 4168 7472 4196
rect 3200 4156 3206 4168
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 3418 4128 3424 4140
rect 2777 4091 2835 4097
rect 3252 4100 3424 4128
rect 658 4020 664 4072
rect 716 4060 722 4072
rect 1118 4060 1124 4072
rect 716 4032 1124 4060
rect 716 4020 722 4032
rect 1118 4020 1124 4032
rect 1176 4020 1182 4072
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 2130 4060 2136 4072
rect 1719 4032 2136 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3050 4060 3056 4072
rect 2731 4032 3056 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3252 4069 3280 4100
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3602 4128 3608 4140
rect 3563 4100 3608 4128
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3697 4063 3755 4069
rect 3384 4032 3429 4060
rect 3384 4020 3390 4032
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 4338 4060 4344 4072
rect 3743 4032 4344 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5767 4032 6040 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 106 3952 112 4004
rect 164 3992 170 4004
rect 1489 3995 1547 4001
rect 1489 3992 1501 3995
rect 164 3964 1501 3992
rect 164 3952 170 3964
rect 1489 3961 1501 3964
rect 1535 3961 1547 3995
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 1489 3955 1547 3961
rect 1596 3964 1869 3992
rect 14 3884 20 3936
rect 72 3924 78 3936
rect 1596 3924 1624 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 1857 3955 1915 3961
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 3942 3995 4000 4001
rect 3942 3992 3954 3995
rect 3651 3964 3954 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 3942 3961 3954 3964
rect 3988 3961 4000 3995
rect 3942 3955 4000 3961
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5902 3992 5908 4004
rect 4764 3964 5908 3992
rect 4764 3952 4770 3964
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 1946 3924 1952 3936
rect 72 3896 1624 3924
rect 1907 3896 1952 3924
rect 72 3884 78 3896
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 3844 3896 5089 3924
rect 3844 3884 3850 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 6012 3924 6040 4032
rect 6104 3992 6132 4168
rect 7466 4156 7472 4168
rect 7524 4196 7530 4208
rect 9033 4199 9091 4205
rect 9033 4196 9045 4199
rect 7524 4168 9045 4196
rect 7524 4156 7530 4168
rect 9033 4165 9045 4168
rect 9079 4196 9091 4199
rect 9324 4196 9352 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9079 4168 9352 4196
rect 9079 4165 9091 4168
rect 9033 4159 9091 4165
rect 6744 4131 6802 4137
rect 6744 4097 6756 4131
rect 6790 4128 6802 4131
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6790 4100 6929 4128
rect 6790 4097 6802 4100
rect 6744 4091 6802 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7423 4100 8248 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 6270 4060 6276 4072
rect 6231 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 6454 4060 6460 4072
rect 6415 4032 6460 4060
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 6104 3964 6684 3992
rect 6178 3924 6184 3936
rect 6012 3896 6184 3924
rect 5077 3887 5135 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6656 3924 6684 3964
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7024 3992 7052 4023
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 7524 4032 7569 4060
rect 7524 4020 7530 4032
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7929 4023 7987 4029
rect 8036 4032 8125 4060
rect 6972 3964 7052 3992
rect 6972 3952 6978 3964
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 6656 3896 6745 3924
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8036 3924 8064 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8220 4060 8248 4100
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 9217 4131 9275 4137
rect 8352 4100 8708 4128
rect 8352 4088 8358 4100
rect 8680 4069 8708 4100
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 11149 4131 11207 4137
rect 9263 4100 9444 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 8665 4063 8723 4069
rect 8220 4032 8616 4060
rect 8113 4023 8171 4029
rect 8297 3995 8355 4001
rect 8297 3961 8309 3995
rect 8343 3992 8355 3995
rect 8386 3992 8392 4004
rect 8343 3964 8392 3992
rect 8343 3961 8355 3964
rect 8297 3955 8355 3961
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 8588 3992 8616 4032
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 8938 4060 8944 4072
rect 8899 4032 8944 4060
rect 8665 4023 8723 4029
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9416 4060 9444 4100
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 12618 4128 12624 4140
rect 11195 4100 12624 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 9858 4060 9864 4072
rect 9416 4032 9864 4060
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11422 4060 11428 4072
rect 11011 4032 11428 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 11882 4060 11888 4072
rect 11839 4032 11888 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 9217 3995 9275 4001
rect 8588 3964 9176 3992
rect 7984 3896 8064 3924
rect 7984 3884 7990 3896
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8757 3927 8815 3933
rect 8168 3896 8213 3924
rect 8168 3884 8174 3896
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 8938 3924 8944 3936
rect 8803 3896 8944 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9148 3924 9176 3964
rect 9217 3961 9229 3995
rect 9263 3992 9275 3995
rect 9554 3995 9612 4001
rect 9554 3992 9566 3995
rect 9263 3964 9566 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 9554 3961 9566 3964
rect 9600 3961 9612 3995
rect 11330 3992 11336 4004
rect 11291 3964 11336 3992
rect 9554 3955 9612 3961
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 11517 3995 11575 4001
rect 11517 3961 11529 3995
rect 11563 3992 11575 3995
rect 12066 3992 12072 4004
rect 11563 3964 12072 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 9306 3924 9312 3936
rect 9148 3896 9312 3924
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 10686 3924 10692 3936
rect 10647 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11756 3896 11897 3924
rect 11756 3884 11762 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 109 3859 167 3865
rect 109 3825 121 3859
rect 155 3856 167 3859
rect 382 3856 388 3868
rect 155 3828 388 3856
rect 155 3825 167 3828
rect 109 3819 167 3825
rect 382 3816 388 3828
rect 440 3816 446 3868
rect 1104 3834 12328 3856
rect 1104 3782 4723 3834
rect 4775 3782 4787 3834
rect 4839 3782 4851 3834
rect 4903 3782 4915 3834
rect 4967 3782 8464 3834
rect 8516 3782 8528 3834
rect 8580 3782 8592 3834
rect 8644 3782 8656 3834
rect 8708 3782 12328 3834
rect 1104 3760 12328 3782
rect 474 3680 480 3732
rect 532 3720 538 3732
rect 1486 3720 1492 3732
rect 532 3692 1492 3720
rect 532 3680 538 3692
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3050 3720 3056 3732
rect 2823 3692 3056 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3602 3720 3608 3732
rect 3292 3692 3608 3720
rect 3292 3680 3298 3692
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3936 3692 3985 3720
rect 3936 3680 3942 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 3973 3683 4031 3689
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 5626 3720 5632 3732
rect 4212 3692 5632 3720
rect 4212 3680 4218 3692
rect 845 3655 903 3661
rect 845 3621 857 3655
rect 891 3652 903 3655
rect 2590 3652 2596 3664
rect 891 3624 2596 3652
rect 891 3621 903 3624
rect 845 3615 903 3621
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 2746 3624 3157 3652
rect 1210 3544 1216 3596
rect 1268 3584 1274 3596
rect 1397 3587 1455 3593
rect 1397 3584 1409 3587
rect 1268 3556 1409 3584
rect 1268 3544 1274 3556
rect 1397 3553 1409 3556
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1664 3587 1722 3593
rect 1664 3553 1676 3587
rect 1710 3584 1722 3587
rect 2746 3584 2774 3624
rect 3145 3621 3157 3624
rect 3191 3621 3203 3655
rect 3145 3615 3203 3621
rect 1710 3556 2774 3584
rect 2869 3587 2927 3593
rect 1710 3553 1722 3556
rect 1664 3547 1722 3553
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3234 3584 3240 3596
rect 2915 3556 3004 3584
rect 3195 3556 3240 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 2866 3408 2872 3460
rect 2924 3408 2930 3460
rect 2976 3448 3004 3556
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 3513 3587 3571 3593
rect 3513 3584 3525 3587
rect 3476 3556 3525 3584
rect 3476 3544 3482 3556
rect 3513 3553 3525 3556
rect 3559 3553 3571 3587
rect 3878 3584 3884 3596
rect 3839 3556 3884 3584
rect 3513 3547 3571 3553
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 4356 3593 4384 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 7377 3723 7435 3729
rect 6196 3692 6859 3720
rect 5261 3655 5319 3661
rect 5261 3652 5273 3655
rect 4816 3624 5273 3652
rect 4816 3593 4844 3624
rect 5261 3621 5273 3624
rect 5307 3621 5319 3655
rect 5261 3615 5319 3621
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3553 4399 3587
rect 4341 3547 4399 3553
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 4801 3547 4859 3553
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 4172 3516 4200 3547
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5626 3584 5632 3596
rect 5587 3556 5632 3584
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3584 5963 3587
rect 6196 3584 6224 3692
rect 6733 3655 6791 3661
rect 6733 3652 6745 3655
rect 6288 3624 6745 3652
rect 6288 3593 6316 3624
rect 6733 3621 6745 3624
rect 6779 3621 6791 3655
rect 6831 3652 6859 3692
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 7466 3720 7472 3732
rect 7423 3692 7472 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7742 3720 7748 3732
rect 7703 3692 7748 3720
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8527 3692 8585 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 9674 3720 9680 3732
rect 8573 3683 8631 3689
rect 8680 3692 9260 3720
rect 9635 3692 9680 3720
rect 8680 3652 8708 3692
rect 9232 3661 9260 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10413 3723 10471 3729
rect 10413 3689 10425 3723
rect 10459 3720 10471 3723
rect 12710 3720 12716 3732
rect 10459 3692 12716 3720
rect 10459 3689 10471 3692
rect 10413 3683 10471 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 6831 3624 8708 3652
rect 9217 3655 9275 3661
rect 6733 3615 6791 3621
rect 9217 3621 9229 3655
rect 9263 3621 9275 3655
rect 9217 3615 9275 3621
rect 9416 3624 9720 3652
rect 5951 3556 6224 3584
rect 6273 3587 6331 3593
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6512 3556 6653 3584
rect 6512 3544 6518 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7742 3584 7748 3596
rect 7524 3556 7748 3584
rect 7524 3544 7530 3556
rect 7742 3544 7748 3556
rect 7800 3584 7806 3596
rect 8205 3587 8263 3593
rect 7800 3556 7972 3584
rect 7800 3544 7806 3556
rect 4430 3516 4436 3528
rect 4172 3488 4436 3516
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4672 3488 4905 3516
rect 4672 3476 4678 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5123 3488 5549 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6420 3488 6561 3516
rect 6420 3476 6426 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 7834 3516 7840 3528
rect 7795 3488 7840 3516
rect 6549 3479 6607 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 7944 3525 7972 3556
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8294 3584 8300 3596
rect 8251 3556 8300 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8444 3556 8585 3584
rect 8444 3544 8450 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 8754 3584 8760 3596
rect 8715 3556 8760 3584
rect 8573 3547 8631 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9416 3584 9444 3624
rect 9582 3584 9588 3596
rect 8987 3556 9444 3584
rect 9543 3556 9588 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9692 3584 9720 3624
rect 9766 3612 9772 3664
rect 9824 3652 9830 3664
rect 9953 3655 10011 3661
rect 9953 3652 9965 3655
rect 9824 3624 9965 3652
rect 9824 3612 9830 3624
rect 9953 3621 9965 3624
rect 9999 3621 10011 3655
rect 9953 3615 10011 3621
rect 10134 3612 10140 3664
rect 10192 3652 10198 3664
rect 10689 3655 10747 3661
rect 10689 3652 10701 3655
rect 10192 3624 10701 3652
rect 10192 3612 10198 3624
rect 10689 3621 10701 3624
rect 10735 3621 10747 3655
rect 10689 3615 10747 3621
rect 10873 3655 10931 3661
rect 10873 3621 10885 3655
rect 10919 3652 10931 3655
rect 11425 3655 11483 3661
rect 10919 3624 11376 3652
rect 10919 3621 10931 3624
rect 10873 3615 10931 3621
rect 10321 3587 10379 3593
rect 9692 3556 9812 3584
rect 9784 3528 9812 3556
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10962 3584 10968 3596
rect 10367 3556 10968 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11348 3584 11376 3624
rect 11425 3621 11437 3655
rect 11471 3652 11483 3655
rect 11606 3652 11612 3664
rect 11471 3624 11612 3652
rect 11471 3621 11483 3624
rect 11425 3615 11483 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 11974 3652 11980 3664
rect 11839 3624 11980 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12250 3584 12256 3596
rect 11348 3556 12256 3584
rect 11057 3547 11115 3553
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8168 3488 8493 3516
rect 8168 3476 8174 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9674 3516 9680 3528
rect 9447 3488 9680 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 10836 3488 11008 3516
rect 10836 3476 10842 3488
rect 10980 3460 11008 3488
rect 11072 3460 11100 3547
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11882 3516 11888 3528
rect 11287 3488 11888 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 3605 3451 3663 3457
rect 3605 3448 3617 3451
rect 2976 3420 3617 3448
rect 3605 3417 3617 3420
rect 3651 3417 3663 3451
rect 3605 3411 3663 3417
rect 6457 3451 6515 3457
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 6914 3448 6920 3460
rect 6503 3420 6920 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 6914 3408 6920 3420
rect 6972 3408 6978 3460
rect 7285 3451 7343 3457
rect 7285 3417 7297 3451
rect 7331 3448 7343 3451
rect 9582 3448 9588 3460
rect 7331 3420 9588 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 10137 3451 10195 3457
rect 10137 3417 10149 3451
rect 10183 3448 10195 3451
rect 10870 3448 10876 3460
rect 10183 3420 10876 3448
rect 10183 3417 10195 3420
rect 10137 3411 10195 3417
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 10962 3408 10968 3460
rect 11020 3408 11026 3460
rect 11054 3408 11060 3460
rect 11112 3408 11118 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 11480 3420 11989 3448
rect 11480 3408 11486 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 11977 3411 12035 3417
rect 2884 3380 2912 3408
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2884 3352 2973 3380
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 3510 3380 3516 3392
rect 3375 3352 3516 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4709 3383 4767 3389
rect 4709 3349 4721 3383
rect 4755 3380 4767 3383
rect 4890 3380 4896 3392
rect 4755 3352 4896 3380
rect 4755 3349 4767 3352
rect 4709 3343 4767 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5074 3380 5080 3392
rect 5031 3352 5080 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 6178 3380 6184 3392
rect 6139 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 6411 3352 8309 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 8297 3349 8309 3352
rect 8343 3380 8355 3383
rect 9490 3380 9496 3392
rect 8343 3352 9496 3380
rect 8343 3349 8355 3352
rect 8297 3343 8355 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11238 3380 11244 3392
rect 10836 3352 11244 3380
rect 10836 3340 10842 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 11517 3383 11575 3389
rect 11517 3380 11529 3383
rect 11388 3352 11529 3380
rect 11388 3340 11394 3352
rect 11517 3349 11529 3352
rect 11563 3349 11575 3383
rect 11517 3343 11575 3349
rect 1104 3290 12328 3312
rect 1104 3238 2852 3290
rect 2904 3238 2916 3290
rect 2968 3238 2980 3290
rect 3032 3238 3044 3290
rect 3096 3238 6594 3290
rect 6646 3238 6658 3290
rect 6710 3238 6722 3290
rect 6774 3238 6786 3290
rect 6838 3238 10335 3290
rect 10387 3238 10399 3290
rect 10451 3238 10463 3290
rect 10515 3238 10527 3290
rect 10579 3238 12328 3290
rect 1104 3216 12328 3238
rect 1946 3176 1952 3188
rect 1872 3148 1952 3176
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1872 2981 1900 3148
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 3234 3176 3240 3188
rect 2731 3148 3240 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3694 3176 3700 3188
rect 3344 3148 3700 3176
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 2866 3108 2872 3120
rect 2556 3080 2872 3108
rect 2556 3068 2562 3080
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 3344 3108 3372 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3878 3176 3884 3188
rect 3839 3148 3884 3176
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 5442 3176 5448 3188
rect 4755 3148 5448 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 5442 3136 5448 3148
rect 5500 3176 5506 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5500 3148 6193 3176
rect 5500 3136 5506 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3145 6331 3179
rect 6454 3176 6460 3188
rect 6415 3148 6460 3176
rect 6273 3139 6331 3145
rect 3160 3080 3372 3108
rect 3605 3111 3663 3117
rect 2038 3040 2044 3052
rect 1999 3012 2044 3040
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 2130 2972 2136 2984
rect 2091 2944 2136 2972
rect 1857 2935 1915 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2498 2972 2504 2984
rect 2372 2944 2504 2972
rect 2372 2932 2378 2944
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 3160 2972 3188 3080
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 4614 3108 4620 3120
rect 3651 3080 4620 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 6288 3108 6316 3139
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8849 3179 8907 3185
rect 8849 3176 8861 3179
rect 7892 3148 8861 3176
rect 7892 3136 7898 3148
rect 8849 3145 8861 3148
rect 8895 3145 8907 3179
rect 8849 3139 8907 3145
rect 9324 3148 10548 3176
rect 7466 3108 7472 3120
rect 6288 3080 7472 3108
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3789 3043 3847 3049
rect 3375 3012 3648 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3620 2984 3648 3012
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4246 3040 4252 3052
rect 3835 3012 4252 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4525 3003 4583 3009
rect 3510 2972 3516 2984
rect 3099 2944 3188 2972
rect 3471 2944 3516 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 4540 2972 4568 3003
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 7024 3049 7052 3080
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 8662 3068 8668 3120
rect 8720 3108 8726 3120
rect 9324 3108 9352 3148
rect 10520 3120 10548 3148
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11296 3148 11897 3176
rect 11296 3136 11302 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 8720 3080 9352 3108
rect 8720 3068 8726 3080
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 10410 3108 10416 3120
rect 9456 3080 10416 3108
rect 9456 3068 9462 3080
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 10502 3068 10508 3120
rect 10560 3068 10566 3120
rect 10597 3111 10655 3117
rect 10597 3077 10609 3111
rect 10643 3108 10655 3111
rect 11974 3108 11980 3120
rect 10643 3080 11980 3108
rect 10643 3077 10655 3080
rect 10597 3071 10655 3077
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6328 3012 6929 3040
rect 6328 3000 6334 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9490 3040 9496 3052
rect 9355 3012 9496 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9600 3012 11836 3040
rect 5074 2981 5080 2984
rect 5068 2972 5080 2981
rect 3660 2944 4844 2972
rect 5035 2944 5080 2972
rect 3660 2932 3666 2944
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 3878 2904 3884 2916
rect 3191 2876 3884 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 4249 2907 4307 2913
rect 4249 2904 4261 2907
rect 4120 2876 4261 2904
rect 4120 2864 4126 2876
rect 4249 2873 4261 2876
rect 4295 2873 4307 2907
rect 4249 2867 4307 2873
rect 290 2796 296 2848
rect 348 2836 354 2848
rect 2038 2836 2044 2848
rect 348 2808 2044 2836
rect 348 2796 354 2808
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 3789 2839 3847 2845
rect 3789 2805 3801 2839
rect 3835 2836 3847 2839
rect 4154 2836 4160 2848
rect 3835 2808 4160 2836
rect 3835 2805 3847 2808
rect 3789 2799 3847 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4387 2808 4721 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 4816 2836 4844 2944
rect 5068 2935 5080 2944
rect 5074 2932 5080 2935
rect 5132 2932 5138 2984
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5626 2972 5632 2984
rect 5500 2944 5632 2972
rect 5500 2932 5506 2944
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6236 2944 7389 2972
rect 6236 2932 6242 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2972 7527 2975
rect 7558 2972 7564 2984
rect 7515 2944 7564 2972
rect 7515 2941 7527 2944
rect 7469 2935 7527 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 9600 2972 9628 3012
rect 10042 2972 10048 2984
rect 7668 2944 9628 2972
rect 10003 2944 10048 2972
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 7668 2904 7696 2944
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10192 2944 10793 2972
rect 10192 2932 10198 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 11606 2972 11612 2984
rect 11011 2944 11612 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 11808 2981 11836 3012
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 4948 2876 7696 2904
rect 7736 2907 7794 2913
rect 4948 2864 4954 2876
rect 7736 2873 7748 2907
rect 7782 2904 7794 2907
rect 8386 2904 8392 2916
rect 7782 2876 8392 2904
rect 7782 2873 7794 2876
rect 7736 2867 7794 2873
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 9125 2907 9183 2913
rect 9125 2904 9137 2907
rect 8496 2876 9137 2904
rect 5626 2836 5632 2848
rect 4816 2808 5632 2836
rect 4709 2799 4767 2805
rect 5626 2796 5632 2808
rect 5684 2836 5690 2848
rect 6273 2839 6331 2845
rect 6273 2836 6285 2839
rect 5684 2808 6285 2836
rect 5684 2796 5690 2808
rect 6273 2805 6285 2808
rect 6319 2805 6331 2839
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6273 2799 6331 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 7377 2839 7435 2845
rect 7377 2805 7389 2839
rect 7423 2836 7435 2839
rect 8496 2836 8524 2876
rect 9125 2873 9137 2876
rect 9171 2873 9183 2907
rect 9125 2867 9183 2873
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 9493 2907 9551 2913
rect 9493 2904 9505 2907
rect 9364 2876 9505 2904
rect 9364 2864 9370 2876
rect 9493 2873 9505 2876
rect 9539 2873 9551 2907
rect 9493 2867 9551 2873
rect 10229 2907 10287 2913
rect 10229 2873 10241 2907
rect 10275 2904 10287 2907
rect 10318 2904 10324 2916
rect 10275 2876 10324 2904
rect 10275 2873 10287 2876
rect 10229 2867 10287 2873
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 10410 2864 10416 2916
rect 10468 2904 10474 2916
rect 11149 2907 11207 2913
rect 11149 2904 11161 2907
rect 10468 2876 10513 2904
rect 10980 2876 11161 2904
rect 10468 2864 10474 2876
rect 10980 2848 11008 2876
rect 11149 2873 11161 2876
rect 11195 2873 11207 2907
rect 11149 2867 11207 2873
rect 7423 2808 8524 2836
rect 7423 2805 7435 2808
rect 7377 2799 7435 2805
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 9456 2808 9597 2836
rect 9456 2796 9462 2808
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 11112 2808 11253 2836
rect 11112 2796 11118 2808
rect 11241 2805 11253 2808
rect 11287 2805 11299 2839
rect 11241 2799 11299 2805
rect 1104 2746 12328 2768
rect 1104 2694 4723 2746
rect 4775 2694 4787 2746
rect 4839 2694 4851 2746
rect 4903 2694 4915 2746
rect 4967 2694 8464 2746
rect 8516 2694 8528 2746
rect 8580 2694 8592 2746
rect 8644 2694 8656 2746
rect 8708 2694 12328 2746
rect 1104 2672 12328 2694
rect 753 2635 811 2641
rect 753 2601 765 2635
rect 799 2632 811 2635
rect 1118 2632 1124 2644
rect 799 2604 1124 2632
rect 799 2601 811 2604
rect 753 2595 811 2601
rect 1118 2592 1124 2604
rect 1176 2592 1182 2644
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2601 3019 2635
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 2961 2595 3019 2601
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 2866 2564 2872 2576
rect 2823 2536 2872 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 2866 2524 2872 2536
rect 2924 2524 2930 2576
rect 2976 2564 3004 2595
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5224 2604 5365 2632
rect 5224 2592 5230 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5353 2595 5411 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 6472 2604 7941 2632
rect 3418 2564 3424 2576
rect 2976 2536 3424 2564
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 4154 2573 4160 2576
rect 4148 2564 4160 2573
rect 4115 2536 4160 2564
rect 4148 2527 4160 2536
rect 4154 2524 4160 2527
rect 4212 2524 4218 2576
rect 4338 2524 4344 2576
rect 4396 2564 4402 2576
rect 5442 2564 5448 2576
rect 4396 2536 5448 2564
rect 4396 2524 4402 2536
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 6472 2564 6500 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8352 2604 8953 2632
rect 8352 2592 8358 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10045 2635 10103 2641
rect 10045 2632 10057 2635
rect 9916 2604 10057 2632
rect 9916 2592 9922 2604
rect 10045 2601 10057 2604
rect 10091 2601 10103 2635
rect 10045 2595 10103 2601
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 12342 2632 12348 2644
rect 10376 2604 12348 2632
rect 10376 2592 10382 2604
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 6196 2536 6500 2564
rect 6816 2567 6874 2573
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2130 2496 2136 2508
rect 2091 2468 2136 2496
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 3602 2496 3608 2508
rect 2731 2468 3608 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 3878 2496 3884 2508
rect 3839 2468 3884 2496
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4430 2496 4436 2508
rect 3988 2468 4436 2496
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3620 2428 3648 2456
rect 3988 2428 4016 2468
rect 4430 2456 4436 2468
rect 4488 2496 4494 2508
rect 4488 2468 5304 2496
rect 4488 2456 4494 2468
rect 3559 2400 3648 2428
rect 3896 2400 4016 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 2774 2320 2780 2372
rect 2832 2320 2838 2372
rect 3050 2320 3056 2372
rect 3108 2360 3114 2372
rect 3326 2360 3332 2372
rect 3108 2332 3332 2360
rect 3108 2320 3114 2332
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 3436 2360 3464 2391
rect 3896 2360 3924 2400
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5166 2428 5172 2440
rect 5040 2400 5172 2428
rect 5040 2388 5046 2400
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5276 2369 5304 2468
rect 5626 2456 5632 2508
rect 5684 2456 5690 2508
rect 6196 2505 6224 2536
rect 6816 2533 6828 2567
rect 6862 2564 6874 2567
rect 6914 2564 6920 2576
rect 6862 2536 6920 2564
rect 6862 2533 6874 2536
rect 6816 2527 6874 2533
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 7282 2524 7288 2576
rect 7340 2564 7346 2576
rect 7466 2564 7472 2576
rect 7340 2536 7472 2564
rect 7340 2524 7346 2536
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 8754 2564 8760 2576
rect 8435 2536 8760 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 9309 2567 9367 2573
rect 9309 2564 9321 2567
rect 9272 2536 9321 2564
rect 9272 2524 9278 2536
rect 9309 2533 9321 2536
rect 9355 2533 9367 2567
rect 9309 2527 9367 2533
rect 9582 2524 9588 2576
rect 9640 2564 9646 2576
rect 9677 2567 9735 2573
rect 9677 2564 9689 2567
rect 9640 2536 9689 2564
rect 9640 2524 9646 2536
rect 9677 2533 9689 2536
rect 9723 2533 9735 2567
rect 10594 2564 10600 2576
rect 9677 2527 9735 2533
rect 9968 2536 10600 2564
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 5859 2468 6193 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 7650 2496 7656 2508
rect 6595 2468 7656 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 5644 2428 5672 2456
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5644 2400 5917 2428
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 6380 2428 6408 2459
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8662 2496 8668 2508
rect 8527 2468 8668 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 8849 2499 8907 2505
rect 8849 2496 8861 2499
rect 8772 2468 8861 2496
rect 6380 2400 6592 2428
rect 5905 2391 5963 2397
rect 6564 2372 6592 2400
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7800 2400 8585 2428
rect 7800 2388 7806 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 3436 2332 3924 2360
rect 5261 2363 5319 2369
rect 5261 2329 5273 2363
rect 5307 2329 5319 2363
rect 5261 2323 5319 2329
rect 6546 2320 6552 2372
rect 6604 2320 6610 2372
rect 8021 2363 8079 2369
rect 8021 2329 8033 2363
rect 8067 2360 8079 2363
rect 8772 2360 8800 2468
rect 8849 2465 8861 2468
rect 8895 2465 8907 2499
rect 8849 2459 8907 2465
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 9968 2505 9996 2536
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 11057 2567 11115 2573
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 11146 2564 11152 2576
rect 11103 2536 11152 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11425 2567 11483 2573
rect 11425 2533 11437 2567
rect 11471 2564 11483 2567
rect 11514 2564 11520 2576
rect 11471 2536 11520 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9916 2468 9965 2496
rect 9916 2456 9922 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2465 10195 2499
rect 10318 2496 10324 2508
rect 10279 2468 10324 2496
rect 10137 2459 10195 2465
rect 10152 2428 10180 2459
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10560 2468 10701 2496
rect 10560 2456 10566 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 8067 2332 8800 2360
rect 8956 2400 10180 2428
rect 8067 2329 8079 2332
rect 8021 2323 8079 2329
rect 2792 2292 2820 2320
rect 3418 2292 3424 2304
rect 2792 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8956 2292 8984 2400
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 12986 2428 12992 2440
rect 10928 2400 12992 2428
rect 10928 2388 10934 2400
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 9306 2320 9312 2372
rect 9364 2360 9370 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 9364 2332 9873 2360
rect 9364 2320 9370 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 10962 2360 10968 2372
rect 10551 2332 10968 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 7984 2264 8984 2292
rect 7984 2252 7990 2264
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9180 2264 9413 2292
rect 9180 2252 9186 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 10686 2252 10692 2304
rect 10744 2292 10750 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10744 2264 10793 2292
rect 10744 2252 10750 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 10928 2264 11161 2292
rect 10928 2252 10934 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 11149 2255 11207 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 1104 2202 12328 2224
rect 1104 2150 2852 2202
rect 2904 2150 2916 2202
rect 2968 2150 2980 2202
rect 3032 2150 3044 2202
rect 3096 2150 6594 2202
rect 6646 2150 6658 2202
rect 6710 2150 6722 2202
rect 6774 2150 6786 2202
rect 6838 2150 10335 2202
rect 10387 2150 10399 2202
rect 10451 2150 10463 2202
rect 10515 2150 10527 2202
rect 10579 2150 12328 2202
rect 1104 2128 12328 2150
rect 6362 2048 6368 2100
rect 6420 2088 6426 2100
rect 6420 2060 6592 2088
rect 6420 2048 6426 2060
rect 6564 2032 6592 2060
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 4062 2020 4068 2032
rect 3016 1992 4068 2020
rect 3016 1980 3022 1992
rect 4062 1980 4068 1992
rect 4120 1980 4126 2032
rect 5902 1980 5908 2032
rect 5960 2020 5966 2032
rect 6454 2020 6460 2032
rect 5960 1992 6460 2020
rect 5960 1980 5966 1992
rect 6454 1980 6460 1992
rect 6512 1980 6518 2032
rect 6546 1980 6552 2032
rect 6604 1980 6610 2032
rect 8938 1980 8944 2032
rect 8996 2020 9002 2032
rect 10042 2020 10048 2032
rect 8996 1992 10048 2020
rect 8996 1980 9002 1992
rect 10042 1980 10048 1992
rect 10100 1980 10106 2032
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 6822 1952 6828 1964
rect 6052 1924 6828 1952
rect 6052 1912 6058 1924
rect 6822 1912 6828 1924
rect 6880 1912 6886 1964
rect 661 1819 719 1825
rect 661 1785 673 1819
rect 707 1816 719 1819
rect 6178 1816 6184 1828
rect 707 1788 6184 1816
rect 707 1785 719 1788
rect 661 1779 719 1785
rect 6178 1776 6184 1788
rect 6236 1776 6242 1828
rect 9214 1708 9220 1760
rect 9272 1748 9278 1760
rect 10410 1748 10416 1760
rect 9272 1720 10416 1748
rect 9272 1708 9278 1720
rect 10410 1708 10416 1720
rect 10468 1708 10474 1760
rect 937 1411 995 1417
rect 937 1377 949 1411
rect 983 1408 995 1411
rect 983 1380 4752 1408
rect 983 1377 995 1380
rect 937 1371 995 1377
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 4614 1340 4620 1352
rect 4304 1312 4620 1340
rect 4304 1300 4310 1312
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 4724 1340 4752 1380
rect 4798 1368 4804 1420
rect 4856 1408 4862 1420
rect 5534 1408 5540 1420
rect 4856 1380 5540 1408
rect 4856 1368 4862 1380
rect 5534 1368 5540 1380
rect 5592 1368 5598 1420
rect 7742 1368 7748 1420
rect 7800 1408 7806 1420
rect 8846 1408 8852 1420
rect 7800 1380 8852 1408
rect 7800 1368 7806 1380
rect 8846 1368 8852 1380
rect 8904 1368 8910 1420
rect 5442 1340 5448 1352
rect 4724 1312 5448 1340
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 4890 1164 4896 1216
rect 4948 1204 4954 1216
rect 6362 1204 6368 1216
rect 4948 1176 6368 1204
rect 4948 1164 4954 1176
rect 6362 1164 6368 1176
rect 6420 1164 6426 1216
rect 10778 892 10784 944
rect 10836 932 10842 944
rect 11514 932 11520 944
rect 10836 904 11520 932
rect 10836 892 10842 904
rect 11514 892 11520 904
rect 11572 892 11578 944
<< via1 >>
rect 2688 13472 2740 13524
rect 10048 13472 10100 13524
rect 664 13404 716 13456
rect 9036 13404 9088 13456
rect 480 13336 532 13388
rect 8116 13336 8168 13388
rect 2320 13200 2372 13252
rect 7932 13200 7984 13252
rect 388 13132 440 13184
rect 6184 13132 6236 13184
rect 2852 13030 2904 13082
rect 2916 13030 2968 13082
rect 2980 13030 3032 13082
rect 3044 13030 3096 13082
rect 6594 13030 6646 13082
rect 6658 13030 6710 13082
rect 6722 13030 6774 13082
rect 6786 13030 6838 13082
rect 10335 13030 10387 13082
rect 10399 13030 10451 13082
rect 10463 13030 10515 13082
rect 10527 13030 10579 13082
rect 5172 12928 5224 12980
rect 6920 12928 6972 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 3424 12860 3476 12912
rect 4344 12860 4396 12912
rect 296 12792 348 12844
rect 1860 12724 1912 12776
rect 2412 12724 2464 12776
rect 4528 12792 4580 12844
rect 5264 12792 5316 12844
rect 5448 12792 5500 12844
rect 9680 12928 9732 12980
rect 11244 12928 11296 12980
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 11152 12860 11204 12912
rect 940 12656 992 12708
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5172 12724 5224 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 6184 12724 6236 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8852 12792 8904 12844
rect 9128 12792 9180 12844
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 12624 12792 12676 12844
rect 7104 12656 7156 12708
rect 8208 12656 8260 12708
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 2044 12588 2096 12640
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 2596 12588 2648 12640
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 4252 12588 4304 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 8024 12588 8076 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 9496 12588 9548 12640
rect 11612 12656 11664 12708
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 4723 12486 4775 12538
rect 4787 12486 4839 12538
rect 4851 12486 4903 12538
rect 4915 12486 4967 12538
rect 8464 12486 8516 12538
rect 8528 12486 8580 12538
rect 8592 12486 8644 12538
rect 8656 12486 8708 12538
rect 2412 12384 2464 12436
rect 1676 12291 1728 12300
rect 1676 12257 1710 12291
rect 1710 12257 1728 12291
rect 5632 12384 5684 12436
rect 6368 12384 6420 12436
rect 3700 12359 3752 12368
rect 3700 12325 3709 12359
rect 3709 12325 3743 12359
rect 3743 12325 3752 12359
rect 3700 12316 3752 12325
rect 4252 12316 4304 12368
rect 5172 12316 5224 12368
rect 1676 12248 1728 12257
rect 4436 12248 4488 12300
rect 1768 12044 1820 12096
rect 2136 12044 2188 12096
rect 3792 12044 3844 12096
rect 5908 12248 5960 12300
rect 7288 12316 7340 12368
rect 8760 12384 8812 12436
rect 8852 12384 8904 12436
rect 9588 12384 9640 12436
rect 11612 12384 11664 12436
rect 9772 12316 9824 12368
rect 6920 12248 6972 12300
rect 8944 12248 8996 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 9864 12291 9916 12300
rect 9864 12257 9879 12291
rect 9879 12257 9913 12291
rect 9913 12257 9916 12291
rect 9864 12248 9916 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 11612 12291 11664 12300
rect 10048 12248 10100 12257
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 9404 12180 9456 12232
rect 9956 12180 10008 12232
rect 6368 12112 6420 12164
rect 8116 12112 8168 12164
rect 4988 12044 5040 12096
rect 7012 12044 7064 12096
rect 7196 12044 7248 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8944 12044 8996 12096
rect 9772 12044 9824 12096
rect 10784 12044 10836 12096
rect 2852 11942 2904 11994
rect 2916 11942 2968 11994
rect 2980 11942 3032 11994
rect 3044 11942 3096 11994
rect 6594 11942 6646 11994
rect 6658 11942 6710 11994
rect 6722 11942 6774 11994
rect 6786 11942 6838 11994
rect 10335 11942 10387 11994
rect 10399 11942 10451 11994
rect 10463 11942 10515 11994
rect 10527 11942 10579 11994
rect 1124 11840 1176 11892
rect 1768 11772 1820 11824
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2412 11636 2464 11688
rect 3792 11636 3844 11688
rect 4620 11840 4672 11892
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 5172 11840 5224 11892
rect 5816 11840 5868 11892
rect 6920 11840 6972 11892
rect 7012 11840 7064 11892
rect 9220 11840 9272 11892
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9864 11840 9916 11892
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 2780 11611 2832 11620
rect 2780 11577 2814 11611
rect 2814 11577 2832 11611
rect 5356 11772 5408 11824
rect 4528 11704 4580 11756
rect 5080 11704 5132 11756
rect 5540 11704 5592 11756
rect 4436 11679 4488 11688
rect 4436 11645 4445 11679
rect 4445 11645 4479 11679
rect 4479 11645 4488 11679
rect 4436 11636 4488 11645
rect 5724 11679 5776 11688
rect 2780 11568 2832 11577
rect 1952 11500 2004 11552
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 5632 11568 5684 11620
rect 7748 11772 7800 11824
rect 6368 11704 6420 11756
rect 6276 11679 6328 11688
rect 6276 11645 6285 11679
rect 6285 11645 6319 11679
rect 6319 11645 6328 11679
rect 6276 11636 6328 11645
rect 7196 11636 7248 11688
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 3332 11500 3384 11552
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 7288 11568 7340 11620
rect 8300 11636 8352 11688
rect 9220 11636 9272 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 9956 11636 10008 11688
rect 10508 11704 10560 11756
rect 10416 11679 10468 11688
rect 9772 11568 9824 11620
rect 5908 11500 5960 11552
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 7564 11500 7616 11552
rect 8944 11500 8996 11552
rect 10416 11645 10425 11679
rect 10425 11645 10459 11679
rect 10459 11645 10468 11679
rect 10416 11636 10468 11645
rect 10784 11704 10836 11756
rect 11152 11679 11204 11688
rect 10232 11568 10284 11620
rect 10324 11500 10376 11552
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 11520 11636 11572 11688
rect 10968 11543 11020 11552
rect 10968 11509 10977 11543
rect 10977 11509 11011 11543
rect 11011 11509 11020 11543
rect 10968 11500 11020 11509
rect 4723 11398 4775 11450
rect 4787 11398 4839 11450
rect 4851 11398 4903 11450
rect 4915 11398 4967 11450
rect 8464 11398 8516 11450
rect 8528 11398 8580 11450
rect 8592 11398 8644 11450
rect 8656 11398 8708 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2228 11296 2280 11348
rect 1952 11228 2004 11280
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 5080 11296 5132 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 5632 11296 5684 11348
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 4252 11228 4304 11280
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 2504 11024 2556 11076
rect 3608 11160 3660 11212
rect 4068 11160 4120 11212
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4344 11160 4396 11212
rect 4528 11160 4580 11212
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 5448 11160 5500 11212
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 7104 11296 7156 11348
rect 10048 11296 10100 11348
rect 10600 11296 10652 11348
rect 6552 11228 6604 11280
rect 8300 11228 8352 11280
rect 8484 11271 8536 11280
rect 8484 11237 8493 11271
rect 8493 11237 8527 11271
rect 8527 11237 8536 11271
rect 8484 11228 8536 11237
rect 8944 11228 8996 11280
rect 7288 11160 7340 11212
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 9036 11160 9088 11212
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 3884 10956 3936 11008
rect 5632 11024 5684 11076
rect 6000 11092 6052 11144
rect 5816 11024 5868 11076
rect 4804 10956 4856 11008
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 5724 10956 5776 11008
rect 6000 10956 6052 11008
rect 7932 11024 7984 11076
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 9956 11271 10008 11280
rect 9956 11237 9965 11271
rect 9965 11237 9999 11271
rect 9999 11237 10008 11271
rect 9956 11228 10008 11237
rect 10416 11160 10468 11212
rect 10876 11228 10928 11280
rect 11244 11203 11296 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 9220 10956 9272 11008
rect 9772 10956 9824 11008
rect 10232 10956 10284 11008
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 2852 10854 2904 10906
rect 2916 10854 2968 10906
rect 2980 10854 3032 10906
rect 3044 10854 3096 10906
rect 6594 10854 6646 10906
rect 6658 10854 6710 10906
rect 6722 10854 6774 10906
rect 6786 10854 6838 10906
rect 10335 10854 10387 10906
rect 10399 10854 10451 10906
rect 10463 10854 10515 10906
rect 10527 10854 10579 10906
rect 1768 10752 1820 10804
rect 4620 10752 4672 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 5816 10752 5868 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 6368 10752 6420 10804
rect 2780 10684 2832 10736
rect 5264 10684 5316 10736
rect 6828 10684 6880 10736
rect 8484 10752 8536 10804
rect 10876 10752 10928 10804
rect 11244 10752 11296 10804
rect 9680 10684 9732 10736
rect 9864 10684 9916 10736
rect 2136 10616 2188 10668
rect 2412 10616 2464 10668
rect 3792 10616 3844 10668
rect 5356 10616 5408 10668
rect 2504 10591 2556 10600
rect 112 10480 164 10532
rect 2228 10480 2280 10532
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 2872 10548 2924 10600
rect 3240 10548 3292 10600
rect 3332 10548 3384 10600
rect 4252 10591 4304 10600
rect 4252 10557 4286 10591
rect 4286 10557 4304 10591
rect 4252 10548 4304 10557
rect 4712 10548 4764 10600
rect 5540 10548 5592 10600
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 9772 10659 9824 10668
rect 2964 10480 3016 10532
rect 3700 10480 3752 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3976 10412 4028 10464
rect 4436 10480 4488 10532
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6000 10548 6052 10557
rect 6552 10548 6604 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 8852 10548 8904 10600
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 9220 10548 9272 10600
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 6828 10412 6880 10464
rect 8300 10480 8352 10532
rect 10048 10548 10100 10600
rect 10232 10548 10284 10600
rect 11152 10548 11204 10600
rect 9036 10412 9088 10464
rect 9772 10412 9824 10464
rect 10140 10412 10192 10464
rect 10232 10412 10284 10464
rect 4723 10310 4775 10362
rect 4787 10310 4839 10362
rect 4851 10310 4903 10362
rect 4915 10310 4967 10362
rect 8464 10310 8516 10362
rect 8528 10310 8580 10362
rect 8592 10310 8644 10362
rect 8656 10310 8708 10362
rect 1860 10208 1912 10260
rect 2596 10208 2648 10260
rect 2688 10208 2740 10260
rect 3148 10140 3200 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 2412 10072 2464 10124
rect 2872 10072 2924 10124
rect 3240 10072 3292 10124
rect 3332 10072 3384 10124
rect 3608 10183 3660 10192
rect 3608 10149 3617 10183
rect 3617 10149 3651 10183
rect 3651 10149 3660 10183
rect 3608 10140 3660 10149
rect 3700 10072 3752 10124
rect 4160 10208 4212 10260
rect 4436 10140 4488 10192
rect 7380 10208 7432 10260
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 2964 9936 3016 9988
rect 4160 10072 4212 10124
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 5540 10140 5592 10192
rect 4896 10072 4948 10124
rect 6000 10140 6052 10192
rect 6184 10072 6236 10124
rect 7012 10072 7064 10124
rect 8852 10208 8904 10260
rect 9680 10208 9732 10260
rect 8392 10140 8444 10192
rect 4988 9936 5040 9988
rect 8208 10072 8260 10124
rect 8668 10072 8720 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9404 10072 9456 10124
rect 3608 9868 3660 9920
rect 4068 9868 4120 9920
rect 4436 9868 4488 9920
rect 5540 9868 5592 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 7380 9868 7432 9920
rect 7932 9868 7984 9920
rect 9220 9936 9272 9988
rect 9128 9868 9180 9920
rect 9864 10140 9916 10192
rect 10692 10208 10744 10260
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 9864 10004 9916 10056
rect 11336 10140 11388 10192
rect 10876 10115 10928 10124
rect 10876 10081 10910 10115
rect 10910 10081 10928 10115
rect 10876 10072 10928 10081
rect 10048 9936 10100 9988
rect 9956 9868 10008 9920
rect 2852 9766 2904 9818
rect 2916 9766 2968 9818
rect 2980 9766 3032 9818
rect 3044 9766 3096 9818
rect 6594 9766 6646 9818
rect 6658 9766 6710 9818
rect 6722 9766 6774 9818
rect 6786 9766 6838 9818
rect 10335 9766 10387 9818
rect 10399 9766 10451 9818
rect 10463 9766 10515 9818
rect 10527 9766 10579 9818
rect 1400 9664 1452 9716
rect 2596 9596 2648 9648
rect 1032 9528 1084 9580
rect 2136 9528 2188 9580
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 2596 9460 2648 9512
rect 3516 9528 3568 9580
rect 3700 9664 3752 9716
rect 4804 9664 4856 9716
rect 6184 9664 6236 9716
rect 7012 9664 7064 9716
rect 3884 9596 3936 9648
rect 4620 9596 4672 9648
rect 4896 9596 4948 9648
rect 1400 9367 1452 9376
rect 1400 9333 1409 9367
rect 1409 9333 1443 9367
rect 1443 9333 1452 9367
rect 1400 9324 1452 9333
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 4620 9460 4672 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 6736 9528 6788 9580
rect 6184 9503 6236 9512
rect 5540 9392 5592 9444
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7288 9664 7340 9716
rect 8944 9664 8996 9716
rect 9220 9664 9272 9716
rect 10232 9664 10284 9716
rect 8392 9596 8444 9648
rect 9588 9596 9640 9648
rect 10508 9596 10560 9648
rect 10876 9664 10928 9716
rect 7380 9503 7432 9512
rect 7380 9469 7414 9503
rect 7414 9469 7432 9503
rect 7380 9460 7432 9469
rect 9956 9528 10008 9580
rect 10784 9528 10836 9580
rect 11152 9528 11204 9580
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10232 9460 10284 9512
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 7656 9392 7708 9444
rect 9956 9435 10008 9444
rect 9956 9401 9965 9435
rect 9965 9401 9999 9435
rect 9999 9401 10008 9435
rect 9956 9392 10008 9401
rect 10692 9392 10744 9444
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 5632 9324 5684 9376
rect 6000 9324 6052 9376
rect 6368 9324 6420 9376
rect 10876 9324 10928 9376
rect 4723 9222 4775 9274
rect 4787 9222 4839 9274
rect 4851 9222 4903 9274
rect 4915 9222 4967 9274
rect 8464 9222 8516 9274
rect 8528 9222 8580 9274
rect 8592 9222 8644 9274
rect 8656 9222 8708 9274
rect 1768 9120 1820 9172
rect 2412 9120 2464 9172
rect 1584 9052 1636 9104
rect 4252 9120 4304 9172
rect 5448 9120 5500 9172
rect 6092 9120 6144 9172
rect 6736 9120 6788 9172
rect 8300 9120 8352 9172
rect 1676 9027 1728 9036
rect 1676 8993 1710 9027
rect 1710 8993 1728 9027
rect 1676 8984 1728 8993
rect 2228 8984 2280 9036
rect 3884 9052 3936 9104
rect 4436 9052 4488 9104
rect 5632 9052 5684 9104
rect 7656 9052 7708 9104
rect 9680 9120 9732 9172
rect 3424 8916 3476 8968
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 3884 8916 3936 8925
rect 2596 8848 2648 8900
rect 1400 8780 1452 8832
rect 3516 8780 3568 8832
rect 7012 9027 7064 9036
rect 4988 8916 5040 8968
rect 7012 8993 7021 9027
rect 7021 8993 7055 9027
rect 7055 8993 7064 9027
rect 7012 8984 7064 8993
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 6092 8916 6144 8968
rect 6828 8848 6880 8900
rect 7012 8848 7064 8900
rect 7380 8984 7432 9036
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 8944 8984 8996 9036
rect 10140 9027 10192 9036
rect 9220 8916 9272 8968
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 8668 8848 8720 8900
rect 9312 8848 9364 8900
rect 9772 8916 9824 8968
rect 10508 8848 10560 8900
rect 6276 8780 6328 8832
rect 6920 8780 6972 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 11428 8780 11480 8832
rect 12072 8780 12124 8832
rect 2852 8678 2904 8730
rect 2916 8678 2968 8730
rect 2980 8678 3032 8730
rect 3044 8678 3096 8730
rect 6594 8678 6646 8730
rect 6658 8678 6710 8730
rect 6722 8678 6774 8730
rect 6786 8678 6838 8730
rect 10335 8678 10387 8730
rect 10399 8678 10451 8730
rect 10463 8678 10515 8730
rect 10527 8678 10579 8730
rect 1400 8619 1452 8628
rect 1400 8585 1409 8619
rect 1409 8585 1443 8619
rect 1443 8585 1452 8619
rect 1400 8576 1452 8585
rect 1676 8576 1728 8628
rect 2412 8576 2464 8628
rect 3240 8576 3292 8628
rect 5540 8576 5592 8628
rect 7196 8576 7248 8628
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 9772 8576 9824 8628
rect 1400 8440 1452 8492
rect 2872 8508 2924 8560
rect 6184 8508 6236 8560
rect 6736 8508 6788 8560
rect 9312 8508 9364 8560
rect 848 8372 900 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2136 8372 2188 8424
rect 1492 8304 1544 8356
rect 2780 8440 2832 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 6460 8440 6512 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 8300 8440 8352 8492
rect 5172 8372 5224 8424
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 5540 8372 5592 8424
rect 6644 8415 6696 8424
rect 2504 8254 2556 8306
rect 2964 8304 3016 8356
rect 3056 8304 3108 8356
rect 4252 8304 4304 8356
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7104 8372 7156 8424
rect 10784 8440 10836 8492
rect 9220 8415 9272 8424
rect 6828 8304 6880 8356
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 11888 8415 11940 8424
rect 9864 8372 9916 8381
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 8944 8304 8996 8356
rect 3424 8236 3476 8288
rect 4436 8236 4488 8288
rect 5172 8236 5224 8288
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 4723 8134 4775 8186
rect 4787 8134 4839 8186
rect 4851 8134 4903 8186
rect 4915 8134 4967 8186
rect 8464 8134 8516 8186
rect 8528 8134 8580 8186
rect 8592 8134 8644 8186
rect 8656 8134 8708 8186
rect 1676 7964 1728 8016
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 3884 8032 3936 8084
rect 4252 7964 4304 8016
rect 5356 8032 5408 8084
rect 6644 8032 6696 8084
rect 7748 8032 7800 8084
rect 2044 7828 2096 7880
rect 2320 7828 2372 7880
rect 2688 7896 2740 7948
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 3240 7939 3292 7948
rect 2872 7896 2924 7905
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 4436 7939 4488 7948
rect 2044 7692 2096 7744
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 5632 7964 5684 8016
rect 6184 7964 6236 8016
rect 4804 7896 4856 7948
rect 5816 7896 5868 7948
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6828 7964 6880 8016
rect 9956 8032 10008 8084
rect 3240 7760 3292 7812
rect 4436 7760 4488 7812
rect 9128 7939 9180 7948
rect 6460 7828 6512 7880
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 10048 7964 10100 8016
rect 10692 7964 10744 8016
rect 11060 7896 11112 7948
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 8300 7828 8352 7880
rect 9312 7828 9364 7880
rect 9864 7828 9916 7880
rect 8852 7760 8904 7812
rect 9680 7760 9732 7812
rect 2596 7692 2648 7744
rect 5448 7692 5500 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 7564 7692 7616 7744
rect 9036 7692 9088 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9956 7735 10008 7744
rect 9312 7692 9364 7701
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 10140 7692 10192 7744
rect 10968 7692 11020 7744
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 2852 7590 2904 7642
rect 2916 7590 2968 7642
rect 2980 7590 3032 7642
rect 3044 7590 3096 7642
rect 6594 7590 6646 7642
rect 6658 7590 6710 7642
rect 6722 7590 6774 7642
rect 6786 7590 6838 7642
rect 10335 7590 10387 7642
rect 10399 7590 10451 7642
rect 10463 7590 10515 7642
rect 10527 7590 10579 7642
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 3424 7488 3476 7540
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2320 7284 2372 7336
rect 2964 7420 3016 7472
rect 3056 7463 3108 7472
rect 3056 7429 3065 7463
rect 3065 7429 3099 7463
rect 3099 7429 3108 7463
rect 3056 7420 3108 7429
rect 3240 7420 3292 7472
rect 2688 7352 2740 7404
rect 2872 7284 2924 7336
rect 3976 7352 4028 7404
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4804 7488 4856 7540
rect 5540 7488 5592 7540
rect 6368 7488 6420 7540
rect 7196 7488 7248 7540
rect 4252 7420 4304 7472
rect 4620 7420 4672 7472
rect 4436 7216 4488 7268
rect 4620 7284 4672 7336
rect 7288 7420 7340 7472
rect 9588 7488 9640 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 10692 7488 10744 7540
rect 10324 7463 10376 7472
rect 10324 7429 10333 7463
rect 10333 7429 10367 7463
rect 10367 7429 10376 7463
rect 10324 7420 10376 7429
rect 4988 7284 5040 7336
rect 5540 7284 5592 7336
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 6184 7284 6236 7336
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 5816 7216 5868 7268
rect 6460 7259 6512 7268
rect 2596 7148 2648 7200
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 5632 7148 5684 7200
rect 6460 7225 6469 7259
rect 6469 7225 6503 7259
rect 6503 7225 6512 7259
rect 6460 7216 6512 7225
rect 6920 7148 6972 7200
rect 7196 7148 7248 7200
rect 9312 7284 9364 7336
rect 10600 7327 10652 7336
rect 9864 7216 9916 7268
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 11244 7284 11296 7336
rect 11704 7284 11756 7336
rect 9312 7148 9364 7200
rect 4723 7046 4775 7098
rect 4787 7046 4839 7098
rect 4851 7046 4903 7098
rect 4915 7046 4967 7098
rect 8464 7046 8516 7098
rect 8528 7046 8580 7098
rect 8592 7046 8644 7098
rect 8656 7046 8708 7098
rect 2872 6987 2924 6996
rect 2872 6953 2881 6987
rect 2881 6953 2915 6987
rect 2915 6953 2924 6987
rect 2872 6944 2924 6953
rect 3884 6944 3936 6996
rect 1860 6876 1912 6928
rect 1676 6851 1728 6860
rect 1676 6817 1710 6851
rect 1710 6817 1728 6851
rect 1676 6808 1728 6817
rect 2688 6808 2740 6860
rect 1216 6740 1268 6792
rect 2596 6672 2648 6724
rect 1584 6604 1636 6656
rect 4252 6876 4304 6928
rect 5724 6944 5776 6996
rect 6184 6944 6236 6996
rect 7748 6944 7800 6996
rect 7840 6944 7892 6996
rect 10048 6944 10100 6996
rect 10508 6944 10560 6996
rect 10876 6944 10928 6996
rect 7104 6919 7156 6928
rect 3700 6808 3752 6860
rect 7104 6885 7138 6919
rect 7138 6885 7156 6919
rect 7104 6876 7156 6885
rect 7196 6876 7248 6928
rect 9680 6876 9732 6928
rect 5632 6851 5684 6860
rect 5632 6817 5666 6851
rect 5666 6817 5684 6851
rect 5632 6808 5684 6817
rect 6920 6808 6972 6860
rect 8760 6851 8812 6860
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 9036 6808 9088 6860
rect 9404 6808 9456 6860
rect 8484 6740 8536 6792
rect 3700 6672 3752 6724
rect 8300 6672 8352 6724
rect 9128 6672 9180 6724
rect 10508 6740 10560 6792
rect 11152 6740 11204 6792
rect 3884 6604 3936 6656
rect 8668 6604 8720 6656
rect 9036 6604 9088 6656
rect 10968 6604 11020 6656
rect 11612 6604 11664 6656
rect 2852 6502 2904 6554
rect 2916 6502 2968 6554
rect 2980 6502 3032 6554
rect 3044 6502 3096 6554
rect 6594 6502 6646 6554
rect 6658 6502 6710 6554
rect 6722 6502 6774 6554
rect 6786 6502 6838 6554
rect 10335 6502 10387 6554
rect 10399 6502 10451 6554
rect 10463 6502 10515 6554
rect 10527 6502 10579 6554
rect 1400 6400 1452 6452
rect 1676 6400 1728 6452
rect 3056 6332 3108 6384
rect 3240 6332 3292 6384
rect 3424 6400 3476 6452
rect 4252 6400 4304 6452
rect 5816 6400 5868 6452
rect 6368 6400 6420 6452
rect 8760 6400 8812 6452
rect 5356 6332 5408 6384
rect 2688 6264 2740 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 3424 6264 3476 6316
rect 2596 6196 2648 6205
rect 2964 6196 3016 6248
rect 3240 6196 3292 6248
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 5080 6264 5132 6316
rect 5448 6264 5500 6316
rect 6920 6264 6972 6316
rect 8116 6264 8168 6316
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 9864 6264 9916 6316
rect 11244 6264 11296 6316
rect 4620 6196 4672 6248
rect 1676 6060 1728 6112
rect 2044 6060 2096 6112
rect 2320 6060 2372 6112
rect 5080 6128 5132 6180
rect 6368 6196 6420 6248
rect 5264 6128 5316 6180
rect 6092 6128 6144 6180
rect 6644 6196 6696 6248
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 7840 6196 7892 6248
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 7932 6060 7984 6112
rect 9312 6196 9364 6248
rect 8944 6128 8996 6180
rect 10692 6128 10744 6180
rect 9496 6060 9548 6112
rect 10600 6060 10652 6112
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 4723 5958 4775 6010
rect 4787 5958 4839 6010
rect 4851 5958 4903 6010
rect 4915 5958 4967 6010
rect 8464 5958 8516 6010
rect 8528 5958 8580 6010
rect 8592 5958 8644 6010
rect 8656 5958 8708 6010
rect 1400 5856 1452 5908
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 3148 5856 3200 5908
rect 3608 5856 3660 5908
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 6644 5856 6696 5908
rect 7104 5856 7156 5908
rect 7380 5856 7432 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 8116 5856 8168 5908
rect 9312 5856 9364 5908
rect 10692 5899 10744 5908
rect 2504 5788 2556 5840
rect 3792 5788 3844 5840
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 2688 5720 2740 5772
rect 3148 5720 3200 5772
rect 3056 5695 3108 5704
rect 1584 5584 1636 5636
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 4160 5652 4212 5704
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 2688 5584 2740 5636
rect 5448 5788 5500 5840
rect 6184 5831 6236 5840
rect 6184 5797 6193 5831
rect 6193 5797 6227 5831
rect 6227 5797 6236 5831
rect 6184 5788 6236 5797
rect 6736 5788 6788 5840
rect 8944 5831 8996 5840
rect 8944 5797 8953 5831
rect 8953 5797 8987 5831
rect 8987 5797 8996 5831
rect 8944 5788 8996 5797
rect 9496 5788 9548 5840
rect 4988 5720 5040 5772
rect 5356 5763 5408 5772
rect 5356 5729 5365 5763
rect 5365 5729 5399 5763
rect 5399 5729 5408 5763
rect 5356 5720 5408 5729
rect 5172 5652 5224 5704
rect 5908 5720 5960 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7656 5720 7708 5772
rect 8576 5763 8628 5772
rect 6184 5652 6236 5704
rect 5632 5584 5684 5636
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9128 5763 9180 5772
rect 9128 5729 9145 5763
rect 9145 5729 9179 5763
rect 9179 5729 9180 5763
rect 9588 5763 9640 5772
rect 9128 5720 9180 5729
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 10048 5652 10100 5704
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 10968 5788 11020 5840
rect 11244 5788 11296 5840
rect 11796 5652 11848 5704
rect 9404 5584 9456 5636
rect 9680 5584 9732 5636
rect 10876 5584 10928 5636
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 2412 5516 2464 5568
rect 3240 5516 3292 5568
rect 6092 5516 6144 5568
rect 8116 5516 8168 5568
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 10232 5516 10284 5568
rect 10968 5516 11020 5568
rect 2852 5414 2904 5466
rect 2916 5414 2968 5466
rect 2980 5414 3032 5466
rect 3044 5414 3096 5466
rect 6594 5414 6646 5466
rect 6658 5414 6710 5466
rect 6722 5414 6774 5466
rect 6786 5414 6838 5466
rect 10335 5414 10387 5466
rect 10399 5414 10451 5466
rect 10463 5414 10515 5466
rect 10527 5414 10579 5466
rect 2688 5312 2740 5364
rect 3148 5312 3200 5364
rect 4344 5312 4396 5364
rect 6092 5312 6144 5364
rect 7840 5312 7892 5364
rect 9128 5312 9180 5364
rect 9496 5312 9548 5364
rect 9680 5312 9732 5364
rect 5264 5287 5316 5296
rect 5264 5253 5273 5287
rect 5273 5253 5307 5287
rect 5307 5253 5316 5287
rect 5264 5244 5316 5253
rect 6184 5244 6236 5296
rect 6920 5244 6972 5296
rect 9312 5244 9364 5296
rect 2412 5176 2464 5228
rect 2780 5176 2832 5228
rect 4436 5176 4488 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 1216 4972 1268 5024
rect 2044 5108 2096 5160
rect 2412 5040 2464 5092
rect 3240 5108 3292 5160
rect 6460 5108 6512 5160
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 7840 5108 7892 5160
rect 3884 5040 3936 5092
rect 4436 5040 4488 5092
rect 4988 5040 5040 5092
rect 8576 5108 8628 5160
rect 8944 5108 8996 5160
rect 8760 5040 8812 5092
rect 9312 5108 9364 5160
rect 9864 5176 9916 5228
rect 10048 5108 10100 5160
rect 10232 5108 10284 5160
rect 11520 5108 11572 5160
rect 9680 5040 9732 5092
rect 10968 5040 11020 5092
rect 13268 5040 13320 5092
rect 3424 4972 3476 5024
rect 5632 4972 5684 5024
rect 6920 4972 6972 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 7932 4972 7984 5024
rect 10232 4972 10284 5024
rect 4723 4870 4775 4922
rect 4787 4870 4839 4922
rect 4851 4870 4903 4922
rect 4915 4870 4967 4922
rect 8464 4870 8516 4922
rect 8528 4870 8580 4922
rect 8592 4870 8644 4922
rect 8656 4870 8708 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 4160 4768 4212 4820
rect 204 4632 256 4684
rect 1676 4632 1728 4684
rect 2688 4632 2740 4684
rect 3424 4700 3476 4752
rect 5264 4768 5316 4820
rect 8760 4768 8812 4820
rect 9496 4811 9548 4820
rect 3608 4632 3660 4684
rect 3792 4632 3844 4684
rect 4160 4675 4212 4684
rect 4160 4641 4169 4675
rect 4169 4641 4203 4675
rect 4203 4641 4212 4675
rect 4160 4632 4212 4641
rect 4344 4632 4396 4684
rect 5264 4632 5316 4684
rect 2136 4496 2188 4548
rect 3148 4496 3200 4548
rect 3884 4496 3936 4548
rect 4344 4496 4396 4548
rect 6184 4564 6236 4616
rect 7656 4700 7708 4752
rect 7840 4700 7892 4752
rect 8392 4700 8444 4752
rect 6920 4632 6972 4684
rect 6460 4496 6512 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 1860 4428 1912 4480
rect 2412 4428 2464 4480
rect 3608 4428 3660 4480
rect 4620 4428 4672 4480
rect 6368 4428 6420 4480
rect 6920 4428 6972 4480
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 10048 4768 10100 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 9404 4700 9456 4752
rect 10692 4700 10744 4752
rect 11336 4700 11388 4752
rect 10784 4632 10836 4684
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 11336 4564 11388 4616
rect 12072 4564 12124 4616
rect 12532 4496 12584 4548
rect 7564 4428 7616 4480
rect 8944 4428 8996 4480
rect 9956 4428 10008 4480
rect 12900 4428 12952 4480
rect 2852 4326 2904 4378
rect 2916 4326 2968 4378
rect 2980 4326 3032 4378
rect 3044 4326 3096 4378
rect 6594 4326 6646 4378
rect 6658 4326 6710 4378
rect 6722 4326 6774 4378
rect 6786 4326 6838 4378
rect 10335 4326 10387 4378
rect 10399 4326 10451 4378
rect 10463 4326 10515 4378
rect 10527 4326 10579 4378
rect 1492 4224 1544 4276
rect 2136 4224 2188 4276
rect 2504 4224 2556 4276
rect 1124 4156 1176 4208
rect 112 4131 164 4140
rect 112 4097 121 4131
rect 121 4097 155 4131
rect 155 4097 164 4131
rect 112 4088 164 4097
rect 388 4088 440 4140
rect 1400 4088 1452 4140
rect 1952 4088 2004 4140
rect 2504 4088 2556 4140
rect 2872 4156 2924 4208
rect 3148 4156 3200 4208
rect 4620 4224 4672 4276
rect 5448 4267 5500 4276
rect 5448 4233 5457 4267
rect 5457 4233 5491 4267
rect 5491 4233 5500 4267
rect 5448 4224 5500 4233
rect 5908 4224 5960 4276
rect 6184 4224 6236 4276
rect 6276 4224 6328 4276
rect 6920 4224 6972 4276
rect 7380 4224 7432 4276
rect 9128 4224 9180 4276
rect 664 4020 716 4072
rect 1124 4020 1176 4072
rect 2136 4020 2188 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3424 4088 3476 4140
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 4344 4020 4396 4072
rect 112 3952 164 4004
rect 20 3884 72 3936
rect 4712 3952 4764 4004
rect 5908 3952 5960 4004
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 3792 3884 3844 3936
rect 7472 4156 7524 4208
rect 9496 4224 9548 4276
rect 6276 4063 6328 4072
rect 6276 4029 6285 4063
rect 6285 4029 6319 4063
rect 6319 4029 6328 4063
rect 6276 4020 6328 4029
rect 6460 4063 6512 4072
rect 6460 4029 6469 4063
rect 6469 4029 6503 4063
rect 6503 4029 6512 4063
rect 6460 4020 6512 4029
rect 6644 4020 6696 4072
rect 6184 3884 6236 3936
rect 6920 3952 6972 4004
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7840 4020 7892 4072
rect 7932 3884 7984 3936
rect 8300 4088 8352 4140
rect 8392 3952 8444 4004
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 12624 4088 12676 4140
rect 9864 4020 9916 4072
rect 11428 4020 11480 4072
rect 11888 4020 11940 4072
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 8944 3884 8996 3936
rect 11336 3995 11388 4004
rect 11336 3961 11345 3995
rect 11345 3961 11379 3995
rect 11379 3961 11388 3995
rect 11336 3952 11388 3961
rect 12072 3952 12124 4004
rect 9312 3884 9364 3936
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 11704 3884 11756 3936
rect 388 3816 440 3868
rect 4723 3782 4775 3834
rect 4787 3782 4839 3834
rect 4851 3782 4903 3834
rect 4915 3782 4967 3834
rect 8464 3782 8516 3834
rect 8528 3782 8580 3834
rect 8592 3782 8644 3834
rect 8656 3782 8708 3834
rect 480 3680 532 3732
rect 1492 3680 1544 3732
rect 3056 3680 3108 3732
rect 3240 3680 3292 3732
rect 3608 3680 3660 3732
rect 3884 3680 3936 3732
rect 4160 3680 4212 3732
rect 2596 3612 2648 3664
rect 1216 3544 1268 3596
rect 3240 3587 3292 3596
rect 2872 3408 2924 3460
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 3424 3544 3476 3596
rect 3884 3587 3936 3596
rect 3884 3553 3893 3587
rect 3893 3553 3927 3587
rect 3927 3553 3936 3587
rect 3884 3544 3936 3553
rect 5632 3680 5684 3732
rect 5172 3587 5224 3596
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 7472 3680 7524 3732
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 12716 3680 12768 3732
rect 6460 3544 6512 3596
rect 7472 3544 7524 3596
rect 7748 3544 7800 3596
rect 4436 3476 4488 3528
rect 4620 3476 4672 3528
rect 6368 3476 6420 3528
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8300 3544 8352 3596
rect 8392 3544 8444 3596
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 9772 3612 9824 3664
rect 10140 3612 10192 3664
rect 10968 3544 11020 3596
rect 11612 3612 11664 3664
rect 11980 3612 12032 3664
rect 8116 3476 8168 3528
rect 9680 3476 9732 3528
rect 9772 3476 9824 3528
rect 10784 3476 10836 3528
rect 12256 3544 12308 3596
rect 11888 3476 11940 3528
rect 6920 3408 6972 3460
rect 9588 3408 9640 3460
rect 10876 3408 10928 3460
rect 10968 3408 11020 3460
rect 11060 3408 11112 3460
rect 11428 3408 11480 3460
rect 3516 3340 3568 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 4896 3340 4948 3392
rect 5080 3340 5132 3392
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 9496 3340 9548 3392
rect 10784 3340 10836 3392
rect 11244 3340 11296 3392
rect 11336 3340 11388 3392
rect 2852 3238 2904 3290
rect 2916 3238 2968 3290
rect 2980 3238 3032 3290
rect 3044 3238 3096 3290
rect 6594 3238 6646 3290
rect 6658 3238 6710 3290
rect 6722 3238 6774 3290
rect 6786 3238 6838 3290
rect 10335 3238 10387 3290
rect 10399 3238 10451 3290
rect 10463 3238 10515 3290
rect 10527 3238 10579 3290
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 1952 3136 2004 3188
rect 3240 3136 3292 3188
rect 2504 3068 2556 3120
rect 2872 3068 2924 3120
rect 3700 3136 3752 3188
rect 3884 3179 3936 3188
rect 3884 3145 3893 3179
rect 3893 3145 3927 3179
rect 3927 3145 3936 3179
rect 3884 3136 3936 3145
rect 5448 3136 5500 3188
rect 6460 3179 6512 3188
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 2320 2932 2372 2984
rect 2504 2932 2556 2984
rect 4620 3068 4672 3120
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 7840 3136 7892 3188
rect 4252 3000 4304 3052
rect 4804 3043 4856 3052
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 3608 2932 3660 2984
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 6276 3000 6328 3052
rect 7472 3068 7524 3120
rect 8668 3068 8720 3120
rect 11244 3136 11296 3188
rect 9404 3068 9456 3120
rect 10416 3068 10468 3120
rect 10508 3068 10560 3120
rect 11980 3068 12032 3120
rect 9496 3000 9548 3052
rect 5080 2975 5132 2984
rect 3884 2864 3936 2916
rect 4068 2864 4120 2916
rect 296 2796 348 2848
rect 2044 2796 2096 2848
rect 4160 2796 4212 2848
rect 5080 2941 5114 2975
rect 5114 2941 5132 2975
rect 5080 2932 5132 2941
rect 5448 2932 5500 2984
rect 5632 2932 5684 2984
rect 6184 2932 6236 2984
rect 7564 2932 7616 2984
rect 10048 2975 10100 2984
rect 4896 2864 4948 2916
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 10140 2932 10192 2984
rect 11612 2932 11664 2984
rect 8392 2864 8444 2916
rect 5632 2796 5684 2848
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 9312 2864 9364 2916
rect 10324 2864 10376 2916
rect 10416 2907 10468 2916
rect 10416 2873 10425 2907
rect 10425 2873 10459 2907
rect 10459 2873 10468 2907
rect 10416 2864 10468 2873
rect 9404 2796 9456 2848
rect 10968 2796 11020 2848
rect 11060 2796 11112 2848
rect 4723 2694 4775 2746
rect 4787 2694 4839 2746
rect 4851 2694 4903 2746
rect 4915 2694 4967 2746
rect 8464 2694 8516 2746
rect 8528 2694 8580 2746
rect 8592 2694 8644 2746
rect 8656 2694 8708 2746
rect 1124 2592 1176 2644
rect 3332 2635 3384 2644
rect 2872 2524 2924 2576
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 5172 2592 5224 2644
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 3424 2524 3476 2576
rect 4160 2567 4212 2576
rect 4160 2533 4194 2567
rect 4194 2533 4212 2567
rect 4160 2524 4212 2533
rect 4344 2524 4396 2576
rect 5448 2524 5500 2576
rect 8300 2592 8352 2644
rect 9864 2592 9916 2644
rect 10324 2592 10376 2644
rect 12348 2592 12400 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 2136 2499 2188 2508
rect 2136 2465 2145 2499
rect 2145 2465 2179 2499
rect 2179 2465 2188 2499
rect 2136 2456 2188 2465
rect 3608 2456 3660 2508
rect 3884 2499 3936 2508
rect 3884 2465 3893 2499
rect 3893 2465 3927 2499
rect 3927 2465 3936 2499
rect 3884 2456 3936 2465
rect 4436 2456 4488 2508
rect 2780 2320 2832 2372
rect 3056 2320 3108 2372
rect 3332 2320 3384 2372
rect 4988 2388 5040 2440
rect 5172 2388 5224 2440
rect 5632 2456 5684 2508
rect 6920 2524 6972 2576
rect 7288 2524 7340 2576
rect 7472 2524 7524 2576
rect 8760 2524 8812 2576
rect 9220 2524 9272 2576
rect 9588 2524 9640 2576
rect 7656 2456 7708 2508
rect 8668 2456 8720 2508
rect 7748 2388 7800 2440
rect 6552 2320 6604 2372
rect 9864 2456 9916 2508
rect 10600 2524 10652 2576
rect 11152 2524 11204 2576
rect 11520 2524 11572 2576
rect 10324 2499 10376 2508
rect 10324 2465 10333 2499
rect 10333 2465 10367 2499
rect 10367 2465 10376 2499
rect 10324 2456 10376 2465
rect 10508 2456 10560 2508
rect 3424 2252 3476 2304
rect 7932 2252 7984 2304
rect 10876 2388 10928 2440
rect 12992 2388 13044 2440
rect 9312 2320 9364 2372
rect 10968 2320 11020 2372
rect 9128 2252 9180 2304
rect 10692 2252 10744 2304
rect 10876 2252 10928 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 2852 2150 2904 2202
rect 2916 2150 2968 2202
rect 2980 2150 3032 2202
rect 3044 2150 3096 2202
rect 6594 2150 6646 2202
rect 6658 2150 6710 2202
rect 6722 2150 6774 2202
rect 6786 2150 6838 2202
rect 10335 2150 10387 2202
rect 10399 2150 10451 2202
rect 10463 2150 10515 2202
rect 10527 2150 10579 2202
rect 6368 2048 6420 2100
rect 2964 1980 3016 2032
rect 4068 1980 4120 2032
rect 5908 1980 5960 2032
rect 6460 1980 6512 2032
rect 6552 1980 6604 2032
rect 8944 1980 8996 2032
rect 10048 1980 10100 2032
rect 6000 1912 6052 1964
rect 6828 1912 6880 1964
rect 6184 1776 6236 1828
rect 9220 1708 9272 1760
rect 10416 1708 10468 1760
rect 4252 1300 4304 1352
rect 4620 1300 4672 1352
rect 4804 1368 4856 1420
rect 5540 1368 5592 1420
rect 7748 1368 7800 1420
rect 8852 1368 8904 1420
rect 5448 1300 5500 1352
rect 4896 1164 4948 1216
rect 6368 1164 6420 1216
rect 10784 892 10836 944
rect 11520 892 11572 944
<< metal2 >>
rect 754 14818 810 15618
rect 2226 14818 2282 15618
rect 3698 14818 3754 15618
rect 5170 14818 5226 15618
rect 6642 14818 6698 15618
rect 8206 14818 8262 15618
rect 9678 14818 9734 15618
rect 11150 14818 11206 15618
rect 12622 14818 12678 15618
rect 664 13456 716 13462
rect 664 13398 716 13404
rect 480 13388 532 13394
rect 480 13330 532 13336
rect 388 13184 440 13190
rect 388 13126 440 13132
rect 296 12844 348 12850
rect 296 12786 348 12792
rect 112 10532 164 10538
rect 112 10474 164 10480
rect 124 4146 152 10474
rect 204 4684 256 4690
rect 204 4626 256 4632
rect 112 4140 164 4146
rect 112 4082 164 4088
rect 112 4004 164 4010
rect 112 3946 164 3952
rect 20 3936 72 3942
rect 20 3878 72 3884
rect 32 800 60 3878
rect 124 800 152 3946
rect 216 800 244 4626
rect 308 2854 336 12786
rect 400 4146 428 13126
rect 388 4140 440 4146
rect 388 4082 440 4088
rect 388 3868 440 3874
rect 388 3810 440 3816
rect 296 2848 348 2854
rect 296 2790 348 2796
rect 400 800 428 3810
rect 492 3738 520 13330
rect 570 12472 626 12481
rect 570 12407 626 12416
rect 480 3732 532 3738
rect 480 3674 532 3680
rect 584 2774 612 12407
rect 676 4078 704 13398
rect 768 7313 796 14818
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 940 12708 992 12714
rect 940 12650 992 12656
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 754 7304 810 7313
rect 754 7239 810 7248
rect 664 4072 716 4078
rect 664 4014 716 4020
rect 754 4040 810 4049
rect 754 3975 810 3984
rect 662 2952 718 2961
rect 662 2887 718 2896
rect 492 2746 612 2774
rect 492 800 520 2746
rect 676 800 704 2887
rect 768 800 796 3975
rect 860 800 888 8366
rect 952 2961 980 12650
rect 1872 12646 1900 12718
rect 1860 12640 1912 12646
rect 1858 12608 1860 12617
rect 2044 12640 2096 12646
rect 1912 12608 1914 12617
rect 2044 12582 2096 12588
rect 1858 12543 1914 12552
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1306 12200 1362 12209
rect 1306 12135 1362 12144
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 938 2952 994 2961
rect 938 2887 994 2896
rect 1044 800 1072 9522
rect 1136 4214 1164 11834
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 1228 5030 1256 6734
rect 1216 5024 1268 5030
rect 1216 4966 1268 4972
rect 1124 4208 1176 4214
rect 1124 4150 1176 4156
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 1136 2961 1164 4014
rect 1228 3602 1256 4966
rect 1216 3596 1268 3602
rect 1216 3538 1268 3544
rect 1122 2952 1178 2961
rect 1122 2887 1178 2896
rect 1124 2644 1176 2650
rect 1124 2586 1176 2592
rect 1136 800 1164 2586
rect 1320 800 1348 12135
rect 1688 11354 1716 12242
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11830 1808 12038
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1964 11286 1992 11494
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10130 1532 10950
rect 1780 10810 1808 11154
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1412 9722 1440 10066
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9081 1440 9318
rect 1780 9178 1808 9998
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1584 9104 1636 9110
rect 1398 9072 1454 9081
rect 1584 9046 1636 9052
rect 1398 9007 1454 9016
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1490 8800 1546 8809
rect 1412 8634 1440 8774
rect 1490 8735 1546 8744
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 6458 1440 8434
rect 1504 8362 1532 8735
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5914 1440 6190
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1504 4282 1532 7278
rect 1596 6769 1624 9046
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8634 1716 8978
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 8537 1808 9114
rect 1766 8528 1822 8537
rect 1766 8463 1822 8472
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 8022 1716 8366
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1582 6760 1638 6769
rect 1582 6695 1638 6704
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 5642 1624 6598
rect 1688 6458 1716 6802
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5778 1716 6054
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 800 1440 4082
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1504 800 1532 3674
rect 1596 2990 1624 4422
rect 1688 4049 1716 4626
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1780 3233 1808 7278
rect 1872 6934 1900 10202
rect 1950 10024 2006 10033
rect 1950 9959 2006 9968
rect 1860 6928 1912 6934
rect 1860 6870 1912 6876
rect 1858 6760 1914 6769
rect 1858 6695 1914 6704
rect 1872 4486 1900 6695
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1964 4146 1992 9959
rect 2056 7886 2084 12582
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11762 2176 12038
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11218 2176 11698
rect 2240 11354 2268 14818
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2226 10704 2282 10713
rect 2136 10668 2188 10674
rect 2226 10639 2282 10648
rect 2136 10610 2188 10616
rect 2148 9586 2176 10610
rect 2240 10538 2268 10639
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 8548 2176 9522
rect 2332 9518 2360 13194
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2424 12646 2452 12718
rect 2412 12640 2464 12646
rect 2410 12608 2412 12617
rect 2596 12640 2648 12646
rect 2464 12608 2466 12617
rect 2596 12582 2648 12588
rect 2410 12543 2466 12552
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2424 11694 2452 12378
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 10674 2452 11630
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2516 10606 2544 11018
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10130 2452 10406
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 9178 2452 9318
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8673 2268 8978
rect 2424 8809 2452 9114
rect 2410 8800 2466 8809
rect 2410 8735 2466 8744
rect 2226 8664 2282 8673
rect 2226 8599 2282 8608
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2148 8520 2268 8548
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2240 8378 2268 8520
rect 2148 8072 2176 8366
rect 2240 8350 2360 8378
rect 2148 8044 2268 8072
rect 2134 7984 2190 7993
rect 2134 7919 2190 7928
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 6118 2084 7686
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5166 2084 5510
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2148 4978 2176 7919
rect 2056 4950 2176 4978
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1858 3632 1914 3641
rect 1858 3567 1914 3576
rect 1766 3224 1822 3233
rect 1766 3159 1822 3168
rect 1872 3040 1900 3567
rect 1964 3194 1992 3878
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1688 3012 1900 3040
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2514 1624 2926
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1688 800 1716 3012
rect 1858 2952 1914 2961
rect 1780 2910 1858 2938
rect 1780 800 1808 2910
rect 1858 2887 1914 2896
rect 1858 2816 1914 2825
rect 1858 2751 1914 2760
rect 1872 2394 1900 2751
rect 1964 2514 1992 3130
rect 2056 3058 2084 4950
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 2148 4282 2176 4490
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2148 2990 2176 4014
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1872 2366 1992 2394
rect 1964 800 1992 2366
rect 2056 800 2084 2790
rect 2148 2514 2176 2926
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2240 2394 2268 8044
rect 2332 7886 2360 8350
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2332 7449 2360 7822
rect 2318 7440 2374 7449
rect 2318 7375 2374 7384
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 6225 2360 7278
rect 2318 6216 2374 6225
rect 2318 6151 2374 6160
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 2990 2360 6054
rect 2424 5914 2452 8570
rect 2516 8312 2544 10542
rect 2608 10266 2636 12582
rect 2700 11121 2728 13466
rect 2826 13084 3122 13104
rect 2882 13082 2906 13084
rect 2962 13082 2986 13084
rect 3042 13082 3066 13084
rect 2904 13030 2906 13082
rect 2968 13030 2980 13082
rect 3042 13030 3044 13082
rect 2882 13028 2906 13030
rect 2962 13028 2986 13030
rect 3042 13028 3066 13030
rect 2826 13008 3122 13028
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3436 12434 3464 12854
rect 3436 12406 3556 12434
rect 2826 11996 3122 12016
rect 2882 11994 2906 11996
rect 2962 11994 2986 11996
rect 3042 11994 3066 11996
rect 2904 11942 2906 11994
rect 2968 11942 2980 11994
rect 3042 11942 3044 11994
rect 2882 11940 2906 11942
rect 2962 11940 2986 11942
rect 3042 11940 3066 11942
rect 2826 11920 3122 11940
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2792 11354 2820 11562
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 3344 11218 3372 11494
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2826 10908 3122 10928
rect 2882 10906 2906 10908
rect 2962 10906 2986 10908
rect 3042 10906 3066 10908
rect 2904 10854 2906 10906
rect 2968 10854 2980 10906
rect 3042 10854 3044 10906
rect 2882 10852 2906 10854
rect 2962 10852 2986 10854
rect 3042 10852 3066 10854
rect 2826 10832 3122 10852
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2688 10260 2740 10266
rect 2792 10248 2820 10678
rect 2884 10662 3096 10690
rect 2884 10606 2912 10662
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2872 10464 2924 10470
rect 2870 10432 2872 10441
rect 2924 10432 2926 10441
rect 2870 10367 2926 10376
rect 2792 10220 2912 10248
rect 2688 10202 2740 10208
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2608 9518 2636 9590
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2504 8306 2556 8312
rect 2504 8248 2556 8254
rect 2608 7834 2636 8842
rect 2700 8090 2728 10202
rect 2884 10130 2912 10220
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2976 9994 3004 10474
rect 3068 10010 3096 10662
rect 3344 10606 3372 11154
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3148 10464 3200 10470
rect 3252 10441 3280 10542
rect 3148 10406 3200 10412
rect 3238 10432 3294 10441
rect 3160 10198 3188 10406
rect 3238 10367 3294 10376
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3422 10160 3478 10169
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3332 10124 3384 10130
rect 3422 10095 3478 10104
rect 3332 10066 3384 10072
rect 2964 9988 3016 9994
rect 3068 9982 3188 10010
rect 2964 9930 3016 9936
rect 2826 9820 3122 9840
rect 2882 9818 2906 9820
rect 2962 9818 2986 9820
rect 3042 9818 3066 9820
rect 2904 9766 2906 9818
rect 2968 9766 2980 9818
rect 3042 9766 3044 9818
rect 2882 9764 2906 9766
rect 2962 9764 2986 9766
rect 3042 9764 3066 9766
rect 2826 9744 3122 9764
rect 2826 8732 3122 8752
rect 2882 8730 2906 8732
rect 2962 8730 2986 8732
rect 3042 8730 3066 8732
rect 2904 8678 2906 8730
rect 2968 8678 2980 8730
rect 3042 8678 3044 8730
rect 2882 8676 2906 8678
rect 2962 8676 2986 8678
rect 3042 8676 3066 8678
rect 2826 8656 3122 8676
rect 2872 8560 2924 8566
rect 2778 8528 2834 8537
rect 2872 8502 2924 8508
rect 2778 8463 2780 8472
rect 2832 8463 2834 8472
rect 2780 8434 2832 8440
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2884 7954 2912 8502
rect 2962 8392 3018 8401
rect 2962 8327 2964 8336
rect 3016 8327 3018 8336
rect 3056 8356 3108 8362
rect 2964 8298 3016 8304
rect 3056 8298 3108 8304
rect 3068 8090 3096 8298
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2516 7806 2636 7834
rect 2516 6100 2544 7806
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7206 2636 7686
rect 2700 7546 2728 7890
rect 2826 7644 3122 7664
rect 2882 7642 2906 7644
rect 2962 7642 2986 7644
rect 3042 7642 3066 7644
rect 2904 7590 2906 7642
rect 2968 7590 2980 7642
rect 3042 7590 3044 7642
rect 2882 7588 2906 7590
rect 2962 7588 2986 7590
rect 3042 7588 3066 7590
rect 2826 7568 3122 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2964 7472 3016 7478
rect 2778 7440 2834 7449
rect 2688 7404 2740 7410
rect 3056 7472 3108 7478
rect 2964 7414 3016 7420
rect 3054 7440 3056 7449
rect 3108 7440 3110 7449
rect 2778 7375 2834 7384
rect 2688 7346 2740 7352
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2700 7041 2728 7346
rect 2686 7032 2742 7041
rect 2686 6967 2742 6976
rect 2688 6860 2740 6866
rect 2792 6848 2820 7375
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2884 7002 2912 7278
rect 2976 7041 3004 7414
rect 3054 7375 3110 7384
rect 2962 7032 3018 7041
rect 2872 6996 2924 7002
rect 2962 6967 3018 6976
rect 2872 6938 2924 6944
rect 2740 6820 2820 6848
rect 2688 6802 2740 6808
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2608 6254 2636 6666
rect 2700 6322 2728 6802
rect 2826 6556 3122 6576
rect 2882 6554 2906 6556
rect 2962 6554 2986 6556
rect 3042 6554 3066 6556
rect 2904 6502 2906 6554
rect 2968 6502 2980 6554
rect 3042 6502 3044 6554
rect 2882 6500 2906 6502
rect 2962 6500 2986 6502
rect 3042 6500 3066 6502
rect 2826 6480 3122 6500
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2516 6072 2636 6100
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5234 2452 5510
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2424 4826 2452 5034
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2318 2816 2374 2825
rect 2318 2751 2374 2760
rect 2148 2366 2268 2394
rect 2148 800 2176 2366
rect 2332 800 2360 2751
rect 2424 800 2452 4422
rect 2516 4282 2544 5782
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3126 2544 4082
rect 2608 4078 2636 6072
rect 2700 5778 2728 6258
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2976 5681 3004 6190
rect 3068 5710 3096 6326
rect 3160 5914 3188 9982
rect 3252 8945 3280 10066
rect 3238 8936 3294 8945
rect 3238 8871 3294 8880
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3252 7954 3280 8570
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 7478 3280 7754
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3252 6390 3280 7414
rect 3344 6905 3372 10066
rect 3436 8974 3464 10095
rect 3528 10010 3556 12406
rect 3712 12374 3740 14818
rect 5184 12986 5212 14818
rect 6656 13240 6684 14818
rect 8220 13682 8248 14818
rect 8220 13654 8432 13682
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7932 13252 7984 13258
rect 6656 13212 6960 13240
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4172 12481 4200 12582
rect 4158 12472 4214 12481
rect 4158 12407 4214 12416
rect 4264 12374 4292 12582
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11694 3832 12038
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3620 10198 3648 11154
rect 3804 10674 3832 11630
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3712 10130 3740 10474
rect 3804 10169 3832 10610
rect 3790 10160 3846 10169
rect 3700 10124 3752 10130
rect 3790 10095 3846 10104
rect 3700 10066 3752 10072
rect 3528 9982 3832 10010
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 9489 3556 9522
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7954 3464 8230
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3436 7546 3464 7890
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3330 6896 3386 6905
rect 3330 6831 3386 6840
rect 3330 6760 3386 6769
rect 3330 6695 3386 6704
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5953 3280 6190
rect 3238 5944 3294 5953
rect 3148 5908 3200 5914
rect 3238 5879 3294 5888
rect 3148 5850 3200 5856
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3056 5704 3108 5710
rect 2962 5672 3018 5681
rect 2688 5636 2740 5642
rect 3056 5646 3108 5652
rect 2962 5607 3018 5616
rect 2688 5578 2740 5584
rect 2700 5370 2728 5578
rect 2826 5468 3122 5488
rect 2882 5466 2906 5468
rect 2962 5466 2986 5468
rect 3042 5466 3066 5468
rect 2904 5414 2906 5466
rect 2968 5414 2980 5466
rect 3042 5414 3044 5466
rect 2882 5412 2906 5414
rect 2962 5412 2986 5414
rect 3042 5412 3066 5414
rect 2826 5392 3122 5412
rect 3160 5370 3188 5714
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2700 4690 2728 5306
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2792 4468 2820 5170
rect 3252 5166 3280 5510
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 2700 4440 2820 4468
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2516 1986 2544 2926
rect 2608 2774 2636 3606
rect 2700 2836 2728 4440
rect 2826 4380 3122 4400
rect 2882 4378 2906 4380
rect 2962 4378 2986 4380
rect 3042 4378 3066 4380
rect 2904 4326 2906 4378
rect 2968 4326 2980 4378
rect 3042 4326 3044 4378
rect 2882 4324 2906 4326
rect 2962 4324 2986 4326
rect 3042 4324 3066 4326
rect 2826 4304 3122 4324
rect 3160 4214 3188 4490
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 3148 4208 3200 4214
rect 3344 4162 3372 6695
rect 3436 6458 3464 7278
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5030 3464 6258
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4758 3464 4966
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3148 4150 3200 4156
rect 2884 3466 2912 4150
rect 3252 4134 3372 4162
rect 3436 4146 3464 4694
rect 3424 4140 3476 4146
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3068 3738 3096 4014
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3160 3534 3188 3878
rect 3252 3738 3280 4134
rect 3424 4082 3476 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3344 3913 3372 4014
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3240 3732 3292 3738
rect 3528 3720 3556 8774
rect 3620 6338 3648 9862
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3712 7449 3740 9658
rect 3698 7440 3754 7449
rect 3698 7375 3754 7384
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 6866 3740 7142
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3712 6497 3740 6666
rect 3698 6488 3754 6497
rect 3698 6423 3754 6432
rect 3620 6310 3740 6338
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5914 3648 6190
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3620 4593 3648 4626
rect 3606 4584 3662 4593
rect 3606 4519 3662 4528
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4146 3648 4422
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3240 3674 3292 3680
rect 3344 3692 3556 3720
rect 3608 3732 3660 3738
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2826 3292 3122 3312
rect 2882 3290 2906 3292
rect 2962 3290 2986 3292
rect 3042 3290 3066 3292
rect 2904 3238 2906 3290
rect 2968 3238 2980 3290
rect 3042 3238 3044 3290
rect 2882 3236 2906 3238
rect 2962 3236 2986 3238
rect 3042 3236 3066 3238
rect 2826 3216 3122 3236
rect 3252 3194 3280 3538
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 3238 3088 3294 3097
rect 2700 2808 2820 2836
rect 2608 2746 2728 2774
rect 2700 2088 2728 2746
rect 2792 2378 2820 2808
rect 2884 2774 2912 3062
rect 3238 3023 3294 3032
rect 3146 2952 3202 2961
rect 3146 2887 3202 2896
rect 2884 2746 3096 2774
rect 2872 2576 2924 2582
rect 2870 2544 2872 2553
rect 2924 2544 2926 2553
rect 2870 2479 2926 2488
rect 3068 2378 3096 2746
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 2826 2204 3122 2224
rect 2882 2202 2906 2204
rect 2962 2202 2986 2204
rect 3042 2202 3066 2204
rect 2904 2150 2906 2202
rect 2968 2150 2980 2202
rect 3042 2150 3044 2202
rect 2882 2148 2906 2150
rect 2962 2148 2986 2150
rect 3042 2148 3066 2150
rect 2826 2128 3122 2148
rect 2700 2060 2820 2088
rect 2516 1958 2728 1986
rect 2594 1864 2650 1873
rect 2594 1799 2650 1808
rect 2608 800 2636 1799
rect 2700 800 2728 1958
rect 2792 800 2820 2060
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 2976 800 3004 1974
rect 3160 898 3188 2887
rect 3068 870 3188 898
rect 3068 800 3096 870
rect 3252 800 3280 3023
rect 3344 2650 3372 3692
rect 3608 3674 3660 3680
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2582 3464 3538
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2990 3556 3334
rect 3620 3074 3648 3674
rect 3712 3194 3740 6310
rect 3804 5846 3832 9982
rect 3896 9654 3924 10950
rect 3988 10470 4016 11494
rect 4356 11370 4384 12854
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11694 4476 12242
rect 4540 11762 4568 12786
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4632 11898 4660 12718
rect 4697 12540 4993 12560
rect 4753 12538 4777 12540
rect 4833 12538 4857 12540
rect 4913 12538 4937 12540
rect 4775 12486 4777 12538
rect 4839 12486 4851 12538
rect 4913 12486 4915 12538
rect 4753 12484 4777 12486
rect 4833 12484 4857 12486
rect 4913 12484 4937 12486
rect 4697 12464 4993 12484
rect 5184 12374 5212 12718
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 5000 11642 5028 12038
rect 5078 11928 5134 11937
rect 5078 11863 5080 11872
rect 5132 11863 5134 11872
rect 5172 11892 5224 11898
rect 5080 11834 5132 11840
rect 5172 11834 5224 11840
rect 5184 11778 5212 11834
rect 5092 11762 5212 11778
rect 5080 11756 5212 11762
rect 5132 11750 5212 11756
rect 5080 11698 5132 11704
rect 5000 11614 5212 11642
rect 5078 11520 5134 11529
rect 4697 11452 4993 11472
rect 5078 11455 5134 11464
rect 4753 11450 4777 11452
rect 4833 11450 4857 11452
rect 4913 11450 4937 11452
rect 4775 11398 4777 11450
rect 4839 11398 4851 11450
rect 4913 11398 4915 11450
rect 4753 11396 4777 11398
rect 4833 11396 4857 11398
rect 4913 11396 4937 11398
rect 4697 11376 4993 11396
rect 4356 11342 4660 11370
rect 5092 11354 5120 11455
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4080 10010 4108 11154
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10266 4200 11086
rect 4264 10606 4292 11222
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4250 10432 4306 10441
rect 4250 10367 4306 10376
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3988 9982 4108 10010
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3896 9110 3924 9590
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3896 8537 3924 8910
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3896 8090 3924 8463
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7585 4016 9982
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3974 7576 4030 7585
rect 3974 7511 4030 7520
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3896 6798 3924 6938
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3884 6656 3936 6662
rect 3988 6633 4016 7346
rect 3884 6598 3936 6604
rect 3974 6624 4030 6633
rect 3896 6254 3924 6598
rect 3974 6559 4030 6568
rect 3974 6488 4030 6497
rect 3974 6423 4030 6432
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3988 5896 4016 6423
rect 4080 6089 4108 9862
rect 4066 6080 4122 6089
rect 4066 6015 4122 6024
rect 3896 5868 4016 5896
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3896 5098 3924 5868
rect 4172 5794 4200 10066
rect 4264 9353 4292 10367
rect 4250 9344 4306 9353
rect 4250 9279 4306 9288
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4264 8362 4292 9114
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 8022 4292 8298
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4264 6934 4292 7414
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4250 6624 4306 6633
rect 4250 6559 4306 6568
rect 4264 6458 4292 6559
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 5794 4384 11154
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4448 10538 4476 10639
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4434 10432 4490 10441
rect 4434 10367 4490 10376
rect 4448 10198 4476 10367
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9761 4476 9862
rect 4434 9752 4490 9761
rect 4434 9687 4490 9696
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 9110 4476 9318
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7954 4476 8230
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4448 7585 4476 7754
rect 4434 7576 4490 7585
rect 4434 7511 4490 7520
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 3988 5766 4200 5794
rect 4264 5766 4384 5794
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 3942 3832 4626
rect 3896 4554 3924 5034
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3882 3904 3938 3913
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3620 3046 3740 3074
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3620 2514 3648 2926
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3712 2394 3740 3046
rect 3804 2904 3832 3878
rect 3882 3839 3938 3848
rect 3896 3738 3924 3839
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3896 3194 3924 3538
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3884 2916 3936 2922
rect 3804 2876 3884 2904
rect 3884 2858 3936 2864
rect 3882 2816 3938 2825
rect 3882 2751 3938 2760
rect 3988 2774 4016 5766
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 4826 4200 5646
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4080 2922 4108 4247
rect 4172 3738 4200 4626
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3482 4292 5766
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 5370 4384 5646
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4356 4690 4384 5306
rect 4448 5234 4476 7210
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4448 4593 4476 5034
rect 4434 4584 4490 4593
rect 4344 4548 4396 4554
rect 4434 4519 4490 4528
rect 4344 4490 4396 4496
rect 4356 4078 4384 4490
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3777 4384 4014
rect 4342 3768 4398 3777
rect 4342 3703 4398 3712
rect 4540 3618 4568 11154
rect 4632 10810 4660 11342
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4712 10600 4764 10606
rect 4816 10577 4844 10950
rect 4908 10713 4936 10950
rect 4894 10704 4950 10713
rect 4894 10639 4950 10648
rect 4712 10542 4764 10548
rect 4802 10568 4858 10577
rect 4724 10452 4752 10542
rect 4802 10503 4858 10512
rect 4632 10424 4752 10452
rect 4632 10248 4660 10424
rect 4697 10364 4993 10384
rect 4753 10362 4777 10364
rect 4833 10362 4857 10364
rect 4913 10362 4937 10364
rect 4775 10310 4777 10362
rect 4839 10310 4851 10362
rect 4913 10310 4915 10362
rect 4753 10308 4777 10310
rect 4833 10308 4857 10310
rect 4913 10308 4937 10310
rect 4697 10288 4993 10308
rect 4632 10220 4752 10248
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4632 9654 4660 10066
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4620 9512 4672 9518
rect 4618 9480 4620 9489
rect 4672 9480 4674 9489
rect 4618 9415 4674 9424
rect 4724 9364 4752 10220
rect 4896 10124 4948 10130
rect 4816 10084 4896 10112
rect 4816 9722 4844 10084
rect 4896 10066 4948 10072
rect 4986 10024 5042 10033
rect 4986 9959 4988 9968
rect 5040 9959 5042 9968
rect 4988 9930 5040 9936
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4896 9648 4948 9654
rect 4894 9616 4896 9625
rect 4948 9616 4950 9625
rect 4894 9551 4950 9560
rect 4632 9336 4752 9364
rect 4632 7478 4660 9336
rect 4697 9276 4993 9296
rect 4753 9274 4777 9276
rect 4833 9274 4857 9276
rect 4913 9274 4937 9276
rect 4775 9222 4777 9274
rect 4839 9222 4851 9274
rect 4913 9222 4915 9274
rect 4753 9220 4777 9222
rect 4833 9220 4857 9222
rect 4913 9220 4937 9222
rect 4697 9200 4993 9220
rect 5092 9058 5120 11154
rect 4908 9030 5120 9058
rect 4908 8276 4936 9030
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5000 8498 5028 8910
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8401 5120 8434
rect 5184 8430 5212 11614
rect 5276 11354 5304 12786
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 11830 5396 12582
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5460 11370 5488 12786
rect 6196 12782 6224 13126
rect 6568 13084 6864 13104
rect 6624 13082 6648 13084
rect 6704 13082 6728 13084
rect 6784 13082 6808 13084
rect 6646 13030 6648 13082
rect 6710 13030 6722 13082
rect 6784 13030 6786 13082
rect 6624 13028 6648 13030
rect 6704 13028 6728 13030
rect 6784 13028 6808 13030
rect 6568 13008 6864 13028
rect 6932 12986 6960 13212
rect 7932 13194 7984 13200
rect 7944 12986 7972 13194
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8128 12782 8156 13330
rect 8404 12986 8432 13654
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 5552 12209 5580 12718
rect 5644 12442 5672 12718
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5368 11342 5488 11370
rect 5368 10849 5396 11342
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5354 10840 5410 10849
rect 5354 10775 5410 10784
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5172 8424 5224 8430
rect 5078 8392 5134 8401
rect 5172 8366 5224 8372
rect 5078 8327 5134 8336
rect 5172 8288 5224 8294
rect 4908 8248 5120 8276
rect 4697 8188 4993 8208
rect 4753 8186 4777 8188
rect 4833 8186 4857 8188
rect 4913 8186 4937 8188
rect 4775 8134 4777 8186
rect 4839 8134 4851 8186
rect 4913 8134 4915 8186
rect 4753 8132 4777 8134
rect 4833 8132 4857 8134
rect 4913 8132 4937 8134
rect 4697 8112 4993 8132
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7546 4844 7890
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4986 7440 5042 7449
rect 4986 7375 5042 7384
rect 5000 7342 5028 7375
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4632 6497 4660 7278
rect 4697 7100 4993 7120
rect 4753 7098 4777 7100
rect 4833 7098 4857 7100
rect 4913 7098 4937 7100
rect 4775 7046 4777 7098
rect 4839 7046 4851 7098
rect 4913 7046 4915 7098
rect 4753 7044 4777 7046
rect 4833 7044 4857 7046
rect 4913 7044 4937 7046
rect 4697 7024 4993 7044
rect 5092 6769 5120 8248
rect 5172 8230 5224 8236
rect 5078 6760 5134 6769
rect 5078 6695 5134 6704
rect 4618 6488 4674 6497
rect 4618 6423 4674 6432
rect 5078 6352 5134 6361
rect 5078 6287 5080 6296
rect 5132 6287 5134 6296
rect 5080 6258 5132 6264
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4632 4570 4660 6190
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4697 6012 4993 6032
rect 4753 6010 4777 6012
rect 4833 6010 4857 6012
rect 4913 6010 4937 6012
rect 4775 5958 4777 6010
rect 4839 5958 4851 6010
rect 4913 5958 4915 6010
rect 4753 5956 4777 5958
rect 4833 5956 4857 5958
rect 4913 5956 4937 5958
rect 4697 5936 4993 5956
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5000 5098 5028 5714
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4697 4924 4993 4944
rect 4753 4922 4777 4924
rect 4833 4922 4857 4924
rect 4913 4922 4937 4924
rect 4775 4870 4777 4922
rect 4839 4870 4851 4922
rect 4913 4870 4915 4922
rect 4753 4868 4777 4870
rect 4833 4868 4857 4870
rect 4913 4868 4937 4870
rect 4697 4848 4993 4868
rect 4632 4542 4752 4570
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4282 4660 4422
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4172 3454 4292 3482
rect 4356 3590 4568 3618
rect 4172 2961 4200 3454
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 3058 4292 3334
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4158 2952 4214 2961
rect 4068 2916 4120 2922
rect 4158 2887 4214 2896
rect 4068 2858 4120 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3790 2680 3846 2689
rect 3790 2615 3846 2624
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3620 2366 3740 2394
rect 3344 800 3372 2314
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 800 3464 2246
rect 3620 800 3648 2366
rect 3804 1034 3832 2615
rect 3896 2514 3924 2751
rect 3988 2746 4108 2774
rect 3974 2680 4030 2689
rect 3974 2615 4030 2624
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3988 1442 4016 2615
rect 4080 2038 4108 2746
rect 4172 2582 4200 2790
rect 4356 2774 4384 3590
rect 4632 3534 4660 4218
rect 4724 4010 4752 4542
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4697 3836 4993 3856
rect 4753 3834 4777 3836
rect 4833 3834 4857 3836
rect 4913 3834 4937 3836
rect 4775 3782 4777 3834
rect 4839 3782 4851 3834
rect 4913 3782 4915 3834
rect 4753 3780 4777 3782
rect 4833 3780 4857 3782
rect 4913 3780 4937 3782
rect 4697 3760 4993 3780
rect 4802 3632 4858 3641
rect 4802 3567 4858 3576
rect 4436 3528 4488 3534
rect 4620 3528 4672 3534
rect 4436 3470 4488 3476
rect 4526 3496 4582 3505
rect 4264 2746 4384 2774
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4264 1442 4292 2746
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 3712 1006 3832 1034
rect 3896 1414 4016 1442
rect 4080 1414 4292 1442
rect 3712 800 3740 1006
rect 3896 800 3924 1414
rect 4080 1306 4108 1414
rect 3988 1278 4108 1306
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 3988 800 4016 1278
rect 4066 1184 4122 1193
rect 4066 1119 4122 1128
rect 4080 800 4108 1119
rect 4264 800 4292 1294
rect 4356 800 4384 2518
rect 4448 2514 4476 3470
rect 4620 3470 4672 3476
rect 4526 3431 4582 3440
rect 4540 2904 4568 3431
rect 4632 3126 4660 3470
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4816 3058 4844 3567
rect 5092 3482 5120 6122
rect 5184 6066 5212 8230
rect 5276 6186 5304 10678
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 8514 5396 10610
rect 5460 10588 5488 11154
rect 5552 10810 5580 11698
rect 5644 11626 5672 12378
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5920 11937 5948 12242
rect 6380 12170 6408 12378
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6568 11996 6864 12016
rect 6624 11994 6648 11996
rect 6704 11994 6728 11996
rect 6784 11994 6808 11996
rect 6646 11942 6648 11994
rect 6710 11942 6722 11994
rect 6784 11942 6786 11994
rect 6624 11940 6648 11942
rect 6704 11940 6728 11942
rect 6784 11940 6808 11942
rect 5906 11928 5962 11937
rect 5816 11892 5868 11898
rect 6568 11920 6864 11940
rect 6932 11898 6960 12242
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11898 7052 12038
rect 5906 11863 5962 11872
rect 6920 11892 6972 11898
rect 5816 11834 5868 11840
rect 6920 11834 6972 11840
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5630 11384 5686 11393
rect 5630 11319 5632 11328
rect 5684 11319 5686 11328
rect 5632 11290 5684 11296
rect 5630 11248 5686 11257
rect 5630 11183 5632 11192
rect 5684 11183 5686 11192
rect 5632 11154 5684 11160
rect 5736 11121 5764 11630
rect 5722 11112 5778 11121
rect 5632 11076 5684 11082
rect 5828 11082 5856 11834
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5722 11047 5778 11056
rect 5816 11076 5868 11082
rect 5632 11018 5684 11024
rect 5816 11018 5868 11024
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10600 5592 10606
rect 5460 10560 5540 10588
rect 5460 9518 5488 10560
rect 5540 10542 5592 10548
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5552 9926 5580 10134
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5552 9450 5580 9862
rect 5644 9625 5672 11018
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5630 9616 5686 9625
rect 5630 9551 5686 9560
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5446 9344 5502 9353
rect 5446 9279 5502 9288
rect 5460 9178 5488 9279
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5552 8634 5580 9386
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 9110 5672 9318
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5368 8486 5488 8514
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 8090 5396 8366
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5354 7848 5410 7857
rect 5354 7783 5410 7792
rect 5368 6390 5396 7783
rect 5460 7750 5488 8486
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5552 7546 5580 8366
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8022 5672 8230
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5736 7426 5764 10950
rect 5828 10810 5856 11018
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5814 10024 5870 10033
rect 5814 9959 5870 9968
rect 5828 7954 5856 9959
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5460 7398 5764 7426
rect 5460 6769 5488 7398
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5446 6760 5502 6769
rect 5446 6695 5502 6704
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5460 6322 5488 6559
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5184 6038 5304 6066
rect 5170 5944 5226 5953
rect 5170 5879 5172 5888
rect 5224 5879 5226 5888
rect 5172 5850 5224 5856
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5184 3913 5212 5646
rect 5276 5302 5304 6038
rect 5460 5846 5488 6258
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5276 4826 5304 5238
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5170 3904 5226 3913
rect 5170 3839 5226 3848
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5000 3454 5120 3482
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4816 2961 4844 2994
rect 4802 2952 4858 2961
rect 4540 2876 4660 2904
rect 4908 2922 4936 3334
rect 4802 2887 4858 2896
rect 4896 2916 4948 2922
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4632 1358 4660 2876
rect 4896 2858 4948 2864
rect 5000 2836 5028 3454
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 2990 5120 3334
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5000 2808 5120 2836
rect 4697 2748 4993 2768
rect 4753 2746 4777 2748
rect 4833 2746 4857 2748
rect 4913 2746 4937 2748
rect 4775 2694 4777 2746
rect 4839 2694 4851 2746
rect 4913 2694 4915 2746
rect 4753 2692 4777 2694
rect 4833 2692 4857 2694
rect 4913 2692 4937 2694
rect 4697 2672 4993 2692
rect 5092 2632 5120 2808
rect 5184 2650 5212 3538
rect 5276 3233 5304 4626
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 5000 2604 5120 2632
rect 5172 2644 5224 2650
rect 4710 2544 4766 2553
rect 4710 2479 4766 2488
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 4526 1184 4582 1193
rect 4724 1170 4752 2479
rect 5000 2446 5028 2604
rect 5172 2586 5224 2592
rect 5368 2530 5396 5714
rect 5446 5128 5502 5137
rect 5446 5063 5502 5072
rect 5460 4282 5488 5063
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3194 5488 3538
rect 5552 3233 5580 7278
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 6866 5672 7142
rect 5736 7002 5764 7278
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5722 6760 5778 6769
rect 5722 6695 5778 6704
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5137 5672 5578
rect 5630 5128 5686 5137
rect 5630 5063 5686 5072
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 3738 5672 4966
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5644 3641 5672 3674
rect 5630 3632 5686 3641
rect 5630 3567 5632 3576
rect 5684 3567 5686 3576
rect 5632 3538 5684 3544
rect 5644 3507 5672 3538
rect 5538 3224 5594 3233
rect 5448 3188 5500 3194
rect 5538 3159 5594 3168
rect 5448 3130 5500 3136
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 2582 5488 2926
rect 5092 2502 5396 2530
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5092 2292 5120 2502
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5000 2264 5120 2292
rect 4804 1420 4856 1426
rect 4804 1362 4856 1368
rect 4526 1119 4582 1128
rect 4632 1142 4752 1170
rect 4540 800 4568 1119
rect 4632 800 4660 1142
rect 4816 1034 4844 1362
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 4724 1006 4844 1034
rect 4724 800 4752 1006
rect 4908 800 4936 1158
rect 5000 800 5028 2264
rect 5184 800 5212 2382
rect 5262 1592 5318 1601
rect 5262 1527 5318 1536
rect 5276 800 5304 1527
rect 5552 1426 5580 3023
rect 5632 2984 5684 2990
rect 5736 2972 5764 6695
rect 5828 6458 5856 7210
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5920 5778 5948 11494
rect 6012 11150 6040 11630
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6012 10606 6040 10950
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 6012 9897 6040 10134
rect 5998 9888 6054 9897
rect 5998 9823 6054 9832
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 6012 5534 6040 9318
rect 6104 9178 6132 11494
rect 6182 11112 6238 11121
rect 6182 11047 6238 11056
rect 6196 10810 6224 11047
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 9722 6224 10066
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6184 9512 6236 9518
rect 6182 9480 6184 9489
rect 6236 9480 6238 9489
rect 6182 9415 6238 9424
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8401 6132 8910
rect 6196 8566 6224 9415
rect 6288 8922 6316 11630
rect 6380 10810 6408 11698
rect 6458 11384 6514 11393
rect 7116 11354 7144 12650
rect 7208 12102 7236 12718
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8024 12640 8076 12646
rect 7944 12600 8024 12628
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11694 7236 12038
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7300 11626 7328 12310
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6458 11319 6514 11328
rect 7104 11348 7156 11354
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6472 10010 6500 11319
rect 7104 11290 7156 11296
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6564 11121 6592 11222
rect 7300 11218 7328 11562
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 6550 11112 6606 11121
rect 6550 11047 6606 11056
rect 6568 10908 6864 10928
rect 6624 10906 6648 10908
rect 6704 10906 6728 10908
rect 6784 10906 6808 10908
rect 6646 10854 6648 10906
rect 6710 10854 6722 10906
rect 6784 10854 6786 10906
rect 6624 10852 6648 10854
rect 6704 10852 6728 10854
rect 6784 10852 6808 10854
rect 6568 10832 6864 10852
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6552 10600 6604 10606
rect 6604 10560 6684 10588
rect 6552 10542 6604 10548
rect 6550 10296 6606 10305
rect 6550 10231 6606 10240
rect 6380 9982 6500 10010
rect 6380 9382 6408 9982
rect 6564 9908 6592 10231
rect 6656 10033 6684 10560
rect 6840 10470 6868 10678
rect 7300 10674 7328 11154
rect 7392 11121 7420 11630
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7378 11112 7434 11121
rect 7378 11047 7434 11056
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6932 10033 6960 10542
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6472 9880 6592 9908
rect 6920 9920 6972 9926
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6288 8894 6408 8922
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6090 8392 6146 8401
rect 6090 8327 6146 8336
rect 6196 8022 6224 8502
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 6186 6132 7686
rect 6196 7342 6224 7958
rect 6288 7954 6316 8774
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6380 7698 6408 8894
rect 6472 8616 6500 9880
rect 6920 9862 6972 9868
rect 6568 9820 6864 9840
rect 6624 9818 6648 9820
rect 6704 9818 6728 9820
rect 6784 9818 6808 9820
rect 6646 9766 6648 9818
rect 6710 9766 6722 9818
rect 6784 9766 6786 9818
rect 6624 9764 6648 9766
rect 6704 9764 6728 9766
rect 6784 9764 6808 9766
rect 6568 9744 6864 9764
rect 6932 9674 6960 9862
rect 7024 9722 7052 10066
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 6748 9646 6960 9674
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6748 9586 6776 9646
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9178 6776 9522
rect 6828 9512 6880 9518
rect 7208 9489 7236 9862
rect 7300 9722 7328 10610
rect 7576 10418 7604 11494
rect 7668 11121 7696 11630
rect 7654 11112 7710 11121
rect 7654 11047 7710 11056
rect 7576 10390 7696 10418
rect 7380 10260 7432 10266
rect 7432 10220 7604 10248
rect 7380 10202 7432 10208
rect 7470 10160 7526 10169
rect 7470 10095 7526 10104
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 6828 9454 6880 9460
rect 7194 9480 7250 9489
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 8906 6868 9454
rect 7194 9415 7250 9424
rect 7024 9042 7144 9058
rect 7208 9042 7236 9415
rect 7012 9036 7144 9042
rect 7064 9030 7144 9036
rect 7012 8978 7064 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6568 8732 6864 8752
rect 6624 8730 6648 8732
rect 6704 8730 6728 8732
rect 6784 8730 6808 8732
rect 6646 8678 6648 8730
rect 6710 8678 6722 8730
rect 6784 8678 6786 8730
rect 6624 8676 6648 8678
rect 6704 8676 6728 8678
rect 6784 8676 6808 8678
rect 6568 8656 6864 8676
rect 6472 8588 6592 8616
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 7886 6500 8434
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6564 7732 6592 8588
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 8090 6684 8366
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6748 7868 6776 8502
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6840 8022 6868 8298
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6748 7840 6960 7868
rect 6288 7670 6408 7698
rect 6472 7704 6592 7732
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6196 5846 6224 6938
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 5684 2944 5764 2972
rect 5828 5506 6040 5534
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5632 2926 5684 2932
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2514 5672 2790
rect 5722 2680 5778 2689
rect 5722 2615 5724 2624
rect 5776 2615 5778 2624
rect 5724 2586 5776 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5630 2408 5686 2417
rect 5630 2343 5686 2352
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5538 1320 5594 1329
rect 5460 898 5488 1294
rect 5538 1255 5594 1264
rect 5368 870 5488 898
rect 5368 800 5396 870
rect 5552 800 5580 1255
rect 5644 800 5672 2343
rect 5828 800 5856 5506
rect 5998 5400 6054 5409
rect 6104 5370 6132 5510
rect 5998 5335 6054 5344
rect 6092 5364 6144 5370
rect 5906 4856 5962 4865
rect 5906 4791 5962 4800
rect 5920 4282 5948 4791
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6012 4185 6040 5335
rect 6092 5306 6144 5312
rect 6196 5302 6224 5646
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6288 4808 6316 7670
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6380 6458 6408 7482
rect 6472 7392 6500 7704
rect 6568 7644 6864 7664
rect 6624 7642 6648 7644
rect 6704 7642 6728 7644
rect 6784 7642 6808 7644
rect 6646 7590 6648 7642
rect 6710 7590 6722 7642
rect 6784 7590 6786 7642
rect 6624 7588 6648 7590
rect 6704 7588 6728 7590
rect 6784 7588 6808 7590
rect 6568 7568 6864 7588
rect 6472 7364 6592 7392
rect 6458 7304 6514 7313
rect 6458 7239 6460 7248
rect 6512 7239 6514 7248
rect 6460 7210 6512 7216
rect 6564 6644 6592 7364
rect 6932 7206 6960 7840
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6472 6616 6592 6644
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6196 4780 6316 4808
rect 6196 4729 6224 4780
rect 6380 4729 6408 6190
rect 6472 5166 6500 6616
rect 6568 6556 6864 6576
rect 6624 6554 6648 6556
rect 6704 6554 6728 6556
rect 6784 6554 6808 6556
rect 6646 6502 6648 6554
rect 6710 6502 6722 6554
rect 6784 6502 6786 6554
rect 6624 6500 6648 6502
rect 6704 6500 6728 6502
rect 6784 6500 6808 6502
rect 6568 6480 6864 6500
rect 6932 6440 6960 6802
rect 6564 6412 6960 6440
rect 6564 5778 6592 6412
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 5914 6684 6190
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6748 5846 6776 6054
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6568 5468 6864 5488
rect 6624 5466 6648 5468
rect 6704 5466 6728 5468
rect 6784 5466 6808 5468
rect 6646 5414 6648 5466
rect 6710 5414 6722 5466
rect 6784 5414 6786 5466
rect 6624 5412 6648 5414
rect 6704 5412 6728 5414
rect 6784 5412 6808 5414
rect 6568 5392 6864 5412
rect 6932 5302 6960 6258
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6182 4720 6238 4729
rect 6182 4655 6238 4664
rect 6366 4720 6422 4729
rect 6932 4690 6960 4966
rect 6366 4655 6422 4664
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6274 4584 6330 4593
rect 6090 4448 6146 4457
rect 6090 4383 6146 4392
rect 5998 4176 6054 4185
rect 5998 4111 6054 4120
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5920 2038 5948 3946
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5908 2032 5960 2038
rect 5908 1974 5960 1980
rect 6012 1970 6040 3839
rect 6104 2258 6132 4383
rect 6196 4282 6224 4558
rect 6918 4584 6974 4593
rect 6274 4519 6330 4528
rect 6460 4548 6512 4554
rect 6288 4282 6316 4519
rect 6918 4519 6974 4528
rect 6460 4490 6512 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3505 6224 3878
rect 6288 3777 6316 4014
rect 6380 3890 6408 4422
rect 6472 4078 6500 4490
rect 6932 4486 6960 4519
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6568 4380 6864 4400
rect 6624 4378 6648 4380
rect 6704 4378 6728 4380
rect 6784 4378 6808 4380
rect 6646 4326 6648 4378
rect 6710 4326 6722 4378
rect 6784 4326 6786 4378
rect 6624 4324 6648 4326
rect 6704 4324 6728 4326
rect 6784 4324 6808 4326
rect 6568 4304 6864 4324
rect 6932 4282 6960 4422
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6460 4072 6512 4078
rect 6644 4072 6696 4078
rect 6460 4014 6512 4020
rect 6564 4020 6644 4026
rect 6564 4014 6696 4020
rect 6564 3998 6684 4014
rect 6920 4004 6972 4010
rect 6564 3890 6592 3998
rect 6920 3946 6972 3952
rect 6932 3913 6960 3946
rect 6380 3862 6592 3890
rect 6918 3904 6974 3913
rect 6274 3768 6330 3777
rect 6274 3703 6330 3712
rect 6380 3618 6408 3862
rect 6918 3839 6974 3848
rect 6932 3641 6960 3839
rect 6288 3590 6408 3618
rect 6918 3632 6974 3641
rect 6460 3596 6512 3602
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6196 2990 6224 3334
rect 6288 3058 6316 3590
rect 6918 3567 6974 3576
rect 6460 3538 6512 3544
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6380 2650 6408 3470
rect 6472 3194 6500 3538
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6568 3292 6864 3312
rect 6624 3290 6648 3292
rect 6704 3290 6728 3292
rect 6784 3290 6808 3292
rect 6646 3238 6648 3290
rect 6710 3238 6722 3290
rect 6784 3238 6786 3290
rect 6624 3236 6648 3238
rect 6704 3236 6728 3238
rect 6784 3236 6808 3238
rect 6568 3216 6864 3236
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6458 3088 6514 3097
rect 6458 3023 6514 3032
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6104 2230 6316 2258
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 6184 1828 6236 1834
rect 6184 1770 6236 1776
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 5906 1048 5962 1057
rect 5906 983 5962 992
rect 5920 800 5948 983
rect 6012 800 6040 1663
rect 6196 800 6224 1770
rect 6288 800 6316 2230
rect 6472 2122 6500 3023
rect 6552 2372 6604 2378
rect 6656 2360 6684 3023
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6840 2854 6868 2887
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6932 2582 6960 3402
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7024 2428 7052 8842
rect 7116 8616 7144 9030
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7196 8628 7248 8634
rect 7116 8588 7196 8616
rect 7196 8570 7248 8576
rect 7104 8424 7156 8430
rect 7300 8412 7328 9658
rect 7392 9518 7420 9862
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7156 8384 7328 8412
rect 7104 8366 7156 8372
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 6934 7144 7686
rect 7208 7546 7236 7822
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6934 7236 7142
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7208 6440 7236 6870
rect 7116 6412 7236 6440
rect 7116 6089 7144 6412
rect 7194 6352 7250 6361
rect 7194 6287 7250 6296
rect 7102 6080 7158 6089
rect 7102 6015 7158 6024
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6604 2332 6684 2360
rect 6932 2400 7052 2428
rect 6552 2314 6604 2320
rect 6568 2204 6864 2224
rect 6624 2202 6648 2204
rect 6704 2202 6728 2204
rect 6784 2202 6808 2204
rect 6646 2150 6648 2202
rect 6710 2150 6722 2202
rect 6784 2150 6786 2202
rect 6624 2148 6648 2150
rect 6704 2148 6728 2150
rect 6784 2148 6808 2150
rect 6568 2128 6864 2148
rect 6380 2106 6500 2122
rect 6368 2100 6500 2106
rect 6420 2094 6500 2100
rect 6368 2042 6420 2048
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6734 2000 6790 2009
rect 6366 1864 6422 1873
rect 6366 1799 6422 1808
rect 6380 1222 6408 1799
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6472 800 6500 1974
rect 6564 800 6592 1974
rect 6734 1935 6790 1944
rect 6828 1964 6880 1970
rect 6748 800 6776 1935
rect 6828 1906 6880 1912
rect 6840 800 6868 1906
rect 6932 800 6960 2400
rect 7116 800 7144 5850
rect 7208 800 7236 6287
rect 7300 2582 7328 7414
rect 7392 5914 7420 8978
rect 7484 6254 7512 10095
rect 7576 8401 7604 10220
rect 7668 9450 7696 10390
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7562 8392 7618 8401
rect 7562 8327 7618 8336
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7576 5409 7604 7686
rect 7668 6474 7696 9046
rect 7760 8090 7788 11766
rect 7944 11082 7972 12600
rect 8024 12582 8076 12588
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8128 11529 8156 12106
rect 8220 12102 8248 12650
rect 8588 12628 8616 12854
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8312 12600 8616 12628
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8312 11694 8340 12600
rect 8438 12540 8734 12560
rect 8494 12538 8518 12540
rect 8574 12538 8598 12540
rect 8654 12538 8678 12540
rect 8516 12486 8518 12538
rect 8580 12486 8592 12538
rect 8654 12486 8656 12538
rect 8494 12484 8518 12486
rect 8574 12484 8598 12486
rect 8654 12484 8678 12486
rect 8438 12464 8734 12484
rect 8772 12442 8800 12718
rect 8864 12442 8892 12786
rect 9048 12782 9076 13398
rect 9692 12986 9720 14818
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 12102 8984 12242
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8956 11558 8984 12038
rect 8944 11552 8996 11558
rect 8114 11520 8170 11529
rect 8944 11494 8996 11500
rect 8114 11455 8170 11464
rect 8128 11218 8156 11455
rect 8438 11452 8734 11472
rect 8494 11450 8518 11452
rect 8574 11450 8598 11452
rect 8654 11450 8678 11452
rect 8516 11398 8518 11450
rect 8580 11398 8592 11450
rect 8654 11398 8656 11450
rect 8494 11396 8518 11398
rect 8574 11396 8598 11398
rect 8654 11396 8678 11398
rect 8438 11376 8734 11396
rect 8956 11286 8984 11494
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8944 11280 8996 11286
rect 9140 11268 9168 12786
rect 10060 12782 10088 13466
rect 11164 13138 11192 14818
rect 11164 13110 11284 13138
rect 10309 13084 10605 13104
rect 10365 13082 10389 13084
rect 10445 13082 10469 13084
rect 10525 13082 10549 13084
rect 10387 13030 10389 13082
rect 10451 13030 10463 13082
rect 10525 13030 10527 13082
rect 10365 13028 10389 13030
rect 10445 13028 10469 13030
rect 10525 13028 10549 13030
rect 10309 13008 10605 13028
rect 11256 12986 11284 13110
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9232 11898 9260 12718
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9324 12306 9352 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11898 9444 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9232 11694 9260 11834
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9140 11240 9352 11268
rect 8944 11222 8996 11228
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7838 10568 7894 10577
rect 8312 10538 8340 11222
rect 8496 10810 8524 11222
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8864 10606 8892 10950
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 7838 10503 7894 10512
rect 8300 10532 8352 10538
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7002 7880 10503
rect 8300 10474 8352 10480
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7760 6882 7788 6938
rect 7944 6882 7972 9862
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7760 6854 7972 6882
rect 7668 6446 7788 6474
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7472 5160 7524 5166
rect 7668 5114 7696 5714
rect 7472 5102 7524 5108
rect 7392 4282 7420 5102
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7484 4214 7512 5102
rect 7576 5086 7696 5114
rect 7576 4486 7604 5086
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4758 7696 4966
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7654 4584 7710 4593
rect 7654 4519 7710 4528
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7472 4072 7524 4078
rect 7378 4040 7434 4049
rect 7472 4014 7524 4020
rect 7378 3975 7434 3984
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7392 800 7420 3975
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 3126 7512 3538
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7576 2990 7604 4422
rect 7668 3584 7696 4519
rect 7760 3738 7788 6446
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5370 7880 6190
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5914 7972 6054
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7852 5166 7880 5306
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7838 4856 7894 4865
rect 7838 4791 7894 4800
rect 7852 4758 7880 4791
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7748 3596 7800 3602
rect 7668 3556 7748 3584
rect 7748 3538 7800 3544
rect 7564 2984 7616 2990
rect 7616 2944 7696 2972
rect 7564 2926 7616 2932
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7484 800 7512 2518
rect 7576 800 7604 2751
rect 7668 2514 7696 2944
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7760 2446 7788 3538
rect 7852 3534 7880 4014
rect 7944 3942 7972 4966
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7852 3194 7880 3470
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7838 2544 7894 2553
rect 7838 2479 7894 2488
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7748 1420 7800 1426
rect 7748 1362 7800 1368
rect 7760 800 7788 1362
rect 7852 800 7880 2479
rect 7944 2310 7972 3878
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8036 800 8064 8978
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8128 5914 8156 6258
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 4049 8156 5510
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3534 8156 3878
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8114 2952 8170 2961
rect 8114 2887 8170 2896
rect 8128 800 8156 2887
rect 8220 800 8248 10066
rect 8312 9178 8340 10474
rect 8438 10364 8734 10384
rect 8494 10362 8518 10364
rect 8574 10362 8598 10364
rect 8654 10362 8678 10364
rect 8516 10310 8518 10362
rect 8580 10310 8592 10362
rect 8654 10310 8656 10362
rect 8494 10308 8518 10310
rect 8574 10308 8598 10310
rect 8654 10308 8678 10310
rect 8438 10288 8734 10308
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8404 9654 8432 10134
rect 8668 10124 8720 10130
rect 8720 10084 8800 10112
rect 8668 10066 8720 10072
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8438 9276 8734 9296
rect 8494 9274 8518 9276
rect 8574 9274 8598 9276
rect 8654 9274 8678 9276
rect 8516 9222 8518 9274
rect 8580 9222 8592 9274
rect 8654 9222 8656 9274
rect 8494 9220 8518 9222
rect 8574 9220 8598 9222
rect 8654 9220 8678 9222
rect 8438 9200 8734 9220
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8312 8498 8340 8978
rect 8680 8906 8708 8978
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 7993 8340 8434
rect 8438 8188 8734 8208
rect 8494 8186 8518 8188
rect 8574 8186 8598 8188
rect 8654 8186 8678 8188
rect 8516 8134 8518 8186
rect 8580 8134 8592 8186
rect 8654 8134 8656 8186
rect 8494 8132 8518 8134
rect 8574 8132 8598 8134
rect 8654 8132 8678 8134
rect 8438 8112 8734 8132
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7342 8340 7822
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6730 8340 7278
rect 8438 7100 8734 7120
rect 8494 7098 8518 7100
rect 8574 7098 8598 7100
rect 8654 7098 8678 7100
rect 8516 7046 8518 7098
rect 8580 7046 8592 7098
rect 8654 7046 8656 7098
rect 8494 7044 8518 7046
rect 8574 7044 8598 7046
rect 8654 7044 8678 7046
rect 8438 7024 8734 7044
rect 8772 6984 8800 10084
rect 8864 7993 8892 10202
rect 8956 10130 8984 11222
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9048 10470 9076 11154
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10606 9260 10950
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8956 9722 8984 10066
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9048 9518 9076 10406
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8956 8634 8984 8978
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8850 7984 8906 7993
rect 8850 7919 8906 7928
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8680 6956 8800 6984
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8496 6361 8524 6734
rect 8680 6662 8708 6956
rect 8864 6866 8892 7754
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8772 6458 8800 6802
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8482 6352 8538 6361
rect 8956 6304 8984 8298
rect 9140 8072 9168 9862
rect 9232 9722 9260 9930
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 8430 9260 8910
rect 9324 8906 9352 11240
rect 9416 10130 9444 11834
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9324 8566 9352 8842
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9140 8044 9260 8072
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 6866 9076 7686
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9140 6730 9168 7890
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8482 6287 8484 6296
rect 8536 6287 8538 6296
rect 8484 6258 8536 6264
rect 8864 6276 8984 6304
rect 8438 6012 8734 6032
rect 8494 6010 8518 6012
rect 8574 6010 8598 6012
rect 8654 6010 8678 6012
rect 8516 5958 8518 6010
rect 8580 5958 8592 6010
rect 8654 5958 8656 6010
rect 8494 5956 8518 5958
rect 8574 5956 8598 5958
rect 8654 5956 8678 5958
rect 8438 5936 8734 5956
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8300 5568 8352 5574
rect 8588 5545 8616 5714
rect 8300 5510 8352 5516
rect 8574 5536 8630 5545
rect 8312 4146 8340 5510
rect 8574 5471 8630 5480
rect 8588 5166 8616 5471
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8438 4924 8734 4944
rect 8494 4922 8518 4924
rect 8574 4922 8598 4924
rect 8654 4922 8678 4924
rect 8516 4870 8518 4922
rect 8580 4870 8592 4922
rect 8654 4870 8656 4922
rect 8494 4868 8518 4870
rect 8574 4868 8598 4870
rect 8654 4868 8678 4870
rect 8438 4848 8734 4868
rect 8772 4826 8800 5034
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8404 4010 8432 4694
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 8312 3720 8340 3839
rect 8438 3836 8734 3856
rect 8494 3834 8518 3836
rect 8574 3834 8598 3836
rect 8654 3834 8678 3836
rect 8516 3782 8518 3834
rect 8580 3782 8592 3834
rect 8654 3782 8656 3834
rect 8494 3780 8518 3782
rect 8574 3780 8598 3782
rect 8654 3780 8678 3782
rect 8438 3760 8734 3780
rect 8312 3692 8524 3720
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8312 2650 8340 3538
rect 8404 2922 8432 3538
rect 8496 3097 8524 3692
rect 8758 3632 8814 3641
rect 8758 3567 8760 3576
rect 8812 3567 8814 3576
rect 8760 3538 8812 3544
rect 8666 3496 8722 3505
rect 8666 3431 8722 3440
rect 8680 3126 8708 3431
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8668 3120 8720 3126
rect 8482 3088 8538 3097
rect 8668 3062 8720 3068
rect 8482 3023 8538 3032
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8438 2748 8734 2768
rect 8494 2746 8518 2748
rect 8574 2746 8598 2748
rect 8654 2746 8678 2748
rect 8516 2694 8518 2746
rect 8580 2694 8592 2746
rect 8654 2694 8656 2746
rect 8494 2692 8518 2694
rect 8574 2692 8598 2694
rect 8654 2692 8678 2694
rect 8438 2672 8734 2692
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8772 2582 8800 3159
rect 8760 2576 8812 2582
rect 8482 2544 8538 2553
rect 8482 2479 8538 2488
rect 8666 2544 8722 2553
rect 8760 2518 8812 2524
rect 8666 2479 8668 2488
rect 8390 2408 8446 2417
rect 8390 2343 8446 2352
rect 8404 800 8432 2343
rect 8496 800 8524 2479
rect 8720 2479 8722 2488
rect 8668 2450 8720 2456
rect 8666 2272 8722 2281
rect 8666 2207 8722 2216
rect 8680 800 8708 2207
rect 8758 1728 8814 1737
rect 8758 1663 8814 1672
rect 8772 800 8800 1663
rect 8864 1426 8892 6276
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8956 5846 8984 6122
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8942 5264 8998 5273
rect 8942 5199 8998 5208
rect 8956 5166 8984 5199
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4078 8984 4422
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 2038 8984 3878
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 8852 1420 8904 1426
rect 8852 1362 8904 1368
rect 8850 1320 8906 1329
rect 8850 1255 8906 1264
rect 8864 800 8892 1255
rect 9048 800 9076 6598
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5370 9168 5714
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9126 5264 9182 5273
rect 9126 5199 9128 5208
rect 9180 5199 9182 5208
rect 9128 5170 9180 5176
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9140 2394 9168 4218
rect 9232 2582 9260 8044
rect 9324 7886 9352 8502
rect 9312 7880 9364 7886
rect 9364 7840 9444 7868
rect 9312 7822 9364 7828
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7342 9352 7686
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6254 9352 7142
rect 9416 6866 9444 7840
rect 9508 7528 9536 12582
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9968 12396 10180 12424
rect 9600 9654 9628 12378
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9784 12209 9812 12310
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9770 12200 9826 12209
rect 9770 12135 9826 12144
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9692 11218 9720 11630
rect 9784 11626 9812 12038
rect 9876 11898 9904 12242
rect 9968 12238 9996 12396
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9968 11694 9996 12174
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9784 11257 9812 11562
rect 9876 11268 9904 11630
rect 10060 11354 10088 12242
rect 10152 11608 10180 12396
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10309 11996 10605 12016
rect 10365 11994 10389 11996
rect 10445 11994 10469 11996
rect 10525 11994 10549 11996
rect 10387 11942 10389 11994
rect 10451 11942 10463 11994
rect 10525 11942 10527 11994
rect 10365 11940 10389 11942
rect 10445 11940 10469 11942
rect 10525 11940 10549 11942
rect 10309 11920 10605 11940
rect 10796 11762 10824 12038
rect 10508 11756 10560 11762
rect 10784 11756 10836 11762
rect 10560 11716 10732 11744
rect 10508 11698 10560 11704
rect 10416 11688 10468 11694
rect 10414 11656 10416 11665
rect 10468 11656 10470 11665
rect 10232 11620 10284 11626
rect 10152 11580 10232 11608
rect 10414 11591 10470 11600
rect 10232 11562 10284 11568
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9956 11280 10008 11286
rect 9770 11248 9826 11257
rect 9680 11212 9732 11218
rect 9770 11183 9826 11192
rect 9876 11240 9956 11268
rect 9680 11154 9732 11160
rect 9678 11112 9734 11121
rect 9678 11047 9734 11056
rect 9692 10742 9720 11047
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9784 10674 9812 10950
rect 9876 10742 9904 11240
rect 9956 11222 10008 11228
rect 10046 11248 10102 11257
rect 10046 11183 10102 11192
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9784 10554 9812 10610
rect 10060 10606 10088 11183
rect 10140 11144 10192 11150
rect 10336 11121 10364 11494
rect 10416 11212 10468 11218
rect 10520 11200 10548 11698
rect 10704 11642 10732 11716
rect 10784 11698 10836 11704
rect 11164 11694 11192 12854
rect 12636 12850 12664 14818
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11256 11898 11284 12135
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11532 11694 11560 12582
rect 11624 12442 11652 12650
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 12306 11652 12378
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11152 11688 11204 11694
rect 10704 11614 10824 11642
rect 11520 11688 11572 11694
rect 11152 11630 11204 11636
rect 11242 11656 11298 11665
rect 10600 11348 10652 11354
rect 10652 11308 10732 11336
rect 10600 11290 10652 11296
rect 10468 11172 10548 11200
rect 10416 11154 10468 11160
rect 10140 11086 10192 11092
rect 10322 11112 10378 11121
rect 10048 10600 10100 10606
rect 9692 10266 9720 10542
rect 9784 10526 9904 10554
rect 10048 10542 10100 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9784 10010 9812 10406
rect 9876 10198 9904 10526
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9864 10056 9916 10062
rect 9784 10004 9864 10010
rect 9784 9998 9916 10004
rect 9784 9982 9904 9998
rect 10060 9994 10088 10542
rect 10152 10470 10180 11086
rect 10322 11047 10378 11056
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10606 10272 10950
rect 10309 10908 10605 10928
rect 10365 10906 10389 10908
rect 10445 10906 10469 10908
rect 10525 10906 10549 10908
rect 10387 10854 10389 10906
rect 10451 10854 10463 10906
rect 10525 10854 10527 10906
rect 10365 10852 10389 10854
rect 10445 10852 10469 10854
rect 10525 10852 10549 10854
rect 10309 10832 10605 10852
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10048 9988 10100 9994
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9692 9178 9720 9862
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 8974 9812 9982
rect 10048 9930 10100 9936
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9586 9996 9862
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9450 9996 9522
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10060 9330 10088 9930
rect 10244 9722 10272 10406
rect 10704 10266 10732 11308
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10309 9820 10605 9840
rect 10365 9818 10389 9820
rect 10445 9818 10469 9820
rect 10525 9818 10549 9820
rect 10387 9766 10389 9818
rect 10451 9766 10463 9818
rect 10525 9766 10527 9818
rect 10365 9764 10389 9766
rect 10445 9764 10469 9766
rect 10525 9764 10549 9766
rect 10309 9744 10605 9764
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 9876 9302 10088 9330
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8634 9812 8910
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8430 9904 9302
rect 10152 9042 10180 9454
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9588 7540 9640 7546
rect 9508 7500 9588 7528
rect 9588 7482 9640 7488
rect 9692 7449 9720 7754
rect 9678 7440 9734 7449
rect 9678 7375 9734 7384
rect 9692 6934 9720 7375
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9416 6066 9444 6802
rect 9324 6038 9444 6066
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9324 5914 9352 6038
rect 9508 5930 9536 6054
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5902 9536 5930
rect 9324 5302 9352 5850
rect 9416 5642 9444 5902
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9324 4078 9352 5102
rect 9416 4758 9444 5578
rect 9508 5370 9536 5782
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5534 9628 5714
rect 9692 5642 9720 6870
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9600 5506 9720 5534
rect 9586 5400 9642 5409
rect 9496 5364 9548 5370
rect 9692 5370 9720 5506
rect 9586 5335 9642 5344
rect 9680 5364 9732 5370
rect 9496 5306 9548 5312
rect 9494 4856 9550 4865
rect 9494 4791 9496 4800
rect 9548 4791 9550 4800
rect 9496 4762 9548 4768
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 2922 9352 3878
rect 9416 3126 9444 3975
rect 9508 3398 9536 4218
rect 9600 3602 9628 5335
rect 9680 5306 9732 5312
rect 9692 5273 9720 5306
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9692 4622 9720 5034
rect 9680 4616 9732 4622
rect 9678 4584 9680 4593
rect 9732 4584 9734 4593
rect 9678 4519 9734 4528
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9692 3641 9720 3674
rect 9784 3670 9812 8366
rect 9876 7886 9904 8366
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9864 7880 9916 7886
rect 9968 7857 9996 8026
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9864 7822 9916 7828
rect 9954 7848 10010 7857
rect 9954 7783 10010 7792
rect 9956 7744 10008 7750
rect 9862 7712 9918 7721
rect 9956 7686 10008 7692
rect 9862 7647 9918 7656
rect 9876 7274 9904 7647
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6361 9904 7210
rect 9862 6352 9918 6361
rect 9862 6287 9864 6296
rect 9916 6287 9918 6296
rect 9864 6258 9916 6264
rect 9876 5234 9904 6258
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9968 4570 9996 7686
rect 10060 7546 10088 7958
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10060 7002 10088 7482
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 5545 10088 5646
rect 10046 5536 10102 5545
rect 10046 5471 10102 5480
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4826 10088 5102
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9968 4542 10088 4570
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 3664 9824 3670
rect 9678 3632 9734 3641
rect 9588 3596 9640 3602
rect 9772 3606 9824 3612
rect 9678 3567 9734 3576
rect 9588 3538 9640 3544
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9140 2366 9260 2394
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 800 9168 2246
rect 9232 1766 9260 2366
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 9324 800 9352 2314
rect 9416 800 9444 2790
rect 9508 800 9536 2994
rect 9600 2582 9628 3402
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9692 800 9720 3470
rect 9784 800 9812 3470
rect 9876 2650 9904 4014
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9862 2544 9918 2553
rect 9862 2479 9864 2488
rect 9916 2479 9918 2488
rect 9864 2450 9916 2456
rect 9968 800 9996 4422
rect 10060 3176 10088 4542
rect 10152 3670 10180 7686
rect 10244 5681 10272 9454
rect 10520 8906 10548 9590
rect 10704 9450 10732 10202
rect 10796 9586 10824 11614
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10888 10810 10916 11222
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9722 10916 10066
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10309 8732 10605 8752
rect 10365 8730 10389 8732
rect 10445 8730 10469 8732
rect 10525 8730 10549 8732
rect 10387 8678 10389 8730
rect 10451 8678 10463 8730
rect 10525 8678 10527 8730
rect 10365 8676 10389 8678
rect 10445 8676 10469 8678
rect 10525 8676 10549 8678
rect 10309 8656 10605 8676
rect 10796 8498 10824 8774
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10309 7644 10605 7664
rect 10365 7642 10389 7644
rect 10445 7642 10469 7644
rect 10525 7642 10549 7644
rect 10387 7590 10389 7642
rect 10451 7590 10463 7642
rect 10525 7590 10527 7642
rect 10365 7588 10389 7590
rect 10445 7588 10469 7590
rect 10525 7588 10549 7590
rect 10309 7568 10605 7588
rect 10704 7546 10732 7958
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 7472 10376 7478
rect 10322 7440 10324 7449
rect 10376 7440 10378 7449
rect 10888 7426 10916 9318
rect 10980 7993 11008 11494
rect 11164 10606 11192 11630
rect 11520 11630 11572 11636
rect 11242 11591 11298 11600
rect 11256 11218 11284 11591
rect 11532 11218 11560 11630
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11256 10810 11284 11154
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11348 10198 11376 10950
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10322 7375 10378 7384
rect 10796 7398 10916 7426
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10506 7032 10562 7041
rect 10506 6967 10508 6976
rect 10560 6967 10562 6976
rect 10508 6938 10560 6944
rect 10508 6792 10560 6798
rect 10612 6780 10640 7278
rect 10560 6752 10640 6780
rect 10508 6734 10560 6740
rect 10309 6556 10605 6576
rect 10365 6554 10389 6556
rect 10445 6554 10469 6556
rect 10525 6554 10549 6556
rect 10387 6502 10389 6554
rect 10451 6502 10463 6554
rect 10525 6502 10527 6554
rect 10365 6500 10389 6502
rect 10445 6500 10469 6502
rect 10525 6500 10549 6502
rect 10309 6480 10605 6500
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5794 10640 6054
rect 10704 5914 10732 6122
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10612 5766 10732 5794
rect 10230 5672 10286 5681
rect 10230 5607 10286 5616
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5166 10272 5510
rect 10309 5468 10605 5488
rect 10365 5466 10389 5468
rect 10445 5466 10469 5468
rect 10525 5466 10549 5468
rect 10387 5414 10389 5466
rect 10451 5414 10463 5466
rect 10525 5414 10527 5466
rect 10365 5412 10389 5414
rect 10445 5412 10469 5414
rect 10525 5412 10549 5414
rect 10309 5392 10605 5412
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10598 5128 10654 5137
rect 10598 5063 10654 5072
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10060 3148 10180 3176
rect 10046 3088 10102 3097
rect 10046 3023 10102 3032
rect 10060 2990 10088 3023
rect 10152 2990 10180 3148
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10244 2530 10272 4966
rect 10612 4570 10640 5063
rect 10704 4758 10732 5766
rect 10796 4826 10824 7398
rect 10876 7336 10928 7342
rect 10980 7324 11008 7686
rect 11072 7342 11100 7890
rect 10928 7296 11008 7324
rect 11060 7336 11112 7342
rect 10876 7278 10928 7284
rect 11060 7278 11112 7284
rect 10888 7002 10916 7278
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11164 6882 11192 9522
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11072 6854 11192 6882
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 5846 11008 6598
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10784 4684 10836 4690
rect 10888 4672 10916 5578
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10980 5098 11008 5510
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10836 4644 10916 4672
rect 10784 4626 10836 4632
rect 10968 4616 11020 4622
rect 10966 4584 10968 4593
rect 11020 4584 11022 4593
rect 10612 4542 10824 4570
rect 10309 4380 10605 4400
rect 10365 4378 10389 4380
rect 10445 4378 10469 4380
rect 10525 4378 10549 4380
rect 10387 4326 10389 4378
rect 10451 4326 10463 4378
rect 10525 4326 10527 4378
rect 10365 4324 10389 4326
rect 10445 4324 10469 4326
rect 10525 4324 10549 4326
rect 10309 4304 10605 4324
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10309 3292 10605 3312
rect 10365 3290 10389 3292
rect 10445 3290 10469 3292
rect 10525 3290 10549 3292
rect 10387 3238 10389 3290
rect 10451 3238 10463 3290
rect 10525 3238 10527 3290
rect 10365 3236 10389 3238
rect 10445 3236 10469 3238
rect 10525 3236 10549 3238
rect 10309 3216 10605 3236
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10428 2922 10456 3062
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10336 2650 10364 2858
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10152 2502 10272 2530
rect 10322 2544 10378 2553
rect 10520 2514 10548 3062
rect 10600 2576 10652 2582
rect 10704 2564 10732 3878
rect 10796 3534 10824 4542
rect 10966 4519 11022 4528
rect 10968 3596 11020 3602
rect 11072 3584 11100 6854
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11020 3556 11100 3584
rect 10968 3538 11020 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11058 3496 11114 3505
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10968 3460 11020 3466
rect 11058 3431 11060 3440
rect 10968 3402 11020 3408
rect 11112 3431 11114 3440
rect 11060 3402 11112 3408
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10652 2536 10732 2564
rect 10600 2518 10652 2524
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10060 800 10088 1974
rect 10152 800 10180 2502
rect 10322 2479 10324 2488
rect 10376 2479 10378 2488
rect 10508 2508 10560 2514
rect 10324 2450 10376 2456
rect 10508 2450 10560 2456
rect 10796 2417 10824 3334
rect 10888 2446 10916 3402
rect 10980 2854 11008 3402
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10876 2440 10928 2446
rect 10230 2408 10286 2417
rect 10230 2343 10286 2352
rect 10782 2408 10838 2417
rect 10876 2382 10928 2388
rect 10782 2343 10838 2352
rect 10968 2372 11020 2378
rect 10244 1986 10272 2343
rect 10968 2314 11020 2320
rect 10692 2304 10744 2310
rect 10876 2304 10928 2310
rect 10692 2246 10744 2252
rect 10796 2264 10876 2292
rect 10309 2204 10605 2224
rect 10365 2202 10389 2204
rect 10445 2202 10469 2204
rect 10525 2202 10549 2204
rect 10387 2150 10389 2202
rect 10451 2150 10463 2202
rect 10525 2150 10527 2202
rect 10365 2148 10389 2150
rect 10445 2148 10469 2150
rect 10525 2148 10549 2150
rect 10309 2128 10605 2148
rect 10244 1958 10364 1986
rect 10336 800 10364 1958
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10428 800 10456 1702
rect 10704 1170 10732 2246
rect 10612 1142 10732 1170
rect 10612 800 10640 1142
rect 10796 1034 10824 2264
rect 10876 2246 10928 2252
rect 10704 1006 10824 1034
rect 10704 800 10732 1006
rect 10784 944 10836 950
rect 10784 886 10836 892
rect 10796 800 10824 886
rect 10980 800 11008 2314
rect 11072 800 11100 2790
rect 11164 2582 11192 6734
rect 11256 6322 11284 7278
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11256 3398 11284 5782
rect 11348 4758 11376 8774
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11348 4010 11376 4558
rect 11440 4078 11468 8774
rect 11532 5166 11560 9454
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11624 4672 11652 6598
rect 11532 4644 11652 4672
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11256 800 11284 3130
rect 11348 800 11376 3334
rect 11440 800 11468 3402
rect 11532 2582 11560 4644
rect 11716 4570 11744 7278
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5710 11836 6054
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11624 4542 11744 4570
rect 11624 3670 11652 4542
rect 11900 4078 11928 8366
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 950 11560 2246
rect 11520 944 11572 950
rect 11520 886 11572 892
rect 11624 800 11652 2926
rect 11716 800 11744 3878
rect 11992 3670 12020 7686
rect 12084 4622 12112 8774
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 800 11928 3470
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11992 800 12020 3062
rect 12084 800 12112 3946
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 800 12296 3538
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12360 800 12388 2586
rect 12452 2553 12480 4762
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12438 2544 12494 2553
rect 12438 2479 12494 2488
rect 12544 800 12572 4490
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 800 12664 4082
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 800 12756 3674
rect 12912 800 12940 4422
rect 13174 3632 13230 3641
rect 13174 3567 13230 3576
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13004 800 13032 2382
rect 13188 800 13216 3567
rect 13280 800 13308 5034
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 386 0 442 800
rect 478 0 534 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
<< via2 >>
rect 570 12416 626 12472
rect 754 7248 810 7304
rect 754 3984 810 4040
rect 662 2896 718 2952
rect 1858 12588 1860 12608
rect 1860 12588 1912 12608
rect 1912 12588 1914 12608
rect 1858 12552 1914 12588
rect 1306 12144 1362 12200
rect 938 2896 994 2952
rect 1122 2896 1178 2952
rect 1398 9016 1454 9072
rect 1490 8744 1546 8800
rect 1766 8472 1822 8528
rect 1582 6704 1638 6760
rect 1674 3984 1730 4040
rect 1950 9968 2006 10024
rect 1858 6704 1914 6760
rect 2226 10648 2282 10704
rect 2410 12588 2412 12608
rect 2412 12588 2464 12608
rect 2464 12588 2466 12608
rect 2410 12552 2466 12588
rect 2410 8744 2466 8800
rect 2226 8608 2282 8664
rect 2134 7928 2190 7984
rect 1858 3576 1914 3632
rect 1766 3168 1822 3224
rect 1858 2896 1914 2952
rect 1858 2760 1914 2816
rect 2318 7384 2374 7440
rect 2318 6160 2374 6216
rect 2826 13082 2882 13084
rect 2906 13082 2962 13084
rect 2986 13082 3042 13084
rect 3066 13082 3122 13084
rect 2826 13030 2852 13082
rect 2852 13030 2882 13082
rect 2906 13030 2916 13082
rect 2916 13030 2962 13082
rect 2986 13030 3032 13082
rect 3032 13030 3042 13082
rect 3066 13030 3096 13082
rect 3096 13030 3122 13082
rect 2826 13028 2882 13030
rect 2906 13028 2962 13030
rect 2986 13028 3042 13030
rect 3066 13028 3122 13030
rect 2826 11994 2882 11996
rect 2906 11994 2962 11996
rect 2986 11994 3042 11996
rect 3066 11994 3122 11996
rect 2826 11942 2852 11994
rect 2852 11942 2882 11994
rect 2906 11942 2916 11994
rect 2916 11942 2962 11994
rect 2986 11942 3032 11994
rect 3032 11942 3042 11994
rect 3066 11942 3096 11994
rect 3096 11942 3122 11994
rect 2826 11940 2882 11942
rect 2906 11940 2962 11942
rect 2986 11940 3042 11942
rect 3066 11940 3122 11942
rect 2686 11056 2742 11112
rect 2826 10906 2882 10908
rect 2906 10906 2962 10908
rect 2986 10906 3042 10908
rect 3066 10906 3122 10908
rect 2826 10854 2852 10906
rect 2852 10854 2882 10906
rect 2906 10854 2916 10906
rect 2916 10854 2962 10906
rect 2986 10854 3032 10906
rect 3032 10854 3042 10906
rect 3066 10854 3096 10906
rect 3096 10854 3122 10906
rect 2826 10852 2882 10854
rect 2906 10852 2962 10854
rect 2986 10852 3042 10854
rect 3066 10852 3122 10854
rect 2870 10412 2872 10432
rect 2872 10412 2924 10432
rect 2924 10412 2926 10432
rect 2870 10376 2926 10412
rect 3238 10376 3294 10432
rect 3422 10104 3478 10160
rect 2826 9818 2882 9820
rect 2906 9818 2962 9820
rect 2986 9818 3042 9820
rect 3066 9818 3122 9820
rect 2826 9766 2852 9818
rect 2852 9766 2882 9818
rect 2906 9766 2916 9818
rect 2916 9766 2962 9818
rect 2986 9766 3032 9818
rect 3032 9766 3042 9818
rect 3066 9766 3096 9818
rect 3096 9766 3122 9818
rect 2826 9764 2882 9766
rect 2906 9764 2962 9766
rect 2986 9764 3042 9766
rect 3066 9764 3122 9766
rect 2826 8730 2882 8732
rect 2906 8730 2962 8732
rect 2986 8730 3042 8732
rect 3066 8730 3122 8732
rect 2826 8678 2852 8730
rect 2852 8678 2882 8730
rect 2906 8678 2916 8730
rect 2916 8678 2962 8730
rect 2986 8678 3032 8730
rect 3032 8678 3042 8730
rect 3066 8678 3096 8730
rect 3096 8678 3122 8730
rect 2826 8676 2882 8678
rect 2906 8676 2962 8678
rect 2986 8676 3042 8678
rect 3066 8676 3122 8678
rect 2778 8492 2834 8528
rect 2778 8472 2780 8492
rect 2780 8472 2832 8492
rect 2832 8472 2834 8492
rect 2962 8356 3018 8392
rect 2962 8336 2964 8356
rect 2964 8336 3016 8356
rect 3016 8336 3018 8356
rect 2826 7642 2882 7644
rect 2906 7642 2962 7644
rect 2986 7642 3042 7644
rect 3066 7642 3122 7644
rect 2826 7590 2852 7642
rect 2852 7590 2882 7642
rect 2906 7590 2916 7642
rect 2916 7590 2962 7642
rect 2986 7590 3032 7642
rect 3032 7590 3042 7642
rect 3066 7590 3096 7642
rect 3096 7590 3122 7642
rect 2826 7588 2882 7590
rect 2906 7588 2962 7590
rect 2986 7588 3042 7590
rect 3066 7588 3122 7590
rect 2778 7384 2834 7440
rect 3054 7420 3056 7440
rect 3056 7420 3108 7440
rect 3108 7420 3110 7440
rect 2686 6976 2742 7032
rect 3054 7384 3110 7420
rect 2962 6976 3018 7032
rect 2826 6554 2882 6556
rect 2906 6554 2962 6556
rect 2986 6554 3042 6556
rect 3066 6554 3122 6556
rect 2826 6502 2852 6554
rect 2852 6502 2882 6554
rect 2906 6502 2916 6554
rect 2916 6502 2962 6554
rect 2986 6502 3032 6554
rect 3032 6502 3042 6554
rect 3066 6502 3096 6554
rect 3096 6502 3122 6554
rect 2826 6500 2882 6502
rect 2906 6500 2962 6502
rect 2986 6500 3042 6502
rect 3066 6500 3122 6502
rect 2318 2760 2374 2816
rect 3238 8880 3294 8936
rect 4158 12416 4214 12472
rect 3790 10104 3846 10160
rect 3514 9424 3570 9480
rect 3330 6840 3386 6896
rect 3330 6704 3386 6760
rect 3238 5888 3294 5944
rect 2962 5616 3018 5672
rect 2826 5466 2882 5468
rect 2906 5466 2962 5468
rect 2986 5466 3042 5468
rect 3066 5466 3122 5468
rect 2826 5414 2852 5466
rect 2852 5414 2882 5466
rect 2906 5414 2916 5466
rect 2916 5414 2962 5466
rect 2986 5414 3032 5466
rect 3032 5414 3042 5466
rect 3066 5414 3096 5466
rect 3096 5414 3122 5466
rect 2826 5412 2882 5414
rect 2906 5412 2962 5414
rect 2986 5412 3042 5414
rect 3066 5412 3122 5414
rect 2826 4378 2882 4380
rect 2906 4378 2962 4380
rect 2986 4378 3042 4380
rect 3066 4378 3122 4380
rect 2826 4326 2852 4378
rect 2852 4326 2882 4378
rect 2906 4326 2916 4378
rect 2916 4326 2962 4378
rect 2986 4326 3032 4378
rect 3032 4326 3042 4378
rect 3066 4326 3096 4378
rect 3096 4326 3122 4378
rect 2826 4324 2882 4326
rect 2906 4324 2962 4326
rect 2986 4324 3042 4326
rect 3066 4324 3122 4326
rect 3330 3848 3386 3904
rect 3698 7384 3754 7440
rect 3698 6432 3754 6488
rect 3606 4528 3662 4584
rect 2826 3290 2882 3292
rect 2906 3290 2962 3292
rect 2986 3290 3042 3292
rect 3066 3290 3122 3292
rect 2826 3238 2852 3290
rect 2852 3238 2882 3290
rect 2906 3238 2916 3290
rect 2916 3238 2962 3290
rect 2986 3238 3032 3290
rect 3032 3238 3042 3290
rect 3066 3238 3096 3290
rect 3096 3238 3122 3290
rect 2826 3236 2882 3238
rect 2906 3236 2962 3238
rect 2986 3236 3042 3238
rect 3066 3236 3122 3238
rect 3238 3032 3294 3088
rect 3146 2896 3202 2952
rect 2870 2524 2872 2544
rect 2872 2524 2924 2544
rect 2924 2524 2926 2544
rect 2870 2488 2926 2524
rect 2826 2202 2882 2204
rect 2906 2202 2962 2204
rect 2986 2202 3042 2204
rect 3066 2202 3122 2204
rect 2826 2150 2852 2202
rect 2852 2150 2882 2202
rect 2906 2150 2916 2202
rect 2916 2150 2962 2202
rect 2986 2150 3032 2202
rect 3032 2150 3042 2202
rect 3066 2150 3096 2202
rect 3096 2150 3122 2202
rect 2826 2148 2882 2150
rect 2906 2148 2962 2150
rect 2986 2148 3042 2150
rect 3066 2148 3122 2150
rect 2594 1808 2650 1864
rect 4697 12538 4753 12540
rect 4777 12538 4833 12540
rect 4857 12538 4913 12540
rect 4937 12538 4993 12540
rect 4697 12486 4723 12538
rect 4723 12486 4753 12538
rect 4777 12486 4787 12538
rect 4787 12486 4833 12538
rect 4857 12486 4903 12538
rect 4903 12486 4913 12538
rect 4937 12486 4967 12538
rect 4967 12486 4993 12538
rect 4697 12484 4753 12486
rect 4777 12484 4833 12486
rect 4857 12484 4913 12486
rect 4937 12484 4993 12486
rect 5078 11892 5134 11928
rect 5078 11872 5080 11892
rect 5080 11872 5132 11892
rect 5132 11872 5134 11892
rect 5078 11464 5134 11520
rect 4697 11450 4753 11452
rect 4777 11450 4833 11452
rect 4857 11450 4913 11452
rect 4937 11450 4993 11452
rect 4697 11398 4723 11450
rect 4723 11398 4753 11450
rect 4777 11398 4787 11450
rect 4787 11398 4833 11450
rect 4857 11398 4903 11450
rect 4903 11398 4913 11450
rect 4937 11398 4967 11450
rect 4967 11398 4993 11450
rect 4697 11396 4753 11398
rect 4777 11396 4833 11398
rect 4857 11396 4913 11398
rect 4937 11396 4993 11398
rect 4250 10376 4306 10432
rect 3882 8472 3938 8528
rect 3974 7520 4030 7576
rect 3974 6568 4030 6624
rect 3974 6432 4030 6488
rect 4066 6024 4122 6080
rect 4250 9288 4306 9344
rect 4250 6568 4306 6624
rect 4434 10648 4490 10704
rect 4434 10376 4490 10432
rect 4434 9696 4490 9752
rect 4434 7520 4490 7576
rect 3882 3848 3938 3904
rect 3882 2760 3938 2816
rect 4066 4256 4122 4312
rect 4434 4528 4490 4584
rect 4342 3712 4398 3768
rect 4894 10648 4950 10704
rect 4802 10512 4858 10568
rect 4697 10362 4753 10364
rect 4777 10362 4833 10364
rect 4857 10362 4913 10364
rect 4937 10362 4993 10364
rect 4697 10310 4723 10362
rect 4723 10310 4753 10362
rect 4777 10310 4787 10362
rect 4787 10310 4833 10362
rect 4857 10310 4903 10362
rect 4903 10310 4913 10362
rect 4937 10310 4967 10362
rect 4967 10310 4993 10362
rect 4697 10308 4753 10310
rect 4777 10308 4833 10310
rect 4857 10308 4913 10310
rect 4937 10308 4993 10310
rect 4618 9460 4620 9480
rect 4620 9460 4672 9480
rect 4672 9460 4674 9480
rect 4618 9424 4674 9460
rect 4986 9988 5042 10024
rect 4986 9968 4988 9988
rect 4988 9968 5040 9988
rect 5040 9968 5042 9988
rect 4894 9596 4896 9616
rect 4896 9596 4948 9616
rect 4948 9596 4950 9616
rect 4894 9560 4950 9596
rect 4697 9274 4753 9276
rect 4777 9274 4833 9276
rect 4857 9274 4913 9276
rect 4937 9274 4993 9276
rect 4697 9222 4723 9274
rect 4723 9222 4753 9274
rect 4777 9222 4787 9274
rect 4787 9222 4833 9274
rect 4857 9222 4903 9274
rect 4903 9222 4913 9274
rect 4937 9222 4967 9274
rect 4967 9222 4993 9274
rect 4697 9220 4753 9222
rect 4777 9220 4833 9222
rect 4857 9220 4913 9222
rect 4937 9220 4993 9222
rect 6568 13082 6624 13084
rect 6648 13082 6704 13084
rect 6728 13082 6784 13084
rect 6808 13082 6864 13084
rect 6568 13030 6594 13082
rect 6594 13030 6624 13082
rect 6648 13030 6658 13082
rect 6658 13030 6704 13082
rect 6728 13030 6774 13082
rect 6774 13030 6784 13082
rect 6808 13030 6838 13082
rect 6838 13030 6864 13082
rect 6568 13028 6624 13030
rect 6648 13028 6704 13030
rect 6728 13028 6784 13030
rect 6808 13028 6864 13030
rect 5538 12144 5594 12200
rect 5354 10784 5410 10840
rect 5078 8336 5134 8392
rect 4697 8186 4753 8188
rect 4777 8186 4833 8188
rect 4857 8186 4913 8188
rect 4937 8186 4993 8188
rect 4697 8134 4723 8186
rect 4723 8134 4753 8186
rect 4777 8134 4787 8186
rect 4787 8134 4833 8186
rect 4857 8134 4903 8186
rect 4903 8134 4913 8186
rect 4937 8134 4967 8186
rect 4967 8134 4993 8186
rect 4697 8132 4753 8134
rect 4777 8132 4833 8134
rect 4857 8132 4913 8134
rect 4937 8132 4993 8134
rect 4986 7384 5042 7440
rect 4697 7098 4753 7100
rect 4777 7098 4833 7100
rect 4857 7098 4913 7100
rect 4937 7098 4993 7100
rect 4697 7046 4723 7098
rect 4723 7046 4753 7098
rect 4777 7046 4787 7098
rect 4787 7046 4833 7098
rect 4857 7046 4903 7098
rect 4903 7046 4913 7098
rect 4937 7046 4967 7098
rect 4967 7046 4993 7098
rect 4697 7044 4753 7046
rect 4777 7044 4833 7046
rect 4857 7044 4913 7046
rect 4937 7044 4993 7046
rect 5078 6704 5134 6760
rect 4618 6432 4674 6488
rect 5078 6316 5134 6352
rect 5078 6296 5080 6316
rect 5080 6296 5132 6316
rect 5132 6296 5134 6316
rect 4697 6010 4753 6012
rect 4777 6010 4833 6012
rect 4857 6010 4913 6012
rect 4937 6010 4993 6012
rect 4697 5958 4723 6010
rect 4723 5958 4753 6010
rect 4777 5958 4787 6010
rect 4787 5958 4833 6010
rect 4857 5958 4903 6010
rect 4903 5958 4913 6010
rect 4937 5958 4967 6010
rect 4967 5958 4993 6010
rect 4697 5956 4753 5958
rect 4777 5956 4833 5958
rect 4857 5956 4913 5958
rect 4937 5956 4993 5958
rect 4697 4922 4753 4924
rect 4777 4922 4833 4924
rect 4857 4922 4913 4924
rect 4937 4922 4993 4924
rect 4697 4870 4723 4922
rect 4723 4870 4753 4922
rect 4777 4870 4787 4922
rect 4787 4870 4833 4922
rect 4857 4870 4903 4922
rect 4903 4870 4913 4922
rect 4937 4870 4967 4922
rect 4967 4870 4993 4922
rect 4697 4868 4753 4870
rect 4777 4868 4833 4870
rect 4857 4868 4913 4870
rect 4937 4868 4993 4870
rect 4158 2896 4214 2952
rect 3790 2624 3846 2680
rect 3974 2624 4030 2680
rect 4697 3834 4753 3836
rect 4777 3834 4833 3836
rect 4857 3834 4913 3836
rect 4937 3834 4993 3836
rect 4697 3782 4723 3834
rect 4723 3782 4753 3834
rect 4777 3782 4787 3834
rect 4787 3782 4833 3834
rect 4857 3782 4903 3834
rect 4903 3782 4913 3834
rect 4937 3782 4967 3834
rect 4967 3782 4993 3834
rect 4697 3780 4753 3782
rect 4777 3780 4833 3782
rect 4857 3780 4913 3782
rect 4937 3780 4993 3782
rect 4802 3576 4858 3632
rect 4066 1128 4122 1184
rect 4526 3440 4582 3496
rect 6568 11994 6624 11996
rect 6648 11994 6704 11996
rect 6728 11994 6784 11996
rect 6808 11994 6864 11996
rect 6568 11942 6594 11994
rect 6594 11942 6624 11994
rect 6648 11942 6658 11994
rect 6658 11942 6704 11994
rect 6728 11942 6774 11994
rect 6774 11942 6784 11994
rect 6808 11942 6838 11994
rect 6838 11942 6864 11994
rect 6568 11940 6624 11942
rect 6648 11940 6704 11942
rect 6728 11940 6784 11942
rect 6808 11940 6864 11942
rect 5906 11872 5962 11928
rect 5630 11348 5686 11384
rect 5630 11328 5632 11348
rect 5632 11328 5684 11348
rect 5684 11328 5686 11348
rect 5630 11212 5686 11248
rect 5630 11192 5632 11212
rect 5632 11192 5684 11212
rect 5684 11192 5686 11212
rect 5722 11056 5778 11112
rect 5630 9560 5686 9616
rect 5446 9288 5502 9344
rect 5354 7792 5410 7848
rect 5814 9968 5870 10024
rect 5446 6704 5502 6760
rect 5446 6568 5502 6624
rect 5170 5908 5226 5944
rect 5170 5888 5172 5908
rect 5172 5888 5224 5908
rect 5224 5888 5226 5908
rect 5170 3848 5226 3904
rect 4802 2896 4858 2952
rect 4697 2746 4753 2748
rect 4777 2746 4833 2748
rect 4857 2746 4913 2748
rect 4937 2746 4993 2748
rect 4697 2694 4723 2746
rect 4723 2694 4753 2746
rect 4777 2694 4787 2746
rect 4787 2694 4833 2746
rect 4857 2694 4903 2746
rect 4903 2694 4913 2746
rect 4937 2694 4967 2746
rect 4967 2694 4993 2746
rect 4697 2692 4753 2694
rect 4777 2692 4833 2694
rect 4857 2692 4913 2694
rect 4937 2692 4993 2694
rect 5262 3168 5318 3224
rect 4710 2488 4766 2544
rect 4526 1128 4582 1184
rect 5446 5072 5502 5128
rect 5722 6704 5778 6760
rect 5630 5072 5686 5128
rect 5630 3596 5686 3632
rect 5630 3576 5632 3596
rect 5632 3576 5684 3596
rect 5684 3576 5686 3596
rect 5538 3168 5594 3224
rect 5538 3032 5594 3088
rect 5262 1536 5318 1592
rect 5998 9832 6054 9888
rect 6182 11056 6238 11112
rect 6182 9460 6184 9480
rect 6184 9460 6236 9480
rect 6236 9460 6238 9480
rect 6182 9424 6238 9460
rect 6458 11328 6514 11384
rect 6550 11056 6606 11112
rect 6568 10906 6624 10908
rect 6648 10906 6704 10908
rect 6728 10906 6784 10908
rect 6808 10906 6864 10908
rect 6568 10854 6594 10906
rect 6594 10854 6624 10906
rect 6648 10854 6658 10906
rect 6658 10854 6704 10906
rect 6728 10854 6774 10906
rect 6774 10854 6784 10906
rect 6808 10854 6838 10906
rect 6838 10854 6864 10906
rect 6568 10852 6624 10854
rect 6648 10852 6704 10854
rect 6728 10852 6784 10854
rect 6808 10852 6864 10854
rect 6550 10240 6606 10296
rect 7378 11056 7434 11112
rect 6642 9968 6698 10024
rect 6918 9968 6974 10024
rect 6090 8336 6146 8392
rect 6568 9818 6624 9820
rect 6648 9818 6704 9820
rect 6728 9818 6784 9820
rect 6808 9818 6864 9820
rect 6568 9766 6594 9818
rect 6594 9766 6624 9818
rect 6648 9766 6658 9818
rect 6658 9766 6704 9818
rect 6728 9766 6774 9818
rect 6774 9766 6784 9818
rect 6808 9766 6838 9818
rect 6838 9766 6864 9818
rect 6568 9764 6624 9766
rect 6648 9764 6704 9766
rect 6728 9764 6784 9766
rect 6808 9764 6864 9766
rect 7654 11056 7710 11112
rect 7470 10104 7526 10160
rect 7194 9424 7250 9480
rect 6568 8730 6624 8732
rect 6648 8730 6704 8732
rect 6728 8730 6784 8732
rect 6808 8730 6864 8732
rect 6568 8678 6594 8730
rect 6594 8678 6624 8730
rect 6648 8678 6658 8730
rect 6658 8678 6704 8730
rect 6728 8678 6774 8730
rect 6774 8678 6784 8730
rect 6808 8678 6838 8730
rect 6838 8678 6864 8730
rect 6568 8676 6624 8678
rect 6648 8676 6704 8678
rect 6728 8676 6784 8678
rect 6808 8676 6864 8678
rect 5722 2644 5778 2680
rect 5722 2624 5724 2644
rect 5724 2624 5776 2644
rect 5776 2624 5778 2644
rect 5630 2352 5686 2408
rect 5538 1264 5594 1320
rect 5998 5344 6054 5400
rect 5906 4800 5962 4856
rect 6568 7642 6624 7644
rect 6648 7642 6704 7644
rect 6728 7642 6784 7644
rect 6808 7642 6864 7644
rect 6568 7590 6594 7642
rect 6594 7590 6624 7642
rect 6648 7590 6658 7642
rect 6658 7590 6704 7642
rect 6728 7590 6774 7642
rect 6774 7590 6784 7642
rect 6808 7590 6838 7642
rect 6838 7590 6864 7642
rect 6568 7588 6624 7590
rect 6648 7588 6704 7590
rect 6728 7588 6784 7590
rect 6808 7588 6864 7590
rect 6458 7268 6514 7304
rect 6458 7248 6460 7268
rect 6460 7248 6512 7268
rect 6512 7248 6514 7268
rect 6568 6554 6624 6556
rect 6648 6554 6704 6556
rect 6728 6554 6784 6556
rect 6808 6554 6864 6556
rect 6568 6502 6594 6554
rect 6594 6502 6624 6554
rect 6648 6502 6658 6554
rect 6658 6502 6704 6554
rect 6728 6502 6774 6554
rect 6774 6502 6784 6554
rect 6808 6502 6838 6554
rect 6838 6502 6864 6554
rect 6568 6500 6624 6502
rect 6648 6500 6704 6502
rect 6728 6500 6784 6502
rect 6808 6500 6864 6502
rect 6568 5466 6624 5468
rect 6648 5466 6704 5468
rect 6728 5466 6784 5468
rect 6808 5466 6864 5468
rect 6568 5414 6594 5466
rect 6594 5414 6624 5466
rect 6648 5414 6658 5466
rect 6658 5414 6704 5466
rect 6728 5414 6774 5466
rect 6774 5414 6784 5466
rect 6808 5414 6838 5466
rect 6838 5414 6864 5466
rect 6568 5412 6624 5414
rect 6648 5412 6704 5414
rect 6728 5412 6784 5414
rect 6808 5412 6864 5414
rect 6182 4664 6238 4720
rect 6366 4664 6422 4720
rect 6090 4392 6146 4448
rect 5998 4120 6054 4176
rect 5998 3848 6054 3904
rect 6274 4528 6330 4584
rect 6918 4528 6974 4584
rect 6568 4378 6624 4380
rect 6648 4378 6704 4380
rect 6728 4378 6784 4380
rect 6808 4378 6864 4380
rect 6568 4326 6594 4378
rect 6594 4326 6624 4378
rect 6648 4326 6658 4378
rect 6658 4326 6704 4378
rect 6728 4326 6774 4378
rect 6774 4326 6784 4378
rect 6808 4326 6838 4378
rect 6838 4326 6864 4378
rect 6568 4324 6624 4326
rect 6648 4324 6704 4326
rect 6728 4324 6784 4326
rect 6808 4324 6864 4326
rect 6274 3712 6330 3768
rect 6918 3848 6974 3904
rect 6182 3440 6238 3496
rect 6918 3576 6974 3632
rect 6568 3290 6624 3292
rect 6648 3290 6704 3292
rect 6728 3290 6784 3292
rect 6808 3290 6864 3292
rect 6568 3238 6594 3290
rect 6594 3238 6624 3290
rect 6648 3238 6658 3290
rect 6658 3238 6704 3290
rect 6728 3238 6774 3290
rect 6774 3238 6784 3290
rect 6808 3238 6838 3290
rect 6838 3238 6864 3290
rect 6568 3236 6624 3238
rect 6648 3236 6704 3238
rect 6728 3236 6784 3238
rect 6808 3236 6864 3238
rect 6458 3032 6514 3088
rect 6642 3032 6698 3088
rect 5998 1672 6054 1728
rect 5906 992 5962 1048
rect 6826 2896 6882 2952
rect 7194 6296 7250 6352
rect 7102 6024 7158 6080
rect 6568 2202 6624 2204
rect 6648 2202 6704 2204
rect 6728 2202 6784 2204
rect 6808 2202 6864 2204
rect 6568 2150 6594 2202
rect 6594 2150 6624 2202
rect 6648 2150 6658 2202
rect 6658 2150 6704 2202
rect 6728 2150 6774 2202
rect 6774 2150 6784 2202
rect 6808 2150 6838 2202
rect 6838 2150 6864 2202
rect 6568 2148 6624 2150
rect 6648 2148 6704 2150
rect 6728 2148 6784 2150
rect 6808 2148 6864 2150
rect 6366 1808 6422 1864
rect 6734 1944 6790 2000
rect 7562 8336 7618 8392
rect 8438 12538 8494 12540
rect 8518 12538 8574 12540
rect 8598 12538 8654 12540
rect 8678 12538 8734 12540
rect 8438 12486 8464 12538
rect 8464 12486 8494 12538
rect 8518 12486 8528 12538
rect 8528 12486 8574 12538
rect 8598 12486 8644 12538
rect 8644 12486 8654 12538
rect 8678 12486 8708 12538
rect 8708 12486 8734 12538
rect 8438 12484 8494 12486
rect 8518 12484 8574 12486
rect 8598 12484 8654 12486
rect 8678 12484 8734 12486
rect 8114 11464 8170 11520
rect 8438 11450 8494 11452
rect 8518 11450 8574 11452
rect 8598 11450 8654 11452
rect 8678 11450 8734 11452
rect 8438 11398 8464 11450
rect 8464 11398 8494 11450
rect 8518 11398 8528 11450
rect 8528 11398 8574 11450
rect 8598 11398 8644 11450
rect 8644 11398 8654 11450
rect 8678 11398 8708 11450
rect 8708 11398 8734 11450
rect 8438 11396 8494 11398
rect 8518 11396 8574 11398
rect 8598 11396 8654 11398
rect 8678 11396 8734 11398
rect 10309 13082 10365 13084
rect 10389 13082 10445 13084
rect 10469 13082 10525 13084
rect 10549 13082 10605 13084
rect 10309 13030 10335 13082
rect 10335 13030 10365 13082
rect 10389 13030 10399 13082
rect 10399 13030 10445 13082
rect 10469 13030 10515 13082
rect 10515 13030 10525 13082
rect 10549 13030 10579 13082
rect 10579 13030 10605 13082
rect 10309 13028 10365 13030
rect 10389 13028 10445 13030
rect 10469 13028 10525 13030
rect 10549 13028 10605 13030
rect 7838 10512 7894 10568
rect 7562 5344 7618 5400
rect 7654 4528 7710 4584
rect 7378 3984 7434 4040
rect 7838 4800 7894 4856
rect 7562 2760 7618 2816
rect 7838 2488 7894 2544
rect 8114 3984 8170 4040
rect 8114 2896 8170 2952
rect 8438 10362 8494 10364
rect 8518 10362 8574 10364
rect 8598 10362 8654 10364
rect 8678 10362 8734 10364
rect 8438 10310 8464 10362
rect 8464 10310 8494 10362
rect 8518 10310 8528 10362
rect 8528 10310 8574 10362
rect 8598 10310 8644 10362
rect 8644 10310 8654 10362
rect 8678 10310 8708 10362
rect 8708 10310 8734 10362
rect 8438 10308 8494 10310
rect 8518 10308 8574 10310
rect 8598 10308 8654 10310
rect 8678 10308 8734 10310
rect 8438 9274 8494 9276
rect 8518 9274 8574 9276
rect 8598 9274 8654 9276
rect 8678 9274 8734 9276
rect 8438 9222 8464 9274
rect 8464 9222 8494 9274
rect 8518 9222 8528 9274
rect 8528 9222 8574 9274
rect 8598 9222 8644 9274
rect 8644 9222 8654 9274
rect 8678 9222 8708 9274
rect 8708 9222 8734 9274
rect 8438 9220 8494 9222
rect 8518 9220 8574 9222
rect 8598 9220 8654 9222
rect 8678 9220 8734 9222
rect 8438 8186 8494 8188
rect 8518 8186 8574 8188
rect 8598 8186 8654 8188
rect 8678 8186 8734 8188
rect 8438 8134 8464 8186
rect 8464 8134 8494 8186
rect 8518 8134 8528 8186
rect 8528 8134 8574 8186
rect 8598 8134 8644 8186
rect 8644 8134 8654 8186
rect 8678 8134 8708 8186
rect 8708 8134 8734 8186
rect 8438 8132 8494 8134
rect 8518 8132 8574 8134
rect 8598 8132 8654 8134
rect 8678 8132 8734 8134
rect 8298 7928 8354 7984
rect 8438 7098 8494 7100
rect 8518 7098 8574 7100
rect 8598 7098 8654 7100
rect 8678 7098 8734 7100
rect 8438 7046 8464 7098
rect 8464 7046 8494 7098
rect 8518 7046 8528 7098
rect 8528 7046 8574 7098
rect 8598 7046 8644 7098
rect 8644 7046 8654 7098
rect 8678 7046 8708 7098
rect 8708 7046 8734 7098
rect 8438 7044 8494 7046
rect 8518 7044 8574 7046
rect 8598 7044 8654 7046
rect 8678 7044 8734 7046
rect 8850 7928 8906 7984
rect 8482 6316 8538 6352
rect 8482 6296 8484 6316
rect 8484 6296 8536 6316
rect 8536 6296 8538 6316
rect 8438 6010 8494 6012
rect 8518 6010 8574 6012
rect 8598 6010 8654 6012
rect 8678 6010 8734 6012
rect 8438 5958 8464 6010
rect 8464 5958 8494 6010
rect 8518 5958 8528 6010
rect 8528 5958 8574 6010
rect 8598 5958 8644 6010
rect 8644 5958 8654 6010
rect 8678 5958 8708 6010
rect 8708 5958 8734 6010
rect 8438 5956 8494 5958
rect 8518 5956 8574 5958
rect 8598 5956 8654 5958
rect 8678 5956 8734 5958
rect 8574 5480 8630 5536
rect 8438 4922 8494 4924
rect 8518 4922 8574 4924
rect 8598 4922 8654 4924
rect 8678 4922 8734 4924
rect 8438 4870 8464 4922
rect 8464 4870 8494 4922
rect 8518 4870 8528 4922
rect 8528 4870 8574 4922
rect 8598 4870 8644 4922
rect 8644 4870 8654 4922
rect 8678 4870 8708 4922
rect 8708 4870 8734 4922
rect 8438 4868 8494 4870
rect 8518 4868 8574 4870
rect 8598 4868 8654 4870
rect 8678 4868 8734 4870
rect 8298 3848 8354 3904
rect 8438 3834 8494 3836
rect 8518 3834 8574 3836
rect 8598 3834 8654 3836
rect 8678 3834 8734 3836
rect 8438 3782 8464 3834
rect 8464 3782 8494 3834
rect 8518 3782 8528 3834
rect 8528 3782 8574 3834
rect 8598 3782 8644 3834
rect 8644 3782 8654 3834
rect 8678 3782 8708 3834
rect 8708 3782 8734 3834
rect 8438 3780 8494 3782
rect 8518 3780 8574 3782
rect 8598 3780 8654 3782
rect 8678 3780 8734 3782
rect 8758 3596 8814 3632
rect 8758 3576 8760 3596
rect 8760 3576 8812 3596
rect 8812 3576 8814 3596
rect 8666 3440 8722 3496
rect 8758 3168 8814 3224
rect 8482 3032 8538 3088
rect 8438 2746 8494 2748
rect 8518 2746 8574 2748
rect 8598 2746 8654 2748
rect 8678 2746 8734 2748
rect 8438 2694 8464 2746
rect 8464 2694 8494 2746
rect 8518 2694 8528 2746
rect 8528 2694 8574 2746
rect 8598 2694 8644 2746
rect 8644 2694 8654 2746
rect 8678 2694 8708 2746
rect 8708 2694 8734 2746
rect 8438 2692 8494 2694
rect 8518 2692 8574 2694
rect 8598 2692 8654 2694
rect 8678 2692 8734 2694
rect 8482 2488 8538 2544
rect 8666 2508 8722 2544
rect 8666 2488 8668 2508
rect 8668 2488 8720 2508
rect 8720 2488 8722 2508
rect 8390 2352 8446 2408
rect 8666 2216 8722 2272
rect 8758 1672 8814 1728
rect 8942 5208 8998 5264
rect 8850 1264 8906 1320
rect 9126 5228 9182 5264
rect 9126 5208 9128 5228
rect 9128 5208 9180 5228
rect 9180 5208 9182 5228
rect 9770 12144 9826 12200
rect 10309 11994 10365 11996
rect 10389 11994 10445 11996
rect 10469 11994 10525 11996
rect 10549 11994 10605 11996
rect 10309 11942 10335 11994
rect 10335 11942 10365 11994
rect 10389 11942 10399 11994
rect 10399 11942 10445 11994
rect 10469 11942 10515 11994
rect 10515 11942 10525 11994
rect 10549 11942 10579 11994
rect 10579 11942 10605 11994
rect 10309 11940 10365 11942
rect 10389 11940 10445 11942
rect 10469 11940 10525 11942
rect 10549 11940 10605 11942
rect 10414 11636 10416 11656
rect 10416 11636 10468 11656
rect 10468 11636 10470 11656
rect 10414 11600 10470 11636
rect 9770 11192 9826 11248
rect 9678 11056 9734 11112
rect 10046 11192 10102 11248
rect 11242 12144 11298 12200
rect 10322 11056 10378 11112
rect 10309 10906 10365 10908
rect 10389 10906 10445 10908
rect 10469 10906 10525 10908
rect 10549 10906 10605 10908
rect 10309 10854 10335 10906
rect 10335 10854 10365 10906
rect 10389 10854 10399 10906
rect 10399 10854 10445 10906
rect 10469 10854 10515 10906
rect 10515 10854 10525 10906
rect 10549 10854 10579 10906
rect 10579 10854 10605 10906
rect 10309 10852 10365 10854
rect 10389 10852 10445 10854
rect 10469 10852 10525 10854
rect 10549 10852 10605 10854
rect 10309 9818 10365 9820
rect 10389 9818 10445 9820
rect 10469 9818 10525 9820
rect 10549 9818 10605 9820
rect 10309 9766 10335 9818
rect 10335 9766 10365 9818
rect 10389 9766 10399 9818
rect 10399 9766 10445 9818
rect 10469 9766 10515 9818
rect 10515 9766 10525 9818
rect 10549 9766 10579 9818
rect 10579 9766 10605 9818
rect 10309 9764 10365 9766
rect 10389 9764 10445 9766
rect 10469 9764 10525 9766
rect 10549 9764 10605 9766
rect 9678 7384 9734 7440
rect 9586 5344 9642 5400
rect 9494 4820 9550 4856
rect 9494 4800 9496 4820
rect 9496 4800 9548 4820
rect 9548 4800 9550 4820
rect 9402 3984 9458 4040
rect 9678 5208 9734 5264
rect 9678 4564 9680 4584
rect 9680 4564 9732 4584
rect 9732 4564 9734 4584
rect 9678 4528 9734 4564
rect 9954 7792 10010 7848
rect 9862 7656 9918 7712
rect 9862 6316 9918 6352
rect 9862 6296 9864 6316
rect 9864 6296 9916 6316
rect 9916 6296 9918 6316
rect 10046 5480 10102 5536
rect 9678 3576 9734 3632
rect 9862 2508 9918 2544
rect 9862 2488 9864 2508
rect 9864 2488 9916 2508
rect 9916 2488 9918 2508
rect 10309 8730 10365 8732
rect 10389 8730 10445 8732
rect 10469 8730 10525 8732
rect 10549 8730 10605 8732
rect 10309 8678 10335 8730
rect 10335 8678 10365 8730
rect 10389 8678 10399 8730
rect 10399 8678 10445 8730
rect 10469 8678 10515 8730
rect 10515 8678 10525 8730
rect 10549 8678 10579 8730
rect 10579 8678 10605 8730
rect 10309 8676 10365 8678
rect 10389 8676 10445 8678
rect 10469 8676 10525 8678
rect 10549 8676 10605 8678
rect 10309 7642 10365 7644
rect 10389 7642 10445 7644
rect 10469 7642 10525 7644
rect 10549 7642 10605 7644
rect 10309 7590 10335 7642
rect 10335 7590 10365 7642
rect 10389 7590 10399 7642
rect 10399 7590 10445 7642
rect 10469 7590 10515 7642
rect 10515 7590 10525 7642
rect 10549 7590 10579 7642
rect 10579 7590 10605 7642
rect 10309 7588 10365 7590
rect 10389 7588 10445 7590
rect 10469 7588 10525 7590
rect 10549 7588 10605 7590
rect 10322 7420 10324 7440
rect 10324 7420 10376 7440
rect 10376 7420 10378 7440
rect 11242 11600 11298 11656
rect 10966 7928 11022 7984
rect 10322 7384 10378 7420
rect 10506 6996 10562 7032
rect 10506 6976 10508 6996
rect 10508 6976 10560 6996
rect 10560 6976 10562 6996
rect 10309 6554 10365 6556
rect 10389 6554 10445 6556
rect 10469 6554 10525 6556
rect 10549 6554 10605 6556
rect 10309 6502 10335 6554
rect 10335 6502 10365 6554
rect 10389 6502 10399 6554
rect 10399 6502 10445 6554
rect 10469 6502 10515 6554
rect 10515 6502 10525 6554
rect 10549 6502 10579 6554
rect 10579 6502 10605 6554
rect 10309 6500 10365 6502
rect 10389 6500 10445 6502
rect 10469 6500 10525 6502
rect 10549 6500 10605 6502
rect 10230 5616 10286 5672
rect 10309 5466 10365 5468
rect 10389 5466 10445 5468
rect 10469 5466 10525 5468
rect 10549 5466 10605 5468
rect 10309 5414 10335 5466
rect 10335 5414 10365 5466
rect 10389 5414 10399 5466
rect 10399 5414 10445 5466
rect 10469 5414 10515 5466
rect 10515 5414 10525 5466
rect 10549 5414 10579 5466
rect 10579 5414 10605 5466
rect 10309 5412 10365 5414
rect 10389 5412 10445 5414
rect 10469 5412 10525 5414
rect 10549 5412 10605 5414
rect 10598 5072 10654 5128
rect 10046 3032 10102 3088
rect 10309 4378 10365 4380
rect 10389 4378 10445 4380
rect 10469 4378 10525 4380
rect 10549 4378 10605 4380
rect 10309 4326 10335 4378
rect 10335 4326 10365 4378
rect 10389 4326 10399 4378
rect 10399 4326 10445 4378
rect 10469 4326 10515 4378
rect 10515 4326 10525 4378
rect 10549 4326 10579 4378
rect 10579 4326 10605 4378
rect 10309 4324 10365 4326
rect 10389 4324 10445 4326
rect 10469 4324 10525 4326
rect 10549 4324 10605 4326
rect 10309 3290 10365 3292
rect 10389 3290 10445 3292
rect 10469 3290 10525 3292
rect 10549 3290 10605 3292
rect 10309 3238 10335 3290
rect 10335 3238 10365 3290
rect 10389 3238 10399 3290
rect 10399 3238 10445 3290
rect 10469 3238 10515 3290
rect 10515 3238 10525 3290
rect 10549 3238 10579 3290
rect 10579 3238 10605 3290
rect 10309 3236 10365 3238
rect 10389 3236 10445 3238
rect 10469 3236 10525 3238
rect 10549 3236 10605 3238
rect 10322 2508 10378 2544
rect 10966 4564 10968 4584
rect 10968 4564 11020 4584
rect 11020 4564 11022 4584
rect 10966 4528 11022 4564
rect 11058 3460 11114 3496
rect 11058 3440 11060 3460
rect 11060 3440 11112 3460
rect 11112 3440 11114 3460
rect 10322 2488 10324 2508
rect 10324 2488 10376 2508
rect 10376 2488 10378 2508
rect 10230 2352 10286 2408
rect 10782 2352 10838 2408
rect 10309 2202 10365 2204
rect 10389 2202 10445 2204
rect 10469 2202 10525 2204
rect 10549 2202 10605 2204
rect 10309 2150 10335 2202
rect 10335 2150 10365 2202
rect 10389 2150 10399 2202
rect 10399 2150 10445 2202
rect 10469 2150 10515 2202
rect 10515 2150 10525 2202
rect 10549 2150 10579 2202
rect 10579 2150 10605 2202
rect 10309 2148 10365 2150
rect 10389 2148 10445 2150
rect 10469 2148 10525 2150
rect 10549 2148 10605 2150
rect 12438 2488 12494 2544
rect 13174 3576 13230 3632
<< metal3 >>
rect 2814 13088 3134 13089
rect 2814 13024 2822 13088
rect 2886 13024 2902 13088
rect 2966 13024 2982 13088
rect 3046 13024 3062 13088
rect 3126 13024 3134 13088
rect 2814 13023 3134 13024
rect 6556 13088 6876 13089
rect 6556 13024 6564 13088
rect 6628 13024 6644 13088
rect 6708 13024 6724 13088
rect 6788 13024 6804 13088
rect 6868 13024 6876 13088
rect 6556 13023 6876 13024
rect 10297 13088 10617 13089
rect 10297 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10465 13088
rect 10529 13024 10545 13088
rect 10609 13024 10617 13088
rect 10297 13023 10617 13024
rect 1853 12610 1919 12613
rect 2405 12612 2471 12613
rect 2078 12610 2084 12612
rect 1853 12608 2084 12610
rect 1853 12552 1858 12608
rect 1914 12552 2084 12608
rect 1853 12550 2084 12552
rect 1853 12547 1919 12550
rect 2078 12548 2084 12550
rect 2148 12548 2154 12612
rect 2405 12610 2452 12612
rect 2360 12608 2452 12610
rect 2360 12552 2410 12608
rect 2360 12550 2452 12552
rect 2405 12548 2452 12550
rect 2516 12548 2522 12612
rect 2405 12547 2471 12548
rect 4685 12544 5005 12545
rect 4685 12480 4693 12544
rect 4757 12480 4773 12544
rect 4837 12480 4853 12544
rect 4917 12480 4933 12544
rect 4997 12480 5005 12544
rect 4685 12479 5005 12480
rect 8426 12544 8746 12545
rect 8426 12480 8434 12544
rect 8498 12480 8514 12544
rect 8578 12480 8594 12544
rect 8658 12480 8674 12544
rect 8738 12480 8746 12544
rect 8426 12479 8746 12480
rect 565 12474 631 12477
rect 4153 12474 4219 12477
rect 565 12472 4219 12474
rect 565 12416 570 12472
rect 626 12416 4158 12472
rect 4214 12416 4219 12472
rect 565 12414 4219 12416
rect 565 12411 631 12414
rect 4153 12411 4219 12414
rect 1301 12202 1367 12205
rect 5533 12202 5599 12205
rect 1301 12200 5599 12202
rect 1301 12144 1306 12200
rect 1362 12144 5538 12200
rect 5594 12144 5599 12200
rect 1301 12142 5599 12144
rect 1301 12139 1367 12142
rect 5533 12139 5599 12142
rect 9765 12202 9831 12205
rect 11237 12202 11303 12205
rect 9765 12200 11303 12202
rect 9765 12144 9770 12200
rect 9826 12144 11242 12200
rect 11298 12144 11303 12200
rect 9765 12142 11303 12144
rect 9765 12139 9831 12142
rect 11237 12139 11303 12142
rect 2814 12000 3134 12001
rect 2814 11936 2822 12000
rect 2886 11936 2902 12000
rect 2966 11936 2982 12000
rect 3046 11936 3062 12000
rect 3126 11936 3134 12000
rect 2814 11935 3134 11936
rect 6556 12000 6876 12001
rect 6556 11936 6564 12000
rect 6628 11936 6644 12000
rect 6708 11936 6724 12000
rect 6788 11936 6804 12000
rect 6868 11936 6876 12000
rect 6556 11935 6876 11936
rect 10297 12000 10617 12001
rect 10297 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10545 12000
rect 10609 11936 10617 12000
rect 10297 11935 10617 11936
rect 5073 11930 5139 11933
rect 5901 11930 5967 11933
rect 5073 11928 5967 11930
rect 5073 11872 5078 11928
rect 5134 11872 5906 11928
rect 5962 11872 5967 11928
rect 5073 11870 5967 11872
rect 5073 11867 5139 11870
rect 5901 11867 5967 11870
rect 10409 11658 10475 11661
rect 11237 11658 11303 11661
rect 10409 11656 11303 11658
rect 10409 11600 10414 11656
rect 10470 11600 11242 11656
rect 11298 11600 11303 11656
rect 10409 11598 11303 11600
rect 10409 11595 10475 11598
rect 11237 11595 11303 11598
rect 5073 11522 5139 11525
rect 8109 11522 8175 11525
rect 5073 11520 8175 11522
rect 5073 11464 5078 11520
rect 5134 11464 8114 11520
rect 8170 11464 8175 11520
rect 5073 11462 8175 11464
rect 5073 11459 5139 11462
rect 8109 11459 8175 11462
rect 4685 11456 5005 11457
rect 4685 11392 4693 11456
rect 4757 11392 4773 11456
rect 4837 11392 4853 11456
rect 4917 11392 4933 11456
rect 4997 11392 5005 11456
rect 4685 11391 5005 11392
rect 8426 11456 8746 11457
rect 8426 11392 8434 11456
rect 8498 11392 8514 11456
rect 8578 11392 8594 11456
rect 8658 11392 8674 11456
rect 8738 11392 8746 11456
rect 8426 11391 8746 11392
rect 5625 11386 5691 11389
rect 6453 11386 6519 11389
rect 5625 11384 6519 11386
rect 5625 11328 5630 11384
rect 5686 11328 6458 11384
rect 6514 11328 6519 11384
rect 5625 11326 6519 11328
rect 5625 11323 5691 11326
rect 6453 11323 6519 11326
rect 5625 11252 5691 11253
rect 5574 11250 5580 11252
rect 5534 11190 5580 11250
rect 5644 11248 5691 11252
rect 5686 11192 5691 11248
rect 5574 11188 5580 11190
rect 5644 11188 5691 11192
rect 5625 11187 5691 11188
rect 9765 11250 9831 11253
rect 10041 11250 10107 11253
rect 9765 11248 10107 11250
rect 9765 11192 9770 11248
rect 9826 11192 10046 11248
rect 10102 11192 10107 11248
rect 9765 11190 10107 11192
rect 9765 11187 9831 11190
rect 10041 11187 10107 11190
rect 974 11052 980 11116
rect 1044 11114 1050 11116
rect 2681 11114 2747 11117
rect 1044 11112 2747 11114
rect 1044 11056 2686 11112
rect 2742 11056 2747 11112
rect 1044 11054 2747 11056
rect 1044 11052 1050 11054
rect 2681 11051 2747 11054
rect 5717 11116 5783 11117
rect 5717 11112 5764 11116
rect 5828 11114 5834 11116
rect 6177 11114 6243 11117
rect 6545 11114 6611 11117
rect 5717 11056 5722 11112
rect 5717 11052 5764 11056
rect 5828 11054 5874 11114
rect 6177 11112 6611 11114
rect 6177 11056 6182 11112
rect 6238 11056 6550 11112
rect 6606 11056 6611 11112
rect 6177 11054 6611 11056
rect 5828 11052 5834 11054
rect 5717 11051 5783 11052
rect 6177 11051 6243 11054
rect 6545 11051 6611 11054
rect 7046 11052 7052 11116
rect 7116 11114 7122 11116
rect 7373 11114 7439 11117
rect 7649 11116 7715 11117
rect 7598 11114 7604 11116
rect 7116 11112 7439 11114
rect 7116 11056 7378 11112
rect 7434 11056 7439 11112
rect 7116 11054 7439 11056
rect 7558 11054 7604 11114
rect 7668 11112 7715 11116
rect 7710 11056 7715 11112
rect 7116 11052 7122 11054
rect 7373 11051 7439 11054
rect 7598 11052 7604 11054
rect 7668 11052 7715 11056
rect 7649 11051 7715 11052
rect 9673 11114 9739 11117
rect 10317 11114 10383 11117
rect 9673 11112 10383 11114
rect 9673 11056 9678 11112
rect 9734 11056 10322 11112
rect 10378 11056 10383 11112
rect 9673 11054 10383 11056
rect 9673 11051 9739 11054
rect 10317 11051 10383 11054
rect 2814 10912 3134 10913
rect 2814 10848 2822 10912
rect 2886 10848 2902 10912
rect 2966 10848 2982 10912
rect 3046 10848 3062 10912
rect 3126 10848 3134 10912
rect 2814 10847 3134 10848
rect 6556 10912 6876 10913
rect 6556 10848 6564 10912
rect 6628 10848 6644 10912
rect 6708 10848 6724 10912
rect 6788 10848 6804 10912
rect 6868 10848 6876 10912
rect 6556 10847 6876 10848
rect 10297 10912 10617 10913
rect 10297 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10545 10912
rect 10609 10848 10617 10912
rect 10297 10847 10617 10848
rect 5349 10844 5415 10845
rect 5206 10842 5212 10844
rect 4662 10782 5212 10842
rect 2221 10706 2287 10709
rect 4429 10706 4495 10709
rect 2221 10704 4495 10706
rect 2221 10648 2226 10704
rect 2282 10648 4434 10704
rect 4490 10648 4495 10704
rect 2221 10646 4495 10648
rect 2221 10643 2287 10646
rect 4429 10643 4495 10646
rect 4662 10570 4722 10782
rect 5206 10780 5212 10782
rect 5276 10780 5282 10844
rect 5349 10840 5396 10844
rect 5460 10842 5466 10844
rect 5349 10784 5354 10840
rect 5349 10780 5396 10784
rect 5460 10782 5506 10842
rect 5460 10780 5466 10782
rect 5349 10779 5415 10780
rect 4889 10706 4955 10709
rect 7966 10706 7972 10708
rect 4889 10704 7972 10706
rect 4889 10648 4894 10704
rect 4950 10648 7972 10704
rect 4889 10646 7972 10648
rect 4889 10643 4955 10646
rect 7966 10644 7972 10646
rect 8036 10644 8042 10708
rect 4432 10510 4722 10570
rect 4797 10570 4863 10573
rect 7833 10570 7899 10573
rect 4797 10568 7899 10570
rect 4797 10512 4802 10568
rect 4858 10512 7838 10568
rect 7894 10512 7899 10568
rect 4797 10510 7899 10512
rect 4432 10437 4492 10510
rect 4797 10507 4863 10510
rect 7833 10507 7899 10510
rect 2865 10432 2931 10437
rect 2865 10376 2870 10432
rect 2926 10376 2931 10432
rect 2865 10371 2931 10376
rect 3233 10434 3299 10437
rect 4245 10434 4311 10437
rect 3233 10432 4311 10434
rect 3233 10376 3238 10432
rect 3294 10376 4250 10432
rect 4306 10376 4311 10432
rect 3233 10374 4311 10376
rect 3233 10371 3299 10374
rect 4245 10371 4311 10374
rect 4429 10432 4495 10437
rect 4429 10376 4434 10432
rect 4490 10376 4495 10432
rect 4429 10371 4495 10376
rect 2868 10298 2928 10371
rect 4685 10368 5005 10369
rect 4685 10304 4693 10368
rect 4757 10304 4773 10368
rect 4837 10304 4853 10368
rect 4917 10304 4933 10368
rect 4997 10304 5005 10368
rect 4685 10303 5005 10304
rect 8426 10368 8746 10369
rect 8426 10304 8434 10368
rect 8498 10304 8514 10368
rect 8578 10304 8594 10368
rect 8658 10304 8674 10368
rect 8738 10304 8746 10368
rect 8426 10303 8746 10304
rect 2868 10238 4354 10298
rect 3417 10162 3483 10165
rect 3785 10162 3851 10165
rect 4294 10162 4354 10238
rect 5206 10236 5212 10300
rect 5276 10298 5282 10300
rect 6545 10298 6611 10301
rect 5276 10296 6611 10298
rect 5276 10240 6550 10296
rect 6606 10240 6611 10296
rect 5276 10238 6611 10240
rect 5276 10236 5282 10238
rect 6545 10235 6611 10238
rect 7465 10162 7531 10165
rect 3417 10160 4170 10162
rect 3417 10104 3422 10160
rect 3478 10104 3790 10160
rect 3846 10104 4170 10160
rect 3417 10102 4170 10104
rect 4294 10160 7531 10162
rect 4294 10104 7470 10160
rect 7526 10104 7531 10160
rect 4294 10102 7531 10104
rect 3417 10099 3483 10102
rect 3785 10099 3851 10102
rect 1945 10026 2011 10029
rect 4110 10026 4170 10102
rect 7465 10099 7531 10102
rect 4981 10026 5047 10029
rect 1945 10024 3434 10026
rect 1945 9968 1950 10024
rect 2006 9968 3434 10024
rect 1945 9966 3434 9968
rect 4110 10024 5047 10026
rect 4110 9968 4986 10024
rect 5042 9968 5047 10024
rect 4110 9966 5047 9968
rect 1945 9963 2011 9966
rect 3374 9890 3434 9966
rect 4981 9963 5047 9966
rect 5809 10026 5875 10029
rect 6637 10026 6703 10029
rect 5809 10024 6703 10026
rect 5809 9968 5814 10024
rect 5870 9968 6642 10024
rect 6698 9968 6703 10024
rect 5809 9966 6703 9968
rect 5809 9963 5875 9966
rect 6637 9963 6703 9966
rect 6913 10026 6979 10029
rect 7230 10026 7236 10028
rect 6913 10024 7236 10026
rect 6913 9968 6918 10024
rect 6974 9968 7236 10024
rect 6913 9966 7236 9968
rect 6913 9963 6979 9966
rect 7230 9964 7236 9966
rect 7300 9964 7306 10028
rect 5993 9890 6059 9893
rect 3374 9888 6059 9890
rect 3374 9832 5998 9888
rect 6054 9832 6059 9888
rect 3374 9830 6059 9832
rect 5993 9827 6059 9830
rect 2814 9824 3134 9825
rect 2814 9760 2822 9824
rect 2886 9760 2902 9824
rect 2966 9760 2982 9824
rect 3046 9760 3062 9824
rect 3126 9760 3134 9824
rect 2814 9759 3134 9760
rect 6556 9824 6876 9825
rect 6556 9760 6564 9824
rect 6628 9760 6644 9824
rect 6708 9760 6724 9824
rect 6788 9760 6804 9824
rect 6868 9760 6876 9824
rect 6556 9759 6876 9760
rect 10297 9824 10617 9825
rect 10297 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10545 9824
rect 10609 9760 10617 9824
rect 10297 9759 10617 9760
rect 4429 9754 4495 9757
rect 6310 9754 6316 9756
rect 4429 9752 6316 9754
rect 4429 9696 4434 9752
rect 4490 9696 6316 9752
rect 4429 9694 6316 9696
rect 4429 9691 4495 9694
rect 6310 9692 6316 9694
rect 6380 9692 6386 9756
rect 3366 9556 3372 9620
rect 3436 9618 3442 9620
rect 4889 9618 4955 9621
rect 3436 9616 4955 9618
rect 3436 9560 4894 9616
rect 4950 9560 4955 9616
rect 3436 9558 4955 9560
rect 3436 9556 3442 9558
rect 4889 9555 4955 9558
rect 5625 9618 5691 9621
rect 9622 9618 9628 9620
rect 5625 9616 9628 9618
rect 5625 9560 5630 9616
rect 5686 9560 9628 9616
rect 5625 9558 9628 9560
rect 5625 9555 5691 9558
rect 9622 9556 9628 9558
rect 9692 9556 9698 9620
rect 3509 9482 3575 9485
rect 4470 9482 4476 9484
rect 3509 9480 4476 9482
rect 3509 9424 3514 9480
rect 3570 9424 4476 9480
rect 3509 9422 4476 9424
rect 3509 9419 3575 9422
rect 4470 9420 4476 9422
rect 4540 9420 4546 9484
rect 4613 9482 4679 9485
rect 6177 9482 6243 9485
rect 7189 9482 7255 9485
rect 4613 9480 5458 9482
rect 4613 9424 4618 9480
rect 4674 9424 5458 9480
rect 4613 9422 5458 9424
rect 4613 9419 4679 9422
rect 5398 9349 5458 9422
rect 6177 9480 7255 9482
rect 6177 9424 6182 9480
rect 6238 9424 7194 9480
rect 7250 9424 7255 9480
rect 6177 9422 7255 9424
rect 6177 9419 6243 9422
rect 7189 9419 7255 9422
rect 4245 9348 4311 9349
rect 4245 9344 4292 9348
rect 4356 9346 4362 9348
rect 4245 9288 4250 9344
rect 4245 9284 4292 9288
rect 4356 9286 4402 9346
rect 5398 9344 5507 9349
rect 5398 9288 5446 9344
rect 5502 9288 5507 9344
rect 5398 9286 5507 9288
rect 4356 9284 4362 9286
rect 4245 9283 4311 9284
rect 5441 9283 5507 9286
rect 4685 9280 5005 9281
rect 4685 9216 4693 9280
rect 4757 9216 4773 9280
rect 4837 9216 4853 9280
rect 4917 9216 4933 9280
rect 4997 9216 5005 9280
rect 4685 9215 5005 9216
rect 8426 9280 8746 9281
rect 8426 9216 8434 9280
rect 8498 9216 8514 9280
rect 8578 9216 8594 9280
rect 8658 9216 8674 9280
rect 8738 9216 8746 9280
rect 8426 9215 8746 9216
rect 1393 9074 1459 9077
rect 6126 9074 6132 9076
rect 1393 9072 6132 9074
rect 1393 9016 1398 9072
rect 1454 9016 6132 9072
rect 1393 9014 6132 9016
rect 1393 9011 1459 9014
rect 6126 9012 6132 9014
rect 6196 9012 6202 9076
rect 3233 8938 3299 8941
rect 9438 8938 9444 8940
rect 3233 8936 9444 8938
rect 3233 8880 3238 8936
rect 3294 8880 9444 8936
rect 3233 8878 9444 8880
rect 3233 8875 3299 8878
rect 9438 8876 9444 8878
rect 9508 8876 9514 8940
rect 1485 8802 1551 8805
rect 2405 8802 2471 8805
rect 1485 8800 2471 8802
rect 1485 8744 1490 8800
rect 1546 8744 2410 8800
rect 2466 8744 2471 8800
rect 1485 8742 2471 8744
rect 1485 8739 1551 8742
rect 2405 8739 2471 8742
rect 2814 8736 3134 8737
rect 2814 8672 2822 8736
rect 2886 8672 2902 8736
rect 2966 8672 2982 8736
rect 3046 8672 3062 8736
rect 3126 8672 3134 8736
rect 2814 8671 3134 8672
rect 6556 8736 6876 8737
rect 6556 8672 6564 8736
rect 6628 8672 6644 8736
rect 6708 8672 6724 8736
rect 6788 8672 6804 8736
rect 6868 8672 6876 8736
rect 6556 8671 6876 8672
rect 10297 8736 10617 8737
rect 10297 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10545 8736
rect 10609 8672 10617 8736
rect 10297 8671 10617 8672
rect 2221 8668 2287 8669
rect 2221 8664 2268 8668
rect 2332 8666 2338 8668
rect 2221 8608 2226 8664
rect 2221 8604 2268 8608
rect 2332 8606 2378 8666
rect 2332 8604 2338 8606
rect 2221 8603 2287 8604
rect 1761 8530 1827 8533
rect 2773 8530 2839 8533
rect 3877 8530 3943 8533
rect 1761 8528 3943 8530
rect 1761 8472 1766 8528
rect 1822 8472 2778 8528
rect 2834 8472 3882 8528
rect 3938 8472 3943 8528
rect 1761 8470 3943 8472
rect 1761 8467 1827 8470
rect 2773 8467 2839 8470
rect 3877 8467 3943 8470
rect 2957 8394 3023 8397
rect 4102 8394 4108 8396
rect 2957 8392 4108 8394
rect 2957 8336 2962 8392
rect 3018 8336 4108 8392
rect 2957 8334 4108 8336
rect 2957 8331 3023 8334
rect 4102 8332 4108 8334
rect 4172 8332 4178 8396
rect 4470 8332 4476 8396
rect 4540 8394 4546 8396
rect 5073 8394 5139 8397
rect 5206 8394 5212 8396
rect 4540 8392 5212 8394
rect 4540 8336 5078 8392
rect 5134 8336 5212 8392
rect 4540 8334 5212 8336
rect 4540 8332 4546 8334
rect 5073 8331 5139 8334
rect 5206 8332 5212 8334
rect 5276 8394 5282 8396
rect 6085 8394 6151 8397
rect 5276 8392 6151 8394
rect 5276 8336 6090 8392
rect 6146 8336 6151 8392
rect 5276 8334 6151 8336
rect 5276 8332 5282 8334
rect 6085 8331 6151 8334
rect 7557 8394 7623 8397
rect 8886 8394 8892 8396
rect 7557 8392 8892 8394
rect 7557 8336 7562 8392
rect 7618 8336 8892 8392
rect 7557 8334 8892 8336
rect 7557 8331 7623 8334
rect 8886 8332 8892 8334
rect 8956 8332 8962 8396
rect 4685 8192 5005 8193
rect 4685 8128 4693 8192
rect 4757 8128 4773 8192
rect 4837 8128 4853 8192
rect 4917 8128 4933 8192
rect 4997 8128 5005 8192
rect 4685 8127 5005 8128
rect 8426 8192 8746 8193
rect 8426 8128 8434 8192
rect 8498 8128 8514 8192
rect 8578 8128 8594 8192
rect 8658 8128 8674 8192
rect 8738 8128 8746 8192
rect 8426 8127 8746 8128
rect 2129 7986 2195 7989
rect 8293 7986 8359 7989
rect 2129 7984 8359 7986
rect 2129 7928 2134 7984
rect 2190 7928 8298 7984
rect 8354 7928 8359 7984
rect 2129 7926 8359 7928
rect 2129 7923 2195 7926
rect 8293 7923 8359 7926
rect 8845 7986 8911 7989
rect 9070 7986 9076 7988
rect 8845 7984 9076 7986
rect 8845 7928 8850 7984
rect 8906 7928 9076 7984
rect 8845 7926 9076 7928
rect 8845 7923 8911 7926
rect 9070 7924 9076 7926
rect 9140 7924 9146 7988
rect 10961 7986 11027 7989
rect 9814 7984 11027 7986
rect 9814 7928 10966 7984
rect 11022 7928 11027 7984
rect 9814 7926 11027 7928
rect 5349 7852 5415 7853
rect 5349 7850 5396 7852
rect 5304 7848 5396 7850
rect 5304 7792 5354 7848
rect 5304 7790 5396 7792
rect 5349 7788 5396 7790
rect 5460 7788 5466 7852
rect 5349 7787 5415 7788
rect 9814 7717 9874 7926
rect 10961 7923 11027 7926
rect 9949 7852 10015 7853
rect 9949 7848 9996 7852
rect 10060 7850 10066 7852
rect 9949 7792 9954 7848
rect 9949 7788 9996 7792
rect 10060 7790 10106 7850
rect 10060 7788 10066 7790
rect 9949 7787 10015 7788
rect 9814 7712 9923 7717
rect 9814 7656 9862 7712
rect 9918 7656 9923 7712
rect 9814 7654 9923 7656
rect 9857 7651 9923 7654
rect 2814 7648 3134 7649
rect 2814 7584 2822 7648
rect 2886 7584 2902 7648
rect 2966 7584 2982 7648
rect 3046 7584 3062 7648
rect 3126 7584 3134 7648
rect 2814 7583 3134 7584
rect 6556 7648 6876 7649
rect 6556 7584 6564 7648
rect 6628 7584 6644 7648
rect 6708 7584 6724 7648
rect 6788 7584 6804 7648
rect 6868 7584 6876 7648
rect 6556 7583 6876 7584
rect 10297 7648 10617 7649
rect 10297 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10465 7648
rect 10529 7584 10545 7648
rect 10609 7584 10617 7648
rect 10297 7583 10617 7584
rect 3969 7578 4035 7581
rect 3420 7576 4035 7578
rect 3420 7520 3974 7576
rect 4030 7520 4035 7576
rect 3420 7518 4035 7520
rect 2313 7442 2379 7445
rect 2773 7442 2839 7445
rect 2313 7440 2839 7442
rect 2313 7384 2318 7440
rect 2374 7384 2778 7440
rect 2834 7384 2839 7440
rect 2313 7382 2839 7384
rect 2313 7379 2379 7382
rect 2773 7379 2839 7382
rect 3049 7442 3115 7445
rect 3420 7442 3480 7518
rect 3969 7515 4035 7518
rect 4429 7578 4495 7581
rect 5942 7578 5948 7580
rect 4429 7576 5948 7578
rect 4429 7520 4434 7576
rect 4490 7520 5948 7576
rect 4429 7518 5948 7520
rect 4429 7515 4495 7518
rect 5942 7516 5948 7518
rect 6012 7516 6018 7580
rect 3049 7440 3480 7442
rect 3049 7384 3054 7440
rect 3110 7384 3480 7440
rect 3049 7382 3480 7384
rect 3049 7379 3115 7382
rect 3550 7380 3556 7444
rect 3620 7442 3626 7444
rect 3693 7442 3759 7445
rect 3620 7440 3759 7442
rect 3620 7384 3698 7440
rect 3754 7384 3759 7440
rect 3620 7382 3759 7384
rect 3620 7380 3626 7382
rect 3693 7379 3759 7382
rect 4981 7442 5047 7445
rect 8150 7442 8156 7444
rect 4981 7440 8156 7442
rect 4981 7384 4986 7440
rect 5042 7384 8156 7440
rect 4981 7382 8156 7384
rect 4981 7379 5047 7382
rect 8150 7380 8156 7382
rect 8220 7380 8226 7444
rect 9673 7442 9739 7445
rect 10317 7442 10383 7445
rect 9673 7440 10383 7442
rect 9673 7384 9678 7440
rect 9734 7384 10322 7440
rect 10378 7384 10383 7440
rect 9673 7382 10383 7384
rect 9673 7379 9739 7382
rect 10317 7379 10383 7382
rect 749 7306 815 7309
rect 6453 7306 6519 7309
rect 749 7304 6519 7306
rect 749 7248 754 7304
rect 810 7248 6458 7304
rect 6514 7248 6519 7304
rect 749 7246 6519 7248
rect 749 7243 815 7246
rect 6453 7243 6519 7246
rect 4685 7104 5005 7105
rect 4685 7040 4693 7104
rect 4757 7040 4773 7104
rect 4837 7040 4853 7104
rect 4917 7040 4933 7104
rect 4997 7040 5005 7104
rect 4685 7039 5005 7040
rect 8426 7104 8746 7105
rect 8426 7040 8434 7104
rect 8498 7040 8514 7104
rect 8578 7040 8594 7104
rect 8658 7040 8674 7104
rect 8738 7040 8746 7104
rect 8426 7039 8746 7040
rect 1894 6972 1900 7036
rect 1964 7034 1970 7036
rect 2681 7034 2747 7037
rect 1964 7032 2747 7034
rect 1964 6976 2686 7032
rect 2742 6976 2747 7032
rect 1964 6974 2747 6976
rect 1964 6972 1970 6974
rect 2681 6971 2747 6974
rect 2957 7034 3023 7037
rect 4470 7034 4476 7036
rect 2957 7032 4476 7034
rect 2957 6976 2962 7032
rect 3018 6976 4476 7032
rect 2957 6974 4476 6976
rect 2957 6971 3023 6974
rect 4470 6972 4476 6974
rect 4540 6972 4546 7036
rect 9622 6972 9628 7036
rect 9692 7034 9698 7036
rect 10501 7034 10567 7037
rect 9692 7032 10567 7034
rect 9692 6976 10506 7032
rect 10562 6976 10567 7032
rect 9692 6974 10567 6976
rect 9692 6972 9698 6974
rect 10501 6971 10567 6974
rect 2630 6836 2636 6900
rect 2700 6898 2706 6900
rect 3325 6898 3391 6901
rect 2700 6896 3391 6898
rect 2700 6840 3330 6896
rect 3386 6840 3391 6896
rect 2700 6838 3391 6840
rect 2700 6836 2706 6838
rect 3325 6835 3391 6838
rect 1577 6762 1643 6765
rect 1853 6762 1919 6765
rect 1577 6760 1919 6762
rect 1577 6704 1582 6760
rect 1638 6704 1858 6760
rect 1914 6704 1919 6760
rect 1577 6702 1919 6704
rect 1577 6699 1643 6702
rect 1853 6699 1919 6702
rect 3325 6762 3391 6765
rect 5073 6762 5139 6765
rect 3325 6760 5139 6762
rect 3325 6704 3330 6760
rect 3386 6704 5078 6760
rect 5134 6704 5139 6760
rect 3325 6702 5139 6704
rect 3325 6699 3391 6702
rect 5073 6699 5139 6702
rect 5441 6762 5507 6765
rect 5717 6762 5783 6765
rect 5441 6760 5783 6762
rect 5441 6704 5446 6760
rect 5502 6704 5722 6760
rect 5778 6704 5783 6760
rect 5441 6702 5783 6704
rect 5441 6699 5507 6702
rect 5717 6699 5783 6702
rect 3969 6626 4035 6629
rect 4245 6626 4311 6629
rect 3969 6624 4311 6626
rect 3969 6568 3974 6624
rect 4030 6568 4250 6624
rect 4306 6568 4311 6624
rect 3969 6566 4311 6568
rect 3969 6563 4035 6566
rect 4245 6563 4311 6566
rect 5206 6564 5212 6628
rect 5276 6626 5282 6628
rect 5441 6626 5507 6629
rect 5276 6624 5507 6626
rect 5276 6568 5446 6624
rect 5502 6568 5507 6624
rect 5276 6566 5507 6568
rect 5276 6564 5282 6566
rect 5441 6563 5507 6566
rect 2814 6560 3134 6561
rect 2814 6496 2822 6560
rect 2886 6496 2902 6560
rect 2966 6496 2982 6560
rect 3046 6496 3062 6560
rect 3126 6496 3134 6560
rect 2814 6495 3134 6496
rect 6556 6560 6876 6561
rect 6556 6496 6564 6560
rect 6628 6496 6644 6560
rect 6708 6496 6724 6560
rect 6788 6496 6804 6560
rect 6868 6496 6876 6560
rect 6556 6495 6876 6496
rect 10297 6560 10617 6561
rect 10297 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10465 6560
rect 10529 6496 10545 6560
rect 10609 6496 10617 6560
rect 10297 6495 10617 6496
rect 3693 6490 3759 6493
rect 3969 6490 4035 6493
rect 3693 6488 4035 6490
rect 3693 6432 3698 6488
rect 3754 6432 3974 6488
rect 4030 6432 4035 6488
rect 3693 6430 4035 6432
rect 3693 6427 3759 6430
rect 3969 6427 4035 6430
rect 4613 6490 4679 6493
rect 5390 6490 5396 6492
rect 4613 6488 5396 6490
rect 4613 6432 4618 6488
rect 4674 6432 5396 6488
rect 4613 6430 5396 6432
rect 4613 6427 4679 6430
rect 5390 6428 5396 6430
rect 5460 6428 5466 6492
rect 5073 6354 5139 6357
rect 7189 6354 7255 6357
rect 5073 6352 7255 6354
rect 5073 6296 5078 6352
rect 5134 6296 7194 6352
rect 7250 6296 7255 6352
rect 5073 6294 7255 6296
rect 5073 6291 5139 6294
rect 7189 6291 7255 6294
rect 8477 6354 8543 6357
rect 9857 6354 9923 6357
rect 8477 6352 9923 6354
rect 8477 6296 8482 6352
rect 8538 6296 9862 6352
rect 9918 6296 9923 6352
rect 8477 6294 9923 6296
rect 8477 6291 8543 6294
rect 9857 6291 9923 6294
rect 2313 6218 2379 6221
rect 5206 6218 5212 6220
rect 2313 6216 5212 6218
rect 2313 6160 2318 6216
rect 2374 6160 5212 6216
rect 2313 6158 5212 6160
rect 2313 6155 2379 6158
rect 5206 6156 5212 6158
rect 5276 6156 5282 6220
rect 3918 6020 3924 6084
rect 3988 6082 3994 6084
rect 4061 6082 4127 6085
rect 7097 6082 7163 6085
rect 3988 6080 4127 6082
rect 3988 6024 4066 6080
rect 4122 6024 4127 6080
rect 3988 6022 4127 6024
rect 3988 6020 3994 6022
rect 4061 6019 4127 6022
rect 5214 6080 7163 6082
rect 5214 6024 7102 6080
rect 7158 6024 7163 6080
rect 5214 6022 7163 6024
rect 4685 6016 5005 6017
rect 4685 5952 4693 6016
rect 4757 5952 4773 6016
rect 4837 5952 4853 6016
rect 4917 5952 4933 6016
rect 4997 5952 5005 6016
rect 4685 5951 5005 5952
rect 5214 5949 5274 6022
rect 7097 6019 7163 6022
rect 8426 6016 8746 6017
rect 8426 5952 8434 6016
rect 8498 5952 8514 6016
rect 8578 5952 8594 6016
rect 8658 5952 8674 6016
rect 8738 5952 8746 6016
rect 8426 5951 8746 5952
rect 3233 5946 3299 5949
rect 3233 5944 4584 5946
rect 3233 5888 3238 5944
rect 3294 5888 4584 5944
rect 3233 5886 4584 5888
rect 3233 5883 3299 5886
rect 4524 5810 4584 5886
rect 5165 5944 5274 5949
rect 5165 5888 5170 5944
rect 5226 5888 5274 5944
rect 5165 5886 5274 5888
rect 5165 5883 5231 5886
rect 7782 5810 7788 5812
rect 4524 5750 7788 5810
rect 7782 5748 7788 5750
rect 7852 5748 7858 5812
rect 2957 5674 3023 5677
rect 7414 5674 7420 5676
rect 2957 5672 7420 5674
rect 2957 5616 2962 5672
rect 3018 5616 7420 5672
rect 2957 5614 7420 5616
rect 2957 5611 3023 5614
rect 7414 5612 7420 5614
rect 7484 5612 7490 5676
rect 9806 5612 9812 5676
rect 9876 5674 9882 5676
rect 10225 5674 10291 5677
rect 9876 5672 10291 5674
rect 9876 5616 10230 5672
rect 10286 5616 10291 5672
rect 9876 5614 10291 5616
rect 9876 5612 9882 5614
rect 10225 5611 10291 5614
rect 8569 5538 8635 5541
rect 10041 5538 10107 5541
rect 8569 5536 10107 5538
rect 8569 5480 8574 5536
rect 8630 5480 10046 5536
rect 10102 5480 10107 5536
rect 8569 5478 10107 5480
rect 8569 5475 8635 5478
rect 10041 5475 10107 5478
rect 2814 5472 3134 5473
rect 2814 5408 2822 5472
rect 2886 5408 2902 5472
rect 2966 5408 2982 5472
rect 3046 5408 3062 5472
rect 3126 5408 3134 5472
rect 2814 5407 3134 5408
rect 6556 5472 6876 5473
rect 6556 5408 6564 5472
rect 6628 5408 6644 5472
rect 6708 5408 6724 5472
rect 6788 5408 6804 5472
rect 6868 5408 6876 5472
rect 6556 5407 6876 5408
rect 10297 5472 10617 5473
rect 10297 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10545 5472
rect 10609 5408 10617 5472
rect 10297 5407 10617 5408
rect 5993 5404 6059 5405
rect 5942 5340 5948 5404
rect 6012 5402 6059 5404
rect 7557 5402 7623 5405
rect 9581 5402 9647 5405
rect 6012 5400 6104 5402
rect 6054 5344 6104 5400
rect 6012 5342 6104 5344
rect 7557 5400 9647 5402
rect 7557 5344 7562 5400
rect 7618 5344 9586 5400
rect 9642 5344 9647 5400
rect 7557 5342 9647 5344
rect 6012 5340 6059 5342
rect 5993 5339 6059 5340
rect 7557 5339 7623 5342
rect 9581 5339 9647 5342
rect 5490 5206 7850 5266
rect 5490 5133 5550 5206
rect 5441 5128 5550 5133
rect 5441 5072 5446 5128
rect 5502 5072 5550 5128
rect 5441 5070 5550 5072
rect 5625 5130 5691 5133
rect 5942 5130 5948 5132
rect 5625 5128 5948 5130
rect 5625 5072 5630 5128
rect 5686 5072 5948 5128
rect 5625 5070 5948 5072
rect 5441 5067 5507 5070
rect 5625 5067 5691 5070
rect 5942 5068 5948 5070
rect 6012 5068 6018 5132
rect 7790 5130 7850 5206
rect 7966 5204 7972 5268
rect 8036 5266 8042 5268
rect 8937 5266 9003 5269
rect 8036 5264 9003 5266
rect 8036 5208 8942 5264
rect 8998 5208 9003 5264
rect 8036 5206 9003 5208
rect 8036 5204 8042 5206
rect 8937 5203 9003 5206
rect 9121 5266 9187 5269
rect 9673 5266 9739 5269
rect 9121 5264 9739 5266
rect 9121 5208 9126 5264
rect 9182 5208 9678 5264
rect 9734 5208 9739 5264
rect 9121 5206 9739 5208
rect 9121 5203 9187 5206
rect 9673 5203 9739 5206
rect 10593 5130 10659 5133
rect 7790 5128 10659 5130
rect 7790 5072 10598 5128
rect 10654 5072 10659 5128
rect 7790 5070 10659 5072
rect 10593 5067 10659 5070
rect 5390 4932 5396 4996
rect 5460 4994 5466 4996
rect 7966 4994 7972 4996
rect 5460 4934 7972 4994
rect 5460 4932 5466 4934
rect 7966 4932 7972 4934
rect 8036 4932 8042 4996
rect 4685 4928 5005 4929
rect 4685 4864 4693 4928
rect 4757 4864 4773 4928
rect 4837 4864 4853 4928
rect 4917 4864 4933 4928
rect 4997 4864 5005 4928
rect 4685 4863 5005 4864
rect 8426 4928 8746 4929
rect 8426 4864 8434 4928
rect 8498 4864 8514 4928
rect 8578 4864 8594 4928
rect 8658 4864 8674 4928
rect 8738 4864 8746 4928
rect 8426 4863 8746 4864
rect 5901 4858 5967 4861
rect 7833 4858 7899 4861
rect 9489 4860 9555 4861
rect 5901 4856 7899 4858
rect 5901 4800 5906 4856
rect 5962 4800 7838 4856
rect 7894 4800 7899 4856
rect 5901 4798 7899 4800
rect 5901 4795 5967 4798
rect 7833 4795 7899 4798
rect 9438 4796 9444 4860
rect 9508 4858 9555 4860
rect 9508 4856 9600 4858
rect 9550 4800 9600 4856
rect 9508 4798 9600 4800
rect 9508 4796 9555 4798
rect 9489 4795 9555 4796
rect 5390 4660 5396 4724
rect 5460 4722 5466 4724
rect 6177 4722 6243 4725
rect 5460 4720 6243 4722
rect 5460 4664 6182 4720
rect 6238 4664 6243 4720
rect 5460 4662 6243 4664
rect 5460 4660 5466 4662
rect 6177 4659 6243 4662
rect 6361 4722 6427 4725
rect 10910 4722 10916 4724
rect 6361 4720 10916 4722
rect 6361 4664 6366 4720
rect 6422 4664 10916 4720
rect 6361 4662 10916 4664
rect 6361 4659 6427 4662
rect 10910 4660 10916 4662
rect 10980 4660 10986 4724
rect 3601 4584 3667 4589
rect 3601 4528 3606 4584
rect 3662 4528 3667 4584
rect 3601 4523 3667 4528
rect 3734 4524 3740 4588
rect 3804 4586 3810 4588
rect 4429 4586 4495 4589
rect 3804 4584 4495 4586
rect 3804 4528 4434 4584
rect 4490 4528 4495 4584
rect 3804 4526 4495 4528
rect 3804 4524 3810 4526
rect 4429 4523 4495 4526
rect 6269 4586 6335 4589
rect 6913 4586 6979 4589
rect 6269 4584 6979 4586
rect 6269 4528 6274 4584
rect 6330 4528 6918 4584
rect 6974 4528 6979 4584
rect 6269 4526 6979 4528
rect 6269 4523 6335 4526
rect 6913 4523 6979 4526
rect 7649 4586 7715 4589
rect 9673 4586 9739 4589
rect 10961 4586 11027 4589
rect 7649 4584 11027 4586
rect 7649 4528 7654 4584
rect 7710 4528 9678 4584
rect 9734 4528 10966 4584
rect 11022 4528 11027 4584
rect 7649 4526 11027 4528
rect 7649 4523 7715 4526
rect 9673 4523 9739 4526
rect 10961 4523 11027 4526
rect 3604 4450 3664 4523
rect 6085 4450 6151 4453
rect 3604 4448 6151 4450
rect 3604 4392 6090 4448
rect 6146 4392 6151 4448
rect 3604 4390 6151 4392
rect 6085 4387 6151 4390
rect 2814 4384 3134 4385
rect 2814 4320 2822 4384
rect 2886 4320 2902 4384
rect 2966 4320 2982 4384
rect 3046 4320 3062 4384
rect 3126 4320 3134 4384
rect 2814 4319 3134 4320
rect 6556 4384 6876 4385
rect 6556 4320 6564 4384
rect 6628 4320 6644 4384
rect 6708 4320 6724 4384
rect 6788 4320 6804 4384
rect 6868 4320 6876 4384
rect 6556 4319 6876 4320
rect 10297 4384 10617 4385
rect 10297 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10545 4384
rect 10609 4320 10617 4384
rect 10297 4319 10617 4320
rect 3918 4252 3924 4316
rect 3988 4314 3994 4316
rect 4061 4314 4127 4317
rect 3988 4312 4127 4314
rect 3988 4256 4066 4312
rect 4122 4256 4127 4312
rect 3988 4254 4127 4256
rect 3988 4252 3994 4254
rect 4061 4251 4127 4254
rect 3918 4116 3924 4180
rect 3988 4178 3994 4180
rect 5574 4178 5580 4180
rect 3988 4118 5580 4178
rect 3988 4116 3994 4118
rect 5574 4116 5580 4118
rect 5644 4116 5650 4180
rect 5993 4178 6059 4181
rect 9254 4178 9260 4180
rect 5993 4176 9260 4178
rect 5993 4120 5998 4176
rect 6054 4120 9260 4176
rect 5993 4118 9260 4120
rect 5993 4115 6059 4118
rect 9254 4116 9260 4118
rect 9324 4116 9330 4180
rect 749 4042 815 4045
rect 974 4042 980 4044
rect 749 4040 980 4042
rect 749 3984 754 4040
rect 810 3984 980 4040
rect 749 3982 980 3984
rect 749 3979 815 3982
rect 974 3980 980 3982
rect 1044 3980 1050 4044
rect 1669 4042 1735 4045
rect 7373 4042 7439 4045
rect 1669 4040 7439 4042
rect 1669 3984 1674 4040
rect 1730 3984 7378 4040
rect 7434 3984 7439 4040
rect 1669 3982 7439 3984
rect 1669 3979 1735 3982
rect 7373 3979 7439 3982
rect 8109 4042 8175 4045
rect 9397 4042 9463 4045
rect 8109 4040 9463 4042
rect 8109 3984 8114 4040
rect 8170 3984 9402 4040
rect 9458 3984 9463 4040
rect 8109 3982 9463 3984
rect 8109 3979 8175 3982
rect 9397 3979 9463 3982
rect 3325 3906 3391 3909
rect 3877 3906 3943 3909
rect 3325 3904 3943 3906
rect 3325 3848 3330 3904
rect 3386 3848 3882 3904
rect 3938 3848 3943 3904
rect 3325 3846 3943 3848
rect 3325 3843 3391 3846
rect 3877 3843 3943 3846
rect 5165 3906 5231 3909
rect 5993 3906 6059 3909
rect 5165 3904 6059 3906
rect 5165 3848 5170 3904
rect 5226 3848 5998 3904
rect 6054 3848 6059 3904
rect 5165 3846 6059 3848
rect 5165 3843 5231 3846
rect 5993 3843 6059 3846
rect 6913 3906 6979 3909
rect 8293 3906 8359 3909
rect 6913 3904 8359 3906
rect 6913 3848 6918 3904
rect 6974 3848 8298 3904
rect 8354 3848 8359 3904
rect 6913 3846 8359 3848
rect 6913 3843 6979 3846
rect 8293 3843 8359 3846
rect 4685 3840 5005 3841
rect 4685 3776 4693 3840
rect 4757 3776 4773 3840
rect 4837 3776 4853 3840
rect 4917 3776 4933 3840
rect 4997 3776 5005 3840
rect 4685 3775 5005 3776
rect 8426 3840 8746 3841
rect 8426 3776 8434 3840
rect 8498 3776 8514 3840
rect 8578 3776 8594 3840
rect 8658 3776 8674 3840
rect 8738 3776 8746 3840
rect 8426 3775 8746 3776
rect 4337 3770 4403 3773
rect 6269 3770 6335 3773
rect 4337 3768 4584 3770
rect 4337 3712 4342 3768
rect 4398 3712 4584 3768
rect 4337 3710 4584 3712
rect 4337 3707 4403 3710
rect 1853 3634 1919 3637
rect 2078 3634 2084 3636
rect 1853 3632 2084 3634
rect 1853 3576 1858 3632
rect 1914 3576 2084 3632
rect 1853 3574 2084 3576
rect 1853 3571 1919 3574
rect 2078 3572 2084 3574
rect 2148 3572 2154 3636
rect 4524 3634 4584 3710
rect 6269 3768 7666 3770
rect 6269 3712 6274 3768
rect 6330 3712 7666 3768
rect 6269 3710 7666 3712
rect 6269 3707 6335 3710
rect 4797 3634 4863 3637
rect 4524 3632 4863 3634
rect 4524 3576 4802 3632
rect 4858 3576 4863 3632
rect 4524 3574 4863 3576
rect 4797 3571 4863 3574
rect 5625 3634 5691 3637
rect 6913 3634 6979 3637
rect 5625 3632 6979 3634
rect 5625 3576 5630 3632
rect 5686 3576 6918 3632
rect 6974 3576 6979 3632
rect 5625 3574 6979 3576
rect 7606 3634 7666 3710
rect 8753 3634 8819 3637
rect 7606 3632 8819 3634
rect 7606 3576 8758 3632
rect 8814 3576 8819 3632
rect 7606 3574 8819 3576
rect 5625 3571 5691 3574
rect 6913 3571 6979 3574
rect 8753 3571 8819 3574
rect 9673 3634 9739 3637
rect 13169 3634 13235 3637
rect 9673 3632 13235 3634
rect 9673 3576 9678 3632
rect 9734 3576 13174 3632
rect 13230 3576 13235 3632
rect 9673 3574 13235 3576
rect 9673 3571 9739 3574
rect 13169 3571 13235 3574
rect 4286 3436 4292 3500
rect 4356 3498 4362 3500
rect 4521 3498 4587 3501
rect 4356 3496 4587 3498
rect 4356 3440 4526 3496
rect 4582 3440 4587 3496
rect 4356 3438 4587 3440
rect 4356 3436 4362 3438
rect 4521 3435 4587 3438
rect 6177 3498 6243 3501
rect 8661 3498 8727 3501
rect 6177 3496 8727 3498
rect 6177 3440 6182 3496
rect 6238 3440 8666 3496
rect 8722 3440 8727 3496
rect 6177 3438 8727 3440
rect 6177 3435 6243 3438
rect 8661 3435 8727 3438
rect 10910 3436 10916 3500
rect 10980 3498 10986 3500
rect 11053 3498 11119 3501
rect 10980 3496 11119 3498
rect 10980 3440 11058 3496
rect 11114 3440 11119 3496
rect 10980 3438 11119 3440
rect 10980 3436 10986 3438
rect 11053 3435 11119 3438
rect 2814 3296 3134 3297
rect 2814 3232 2822 3296
rect 2886 3232 2902 3296
rect 2966 3232 2982 3296
rect 3046 3232 3062 3296
rect 3126 3232 3134 3296
rect 2814 3231 3134 3232
rect 6556 3296 6876 3297
rect 6556 3232 6564 3296
rect 6628 3232 6644 3296
rect 6708 3232 6724 3296
rect 6788 3232 6804 3296
rect 6868 3232 6876 3296
rect 6556 3231 6876 3232
rect 10297 3296 10617 3297
rect 10297 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10545 3296
rect 10609 3232 10617 3296
rect 10297 3231 10617 3232
rect 1761 3228 1827 3229
rect 1710 3226 1716 3228
rect 1670 3166 1716 3226
rect 1780 3224 1827 3228
rect 1822 3168 1827 3224
rect 1710 3164 1716 3166
rect 1780 3164 1827 3168
rect 1761 3163 1827 3164
rect 5257 3226 5323 3229
rect 5533 3226 5599 3229
rect 8753 3226 8819 3229
rect 8886 3226 8892 3228
rect 5257 3224 5458 3226
rect 5257 3168 5262 3224
rect 5318 3168 5458 3224
rect 5257 3166 5458 3168
rect 5257 3163 5323 3166
rect 3233 3090 3299 3093
rect 3366 3090 3372 3092
rect 3233 3088 3372 3090
rect 3233 3032 3238 3088
rect 3294 3032 3372 3088
rect 3233 3030 3372 3032
rect 3233 3027 3299 3030
rect 3366 3028 3372 3030
rect 3436 3028 3442 3092
rect 657 2954 723 2957
rect 933 2954 999 2957
rect 657 2952 999 2954
rect 657 2896 662 2952
rect 718 2896 938 2952
rect 994 2896 999 2952
rect 657 2894 999 2896
rect 657 2891 723 2894
rect 933 2891 999 2894
rect 1117 2954 1183 2957
rect 1853 2954 1919 2957
rect 2446 2954 2452 2956
rect 1117 2952 1410 2954
rect 1117 2896 1122 2952
rect 1178 2896 1410 2952
rect 1117 2894 1410 2896
rect 1117 2891 1183 2894
rect 1350 2818 1410 2894
rect 1853 2952 2452 2954
rect 1853 2896 1858 2952
rect 1914 2896 2452 2952
rect 1853 2894 2452 2896
rect 1853 2891 1919 2894
rect 2446 2892 2452 2894
rect 2516 2892 2522 2956
rect 3141 2954 3207 2957
rect 4153 2956 4219 2957
rect 3550 2954 3556 2956
rect 3141 2952 3556 2954
rect 3141 2896 3146 2952
rect 3202 2896 3556 2952
rect 3141 2894 3556 2896
rect 3141 2891 3207 2894
rect 3550 2892 3556 2894
rect 3620 2892 3626 2956
rect 3918 2954 3924 2956
rect 3742 2894 3924 2954
rect 1853 2818 1919 2821
rect 2313 2820 2379 2821
rect 1350 2816 1919 2818
rect 1350 2760 1858 2816
rect 1914 2760 1919 2816
rect 1350 2758 1919 2760
rect 1853 2755 1919 2758
rect 2262 2756 2268 2820
rect 2332 2818 2379 2820
rect 2332 2816 2424 2818
rect 2374 2760 2424 2816
rect 2332 2758 2424 2760
rect 2332 2756 2379 2758
rect 2313 2755 2379 2756
rect 3742 2685 3802 2894
rect 3918 2892 3924 2894
rect 3988 2892 3994 2956
rect 4102 2954 4108 2956
rect 4062 2894 4108 2954
rect 4172 2952 4219 2956
rect 4797 2954 4863 2957
rect 5398 2956 5458 3166
rect 5533 3224 6378 3226
rect 5533 3168 5538 3224
rect 5594 3168 6378 3224
rect 5533 3166 6378 3168
rect 5533 3163 5599 3166
rect 5533 3092 5599 3093
rect 5533 3088 5580 3092
rect 5644 3090 5650 3092
rect 6318 3090 6378 3166
rect 8753 3224 8892 3226
rect 8753 3168 8758 3224
rect 8814 3168 8892 3224
rect 8753 3166 8892 3168
rect 8753 3163 8819 3166
rect 8886 3164 8892 3166
rect 8956 3164 8962 3228
rect 6453 3090 6519 3093
rect 5533 3032 5538 3088
rect 5533 3028 5580 3032
rect 5644 3030 5690 3090
rect 6318 3088 6519 3090
rect 6318 3032 6458 3088
rect 6514 3032 6519 3088
rect 6318 3030 6519 3032
rect 5644 3028 5650 3030
rect 5533 3027 5599 3028
rect 6453 3027 6519 3030
rect 6637 3090 6703 3093
rect 8477 3090 8543 3093
rect 10041 3092 10107 3093
rect 6637 3088 8543 3090
rect 6637 3032 6642 3088
rect 6698 3032 8482 3088
rect 8538 3032 8543 3088
rect 6637 3030 8543 3032
rect 6637 3027 6703 3030
rect 8477 3027 8543 3030
rect 9990 3028 9996 3092
rect 10060 3090 10107 3092
rect 10060 3088 10152 3090
rect 10102 3032 10152 3088
rect 10060 3030 10152 3032
rect 10060 3028 10107 3030
rect 10041 3027 10107 3028
rect 4214 2896 4219 2952
rect 4102 2892 4108 2894
rect 4172 2892 4219 2896
rect 4153 2891 4219 2892
rect 4294 2952 4863 2954
rect 4294 2896 4802 2952
rect 4858 2896 4863 2952
rect 4294 2894 4863 2896
rect 3877 2818 3943 2821
rect 4294 2818 4354 2894
rect 4797 2891 4863 2894
rect 5390 2892 5396 2956
rect 5460 2892 5466 2956
rect 6310 2892 6316 2956
rect 6380 2954 6386 2956
rect 6821 2954 6887 2957
rect 7598 2954 7604 2956
rect 6380 2952 6887 2954
rect 6380 2896 6826 2952
rect 6882 2896 6887 2952
rect 6380 2894 6887 2896
rect 6380 2892 6386 2894
rect 6821 2891 6887 2894
rect 7054 2894 7604 2954
rect 7054 2818 7114 2894
rect 7598 2892 7604 2894
rect 7668 2892 7674 2956
rect 8109 2954 8175 2957
rect 9806 2954 9812 2956
rect 8109 2952 9812 2954
rect 8109 2896 8114 2952
rect 8170 2896 9812 2952
rect 8109 2894 9812 2896
rect 8109 2891 8175 2894
rect 9806 2892 9812 2894
rect 9876 2892 9882 2956
rect 3877 2816 4354 2818
rect 3877 2760 3882 2816
rect 3938 2760 4354 2816
rect 3877 2758 4354 2760
rect 5214 2758 7114 2818
rect 7557 2818 7623 2821
rect 7782 2818 7788 2820
rect 7557 2816 7788 2818
rect 7557 2760 7562 2816
rect 7618 2760 7788 2816
rect 7557 2758 7788 2760
rect 3877 2755 3943 2758
rect 4685 2752 5005 2753
rect 4685 2688 4693 2752
rect 4757 2688 4773 2752
rect 4837 2688 4853 2752
rect 4917 2688 4933 2752
rect 4997 2688 5005 2752
rect 4685 2687 5005 2688
rect 3742 2680 3851 2685
rect 3742 2624 3790 2680
rect 3846 2624 3851 2680
rect 3742 2622 3851 2624
rect 3785 2619 3851 2622
rect 3969 2682 4035 2685
rect 4102 2682 4108 2684
rect 3969 2680 4108 2682
rect 3969 2624 3974 2680
rect 4030 2624 4108 2680
rect 3969 2622 4108 2624
rect 3969 2619 4035 2622
rect 4102 2620 4108 2622
rect 4172 2620 4178 2684
rect 2865 2546 2931 2549
rect 3734 2546 3740 2548
rect 2865 2544 3740 2546
rect 2865 2488 2870 2544
rect 2926 2488 3740 2544
rect 2865 2486 3740 2488
rect 2865 2483 2931 2486
rect 3734 2484 3740 2486
rect 3804 2484 3810 2548
rect 4705 2546 4771 2549
rect 5214 2546 5274 2758
rect 7557 2755 7623 2758
rect 7782 2756 7788 2758
rect 7852 2756 7858 2820
rect 8426 2752 8746 2753
rect 8426 2688 8434 2752
rect 8498 2688 8514 2752
rect 8578 2688 8594 2752
rect 8658 2688 8674 2752
rect 8738 2688 8746 2752
rect 8426 2687 8746 2688
rect 5717 2682 5783 2685
rect 6126 2682 6132 2684
rect 5717 2680 6132 2682
rect 5717 2624 5722 2680
rect 5778 2624 6132 2680
rect 5717 2622 6132 2624
rect 5717 2619 5783 2622
rect 6126 2620 6132 2622
rect 6196 2620 6202 2684
rect 4705 2544 5274 2546
rect 4705 2488 4710 2544
rect 4766 2488 5274 2544
rect 4705 2486 5274 2488
rect 4705 2483 4771 2486
rect 5942 2484 5948 2548
rect 6012 2546 6018 2548
rect 7833 2546 7899 2549
rect 6012 2544 7899 2546
rect 6012 2488 7838 2544
rect 7894 2488 7899 2544
rect 6012 2486 7899 2488
rect 6012 2484 6018 2486
rect 7833 2483 7899 2486
rect 8150 2484 8156 2548
rect 8220 2546 8226 2548
rect 8477 2546 8543 2549
rect 8220 2544 8543 2546
rect 8220 2488 8482 2544
rect 8538 2488 8543 2544
rect 8220 2486 8543 2488
rect 8220 2484 8226 2486
rect 8477 2483 8543 2486
rect 8661 2546 8727 2549
rect 9857 2546 9923 2549
rect 8661 2544 9923 2546
rect 8661 2488 8666 2544
rect 8722 2488 9862 2544
rect 9918 2488 9923 2544
rect 8661 2486 9923 2488
rect 8661 2483 8727 2486
rect 9857 2483 9923 2486
rect 10317 2546 10383 2549
rect 12433 2546 12499 2549
rect 10317 2544 12499 2546
rect 10317 2488 10322 2544
rect 10378 2488 12438 2544
rect 12494 2488 12499 2544
rect 10317 2486 12499 2488
rect 10317 2483 10383 2486
rect 12433 2483 12499 2486
rect 5206 2348 5212 2412
rect 5276 2410 5282 2412
rect 5625 2410 5691 2413
rect 5276 2408 5691 2410
rect 5276 2352 5630 2408
rect 5686 2352 5691 2408
rect 5276 2350 5691 2352
rect 5276 2348 5282 2350
rect 5625 2347 5691 2350
rect 8385 2410 8451 2413
rect 9070 2410 9076 2412
rect 8385 2408 9076 2410
rect 8385 2352 8390 2408
rect 8446 2352 9076 2408
rect 8385 2350 9076 2352
rect 8385 2347 8451 2350
rect 9070 2348 9076 2350
rect 9140 2348 9146 2412
rect 10225 2410 10291 2413
rect 10777 2410 10843 2413
rect 10225 2408 10843 2410
rect 10225 2352 10230 2408
rect 10286 2352 10782 2408
rect 10838 2352 10843 2408
rect 10225 2350 10843 2352
rect 10225 2347 10291 2350
rect 10777 2347 10843 2350
rect 7414 2212 7420 2276
rect 7484 2274 7490 2276
rect 8661 2274 8727 2277
rect 7484 2272 8727 2274
rect 7484 2216 8666 2272
rect 8722 2216 8727 2272
rect 7484 2214 8727 2216
rect 7484 2212 7490 2214
rect 8661 2211 8727 2214
rect 2814 2208 3134 2209
rect 2814 2144 2822 2208
rect 2886 2144 2902 2208
rect 2966 2144 2982 2208
rect 3046 2144 3062 2208
rect 3126 2144 3134 2208
rect 2814 2143 3134 2144
rect 6556 2208 6876 2209
rect 6556 2144 6564 2208
rect 6628 2144 6644 2208
rect 6708 2144 6724 2208
rect 6788 2144 6804 2208
rect 6868 2144 6876 2208
rect 6556 2143 6876 2144
rect 10297 2208 10617 2209
rect 10297 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10545 2208
rect 10609 2144 10617 2208
rect 10297 2143 10617 2144
rect 5390 1940 5396 2004
rect 5460 2002 5466 2004
rect 6729 2002 6795 2005
rect 5460 2000 6795 2002
rect 5460 1944 6734 2000
rect 6790 1944 6795 2000
rect 5460 1942 6795 1944
rect 5460 1940 5466 1942
rect 6729 1939 6795 1942
rect 2589 1868 2655 1869
rect 2589 1866 2636 1868
rect 2544 1864 2636 1866
rect 2544 1808 2594 1864
rect 2544 1806 2636 1808
rect 2589 1804 2636 1806
rect 2700 1804 2706 1868
rect 6361 1866 6427 1869
rect 7046 1866 7052 1868
rect 6361 1864 7052 1866
rect 6361 1808 6366 1864
rect 6422 1808 7052 1864
rect 6361 1806 7052 1808
rect 2589 1803 2655 1804
rect 6361 1803 6427 1806
rect 7046 1804 7052 1806
rect 7116 1804 7122 1868
rect 1710 1668 1716 1732
rect 1780 1730 1786 1732
rect 5993 1730 6059 1733
rect 1780 1728 6059 1730
rect 1780 1672 5998 1728
rect 6054 1672 6059 1728
rect 1780 1670 6059 1672
rect 1780 1668 1786 1670
rect 5993 1667 6059 1670
rect 7966 1668 7972 1732
rect 8036 1730 8042 1732
rect 8753 1730 8819 1733
rect 8036 1728 8819 1730
rect 8036 1672 8758 1728
rect 8814 1672 8819 1728
rect 8036 1670 8819 1672
rect 8036 1668 8042 1670
rect 8753 1667 8819 1670
rect 1894 1532 1900 1596
rect 1964 1594 1970 1596
rect 5257 1594 5323 1597
rect 1964 1592 5323 1594
rect 1964 1536 5262 1592
rect 5318 1536 5323 1592
rect 1964 1534 5323 1536
rect 1964 1532 1970 1534
rect 5257 1531 5323 1534
rect 5758 1458 5764 1460
rect 4110 1398 5764 1458
rect 4110 1189 4170 1398
rect 5758 1396 5764 1398
rect 5828 1396 5834 1460
rect 4470 1260 4476 1324
rect 4540 1322 4546 1324
rect 5533 1322 5599 1325
rect 4540 1320 5599 1322
rect 4540 1264 5538 1320
rect 5594 1264 5599 1320
rect 4540 1262 5599 1264
rect 4540 1260 4546 1262
rect 5533 1259 5599 1262
rect 8845 1322 8911 1325
rect 9254 1322 9260 1324
rect 8845 1320 9260 1322
rect 8845 1264 8850 1320
rect 8906 1264 9260 1320
rect 8845 1262 9260 1264
rect 8845 1259 8911 1262
rect 9254 1260 9260 1262
rect 9324 1260 9330 1324
rect 4061 1184 4170 1189
rect 4061 1128 4066 1184
rect 4122 1128 4170 1184
rect 4061 1126 4170 1128
rect 4521 1186 4587 1189
rect 7230 1186 7236 1188
rect 4521 1184 7236 1186
rect 4521 1128 4526 1184
rect 4582 1128 7236 1184
rect 4521 1126 7236 1128
rect 4061 1123 4127 1126
rect 4521 1123 4587 1126
rect 7230 1124 7236 1126
rect 7300 1124 7306 1188
rect 4286 988 4292 1052
rect 4356 1050 4362 1052
rect 5901 1050 5967 1053
rect 4356 1048 5967 1050
rect 4356 992 5906 1048
rect 5962 992 5967 1048
rect 4356 990 5967 992
rect 4356 988 4362 990
rect 5901 987 5967 990
<< via3 >>
rect 2822 13084 2886 13088
rect 2822 13028 2826 13084
rect 2826 13028 2882 13084
rect 2882 13028 2886 13084
rect 2822 13024 2886 13028
rect 2902 13084 2966 13088
rect 2902 13028 2906 13084
rect 2906 13028 2962 13084
rect 2962 13028 2966 13084
rect 2902 13024 2966 13028
rect 2982 13084 3046 13088
rect 2982 13028 2986 13084
rect 2986 13028 3042 13084
rect 3042 13028 3046 13084
rect 2982 13024 3046 13028
rect 3062 13084 3126 13088
rect 3062 13028 3066 13084
rect 3066 13028 3122 13084
rect 3122 13028 3126 13084
rect 3062 13024 3126 13028
rect 6564 13084 6628 13088
rect 6564 13028 6568 13084
rect 6568 13028 6624 13084
rect 6624 13028 6628 13084
rect 6564 13024 6628 13028
rect 6644 13084 6708 13088
rect 6644 13028 6648 13084
rect 6648 13028 6704 13084
rect 6704 13028 6708 13084
rect 6644 13024 6708 13028
rect 6724 13084 6788 13088
rect 6724 13028 6728 13084
rect 6728 13028 6784 13084
rect 6784 13028 6788 13084
rect 6724 13024 6788 13028
rect 6804 13084 6868 13088
rect 6804 13028 6808 13084
rect 6808 13028 6864 13084
rect 6864 13028 6868 13084
rect 6804 13024 6868 13028
rect 10305 13084 10369 13088
rect 10305 13028 10309 13084
rect 10309 13028 10365 13084
rect 10365 13028 10369 13084
rect 10305 13024 10369 13028
rect 10385 13084 10449 13088
rect 10385 13028 10389 13084
rect 10389 13028 10445 13084
rect 10445 13028 10449 13084
rect 10385 13024 10449 13028
rect 10465 13084 10529 13088
rect 10465 13028 10469 13084
rect 10469 13028 10525 13084
rect 10525 13028 10529 13084
rect 10465 13024 10529 13028
rect 10545 13084 10609 13088
rect 10545 13028 10549 13084
rect 10549 13028 10605 13084
rect 10605 13028 10609 13084
rect 10545 13024 10609 13028
rect 2084 12548 2148 12612
rect 2452 12608 2516 12612
rect 2452 12552 2466 12608
rect 2466 12552 2516 12608
rect 2452 12548 2516 12552
rect 4693 12540 4757 12544
rect 4693 12484 4697 12540
rect 4697 12484 4753 12540
rect 4753 12484 4757 12540
rect 4693 12480 4757 12484
rect 4773 12540 4837 12544
rect 4773 12484 4777 12540
rect 4777 12484 4833 12540
rect 4833 12484 4837 12540
rect 4773 12480 4837 12484
rect 4853 12540 4917 12544
rect 4853 12484 4857 12540
rect 4857 12484 4913 12540
rect 4913 12484 4917 12540
rect 4853 12480 4917 12484
rect 4933 12540 4997 12544
rect 4933 12484 4937 12540
rect 4937 12484 4993 12540
rect 4993 12484 4997 12540
rect 4933 12480 4997 12484
rect 8434 12540 8498 12544
rect 8434 12484 8438 12540
rect 8438 12484 8494 12540
rect 8494 12484 8498 12540
rect 8434 12480 8498 12484
rect 8514 12540 8578 12544
rect 8514 12484 8518 12540
rect 8518 12484 8574 12540
rect 8574 12484 8578 12540
rect 8514 12480 8578 12484
rect 8594 12540 8658 12544
rect 8594 12484 8598 12540
rect 8598 12484 8654 12540
rect 8654 12484 8658 12540
rect 8594 12480 8658 12484
rect 8674 12540 8738 12544
rect 8674 12484 8678 12540
rect 8678 12484 8734 12540
rect 8734 12484 8738 12540
rect 8674 12480 8738 12484
rect 2822 11996 2886 12000
rect 2822 11940 2826 11996
rect 2826 11940 2882 11996
rect 2882 11940 2886 11996
rect 2822 11936 2886 11940
rect 2902 11996 2966 12000
rect 2902 11940 2906 11996
rect 2906 11940 2962 11996
rect 2962 11940 2966 11996
rect 2902 11936 2966 11940
rect 2982 11996 3046 12000
rect 2982 11940 2986 11996
rect 2986 11940 3042 11996
rect 3042 11940 3046 11996
rect 2982 11936 3046 11940
rect 3062 11996 3126 12000
rect 3062 11940 3066 11996
rect 3066 11940 3122 11996
rect 3122 11940 3126 11996
rect 3062 11936 3126 11940
rect 6564 11996 6628 12000
rect 6564 11940 6568 11996
rect 6568 11940 6624 11996
rect 6624 11940 6628 11996
rect 6564 11936 6628 11940
rect 6644 11996 6708 12000
rect 6644 11940 6648 11996
rect 6648 11940 6704 11996
rect 6704 11940 6708 11996
rect 6644 11936 6708 11940
rect 6724 11996 6788 12000
rect 6724 11940 6728 11996
rect 6728 11940 6784 11996
rect 6784 11940 6788 11996
rect 6724 11936 6788 11940
rect 6804 11996 6868 12000
rect 6804 11940 6808 11996
rect 6808 11940 6864 11996
rect 6864 11940 6868 11996
rect 6804 11936 6868 11940
rect 10305 11996 10369 12000
rect 10305 11940 10309 11996
rect 10309 11940 10365 11996
rect 10365 11940 10369 11996
rect 10305 11936 10369 11940
rect 10385 11996 10449 12000
rect 10385 11940 10389 11996
rect 10389 11940 10445 11996
rect 10445 11940 10449 11996
rect 10385 11936 10449 11940
rect 10465 11996 10529 12000
rect 10465 11940 10469 11996
rect 10469 11940 10525 11996
rect 10525 11940 10529 11996
rect 10465 11936 10529 11940
rect 10545 11996 10609 12000
rect 10545 11940 10549 11996
rect 10549 11940 10605 11996
rect 10605 11940 10609 11996
rect 10545 11936 10609 11940
rect 4693 11452 4757 11456
rect 4693 11396 4697 11452
rect 4697 11396 4753 11452
rect 4753 11396 4757 11452
rect 4693 11392 4757 11396
rect 4773 11452 4837 11456
rect 4773 11396 4777 11452
rect 4777 11396 4833 11452
rect 4833 11396 4837 11452
rect 4773 11392 4837 11396
rect 4853 11452 4917 11456
rect 4853 11396 4857 11452
rect 4857 11396 4913 11452
rect 4913 11396 4917 11452
rect 4853 11392 4917 11396
rect 4933 11452 4997 11456
rect 4933 11396 4937 11452
rect 4937 11396 4993 11452
rect 4993 11396 4997 11452
rect 4933 11392 4997 11396
rect 8434 11452 8498 11456
rect 8434 11396 8438 11452
rect 8438 11396 8494 11452
rect 8494 11396 8498 11452
rect 8434 11392 8498 11396
rect 8514 11452 8578 11456
rect 8514 11396 8518 11452
rect 8518 11396 8574 11452
rect 8574 11396 8578 11452
rect 8514 11392 8578 11396
rect 8594 11452 8658 11456
rect 8594 11396 8598 11452
rect 8598 11396 8654 11452
rect 8654 11396 8658 11452
rect 8594 11392 8658 11396
rect 8674 11452 8738 11456
rect 8674 11396 8678 11452
rect 8678 11396 8734 11452
rect 8734 11396 8738 11452
rect 8674 11392 8738 11396
rect 5580 11248 5644 11252
rect 5580 11192 5630 11248
rect 5630 11192 5644 11248
rect 5580 11188 5644 11192
rect 980 11052 1044 11116
rect 5764 11112 5828 11116
rect 5764 11056 5778 11112
rect 5778 11056 5828 11112
rect 5764 11052 5828 11056
rect 7052 11052 7116 11116
rect 7604 11112 7668 11116
rect 7604 11056 7654 11112
rect 7654 11056 7668 11112
rect 7604 11052 7668 11056
rect 2822 10908 2886 10912
rect 2822 10852 2826 10908
rect 2826 10852 2882 10908
rect 2882 10852 2886 10908
rect 2822 10848 2886 10852
rect 2902 10908 2966 10912
rect 2902 10852 2906 10908
rect 2906 10852 2962 10908
rect 2962 10852 2966 10908
rect 2902 10848 2966 10852
rect 2982 10908 3046 10912
rect 2982 10852 2986 10908
rect 2986 10852 3042 10908
rect 3042 10852 3046 10908
rect 2982 10848 3046 10852
rect 3062 10908 3126 10912
rect 3062 10852 3066 10908
rect 3066 10852 3122 10908
rect 3122 10852 3126 10908
rect 3062 10848 3126 10852
rect 6564 10908 6628 10912
rect 6564 10852 6568 10908
rect 6568 10852 6624 10908
rect 6624 10852 6628 10908
rect 6564 10848 6628 10852
rect 6644 10908 6708 10912
rect 6644 10852 6648 10908
rect 6648 10852 6704 10908
rect 6704 10852 6708 10908
rect 6644 10848 6708 10852
rect 6724 10908 6788 10912
rect 6724 10852 6728 10908
rect 6728 10852 6784 10908
rect 6784 10852 6788 10908
rect 6724 10848 6788 10852
rect 6804 10908 6868 10912
rect 6804 10852 6808 10908
rect 6808 10852 6864 10908
rect 6864 10852 6868 10908
rect 6804 10848 6868 10852
rect 10305 10908 10369 10912
rect 10305 10852 10309 10908
rect 10309 10852 10365 10908
rect 10365 10852 10369 10908
rect 10305 10848 10369 10852
rect 10385 10908 10449 10912
rect 10385 10852 10389 10908
rect 10389 10852 10445 10908
rect 10445 10852 10449 10908
rect 10385 10848 10449 10852
rect 10465 10908 10529 10912
rect 10465 10852 10469 10908
rect 10469 10852 10525 10908
rect 10525 10852 10529 10908
rect 10465 10848 10529 10852
rect 10545 10908 10609 10912
rect 10545 10852 10549 10908
rect 10549 10852 10605 10908
rect 10605 10852 10609 10908
rect 10545 10848 10609 10852
rect 5212 10780 5276 10844
rect 5396 10840 5460 10844
rect 5396 10784 5410 10840
rect 5410 10784 5460 10840
rect 5396 10780 5460 10784
rect 7972 10644 8036 10708
rect 4693 10364 4757 10368
rect 4693 10308 4697 10364
rect 4697 10308 4753 10364
rect 4753 10308 4757 10364
rect 4693 10304 4757 10308
rect 4773 10364 4837 10368
rect 4773 10308 4777 10364
rect 4777 10308 4833 10364
rect 4833 10308 4837 10364
rect 4773 10304 4837 10308
rect 4853 10364 4917 10368
rect 4853 10308 4857 10364
rect 4857 10308 4913 10364
rect 4913 10308 4917 10364
rect 4853 10304 4917 10308
rect 4933 10364 4997 10368
rect 4933 10308 4937 10364
rect 4937 10308 4993 10364
rect 4993 10308 4997 10364
rect 4933 10304 4997 10308
rect 8434 10364 8498 10368
rect 8434 10308 8438 10364
rect 8438 10308 8494 10364
rect 8494 10308 8498 10364
rect 8434 10304 8498 10308
rect 8514 10364 8578 10368
rect 8514 10308 8518 10364
rect 8518 10308 8574 10364
rect 8574 10308 8578 10364
rect 8514 10304 8578 10308
rect 8594 10364 8658 10368
rect 8594 10308 8598 10364
rect 8598 10308 8654 10364
rect 8654 10308 8658 10364
rect 8594 10304 8658 10308
rect 8674 10364 8738 10368
rect 8674 10308 8678 10364
rect 8678 10308 8734 10364
rect 8734 10308 8738 10364
rect 8674 10304 8738 10308
rect 5212 10236 5276 10300
rect 7236 9964 7300 10028
rect 2822 9820 2886 9824
rect 2822 9764 2826 9820
rect 2826 9764 2882 9820
rect 2882 9764 2886 9820
rect 2822 9760 2886 9764
rect 2902 9820 2966 9824
rect 2902 9764 2906 9820
rect 2906 9764 2962 9820
rect 2962 9764 2966 9820
rect 2902 9760 2966 9764
rect 2982 9820 3046 9824
rect 2982 9764 2986 9820
rect 2986 9764 3042 9820
rect 3042 9764 3046 9820
rect 2982 9760 3046 9764
rect 3062 9820 3126 9824
rect 3062 9764 3066 9820
rect 3066 9764 3122 9820
rect 3122 9764 3126 9820
rect 3062 9760 3126 9764
rect 6564 9820 6628 9824
rect 6564 9764 6568 9820
rect 6568 9764 6624 9820
rect 6624 9764 6628 9820
rect 6564 9760 6628 9764
rect 6644 9820 6708 9824
rect 6644 9764 6648 9820
rect 6648 9764 6704 9820
rect 6704 9764 6708 9820
rect 6644 9760 6708 9764
rect 6724 9820 6788 9824
rect 6724 9764 6728 9820
rect 6728 9764 6784 9820
rect 6784 9764 6788 9820
rect 6724 9760 6788 9764
rect 6804 9820 6868 9824
rect 6804 9764 6808 9820
rect 6808 9764 6864 9820
rect 6864 9764 6868 9820
rect 6804 9760 6868 9764
rect 10305 9820 10369 9824
rect 10305 9764 10309 9820
rect 10309 9764 10365 9820
rect 10365 9764 10369 9820
rect 10305 9760 10369 9764
rect 10385 9820 10449 9824
rect 10385 9764 10389 9820
rect 10389 9764 10445 9820
rect 10445 9764 10449 9820
rect 10385 9760 10449 9764
rect 10465 9820 10529 9824
rect 10465 9764 10469 9820
rect 10469 9764 10525 9820
rect 10525 9764 10529 9820
rect 10465 9760 10529 9764
rect 10545 9820 10609 9824
rect 10545 9764 10549 9820
rect 10549 9764 10605 9820
rect 10605 9764 10609 9820
rect 10545 9760 10609 9764
rect 6316 9692 6380 9756
rect 3372 9556 3436 9620
rect 9628 9556 9692 9620
rect 4476 9420 4540 9484
rect 4292 9344 4356 9348
rect 4292 9288 4306 9344
rect 4306 9288 4356 9344
rect 4292 9284 4356 9288
rect 4693 9276 4757 9280
rect 4693 9220 4697 9276
rect 4697 9220 4753 9276
rect 4753 9220 4757 9276
rect 4693 9216 4757 9220
rect 4773 9276 4837 9280
rect 4773 9220 4777 9276
rect 4777 9220 4833 9276
rect 4833 9220 4837 9276
rect 4773 9216 4837 9220
rect 4853 9276 4917 9280
rect 4853 9220 4857 9276
rect 4857 9220 4913 9276
rect 4913 9220 4917 9276
rect 4853 9216 4917 9220
rect 4933 9276 4997 9280
rect 4933 9220 4937 9276
rect 4937 9220 4993 9276
rect 4993 9220 4997 9276
rect 4933 9216 4997 9220
rect 8434 9276 8498 9280
rect 8434 9220 8438 9276
rect 8438 9220 8494 9276
rect 8494 9220 8498 9276
rect 8434 9216 8498 9220
rect 8514 9276 8578 9280
rect 8514 9220 8518 9276
rect 8518 9220 8574 9276
rect 8574 9220 8578 9276
rect 8514 9216 8578 9220
rect 8594 9276 8658 9280
rect 8594 9220 8598 9276
rect 8598 9220 8654 9276
rect 8654 9220 8658 9276
rect 8594 9216 8658 9220
rect 8674 9276 8738 9280
rect 8674 9220 8678 9276
rect 8678 9220 8734 9276
rect 8734 9220 8738 9276
rect 8674 9216 8738 9220
rect 6132 9012 6196 9076
rect 9444 8876 9508 8940
rect 2822 8732 2886 8736
rect 2822 8676 2826 8732
rect 2826 8676 2882 8732
rect 2882 8676 2886 8732
rect 2822 8672 2886 8676
rect 2902 8732 2966 8736
rect 2902 8676 2906 8732
rect 2906 8676 2962 8732
rect 2962 8676 2966 8732
rect 2902 8672 2966 8676
rect 2982 8732 3046 8736
rect 2982 8676 2986 8732
rect 2986 8676 3042 8732
rect 3042 8676 3046 8732
rect 2982 8672 3046 8676
rect 3062 8732 3126 8736
rect 3062 8676 3066 8732
rect 3066 8676 3122 8732
rect 3122 8676 3126 8732
rect 3062 8672 3126 8676
rect 6564 8732 6628 8736
rect 6564 8676 6568 8732
rect 6568 8676 6624 8732
rect 6624 8676 6628 8732
rect 6564 8672 6628 8676
rect 6644 8732 6708 8736
rect 6644 8676 6648 8732
rect 6648 8676 6704 8732
rect 6704 8676 6708 8732
rect 6644 8672 6708 8676
rect 6724 8732 6788 8736
rect 6724 8676 6728 8732
rect 6728 8676 6784 8732
rect 6784 8676 6788 8732
rect 6724 8672 6788 8676
rect 6804 8732 6868 8736
rect 6804 8676 6808 8732
rect 6808 8676 6864 8732
rect 6864 8676 6868 8732
rect 6804 8672 6868 8676
rect 10305 8732 10369 8736
rect 10305 8676 10309 8732
rect 10309 8676 10365 8732
rect 10365 8676 10369 8732
rect 10305 8672 10369 8676
rect 10385 8732 10449 8736
rect 10385 8676 10389 8732
rect 10389 8676 10445 8732
rect 10445 8676 10449 8732
rect 10385 8672 10449 8676
rect 10465 8732 10529 8736
rect 10465 8676 10469 8732
rect 10469 8676 10525 8732
rect 10525 8676 10529 8732
rect 10465 8672 10529 8676
rect 10545 8732 10609 8736
rect 10545 8676 10549 8732
rect 10549 8676 10605 8732
rect 10605 8676 10609 8732
rect 10545 8672 10609 8676
rect 2268 8664 2332 8668
rect 2268 8608 2282 8664
rect 2282 8608 2332 8664
rect 2268 8604 2332 8608
rect 4108 8332 4172 8396
rect 4476 8332 4540 8396
rect 5212 8332 5276 8396
rect 8892 8332 8956 8396
rect 4693 8188 4757 8192
rect 4693 8132 4697 8188
rect 4697 8132 4753 8188
rect 4753 8132 4757 8188
rect 4693 8128 4757 8132
rect 4773 8188 4837 8192
rect 4773 8132 4777 8188
rect 4777 8132 4833 8188
rect 4833 8132 4837 8188
rect 4773 8128 4837 8132
rect 4853 8188 4917 8192
rect 4853 8132 4857 8188
rect 4857 8132 4913 8188
rect 4913 8132 4917 8188
rect 4853 8128 4917 8132
rect 4933 8188 4997 8192
rect 4933 8132 4937 8188
rect 4937 8132 4993 8188
rect 4993 8132 4997 8188
rect 4933 8128 4997 8132
rect 8434 8188 8498 8192
rect 8434 8132 8438 8188
rect 8438 8132 8494 8188
rect 8494 8132 8498 8188
rect 8434 8128 8498 8132
rect 8514 8188 8578 8192
rect 8514 8132 8518 8188
rect 8518 8132 8574 8188
rect 8574 8132 8578 8188
rect 8514 8128 8578 8132
rect 8594 8188 8658 8192
rect 8594 8132 8598 8188
rect 8598 8132 8654 8188
rect 8654 8132 8658 8188
rect 8594 8128 8658 8132
rect 8674 8188 8738 8192
rect 8674 8132 8678 8188
rect 8678 8132 8734 8188
rect 8734 8132 8738 8188
rect 8674 8128 8738 8132
rect 9076 7924 9140 7988
rect 5396 7848 5460 7852
rect 5396 7792 5410 7848
rect 5410 7792 5460 7848
rect 5396 7788 5460 7792
rect 9996 7848 10060 7852
rect 9996 7792 10010 7848
rect 10010 7792 10060 7848
rect 9996 7788 10060 7792
rect 2822 7644 2886 7648
rect 2822 7588 2826 7644
rect 2826 7588 2882 7644
rect 2882 7588 2886 7644
rect 2822 7584 2886 7588
rect 2902 7644 2966 7648
rect 2902 7588 2906 7644
rect 2906 7588 2962 7644
rect 2962 7588 2966 7644
rect 2902 7584 2966 7588
rect 2982 7644 3046 7648
rect 2982 7588 2986 7644
rect 2986 7588 3042 7644
rect 3042 7588 3046 7644
rect 2982 7584 3046 7588
rect 3062 7644 3126 7648
rect 3062 7588 3066 7644
rect 3066 7588 3122 7644
rect 3122 7588 3126 7644
rect 3062 7584 3126 7588
rect 6564 7644 6628 7648
rect 6564 7588 6568 7644
rect 6568 7588 6624 7644
rect 6624 7588 6628 7644
rect 6564 7584 6628 7588
rect 6644 7644 6708 7648
rect 6644 7588 6648 7644
rect 6648 7588 6704 7644
rect 6704 7588 6708 7644
rect 6644 7584 6708 7588
rect 6724 7644 6788 7648
rect 6724 7588 6728 7644
rect 6728 7588 6784 7644
rect 6784 7588 6788 7644
rect 6724 7584 6788 7588
rect 6804 7644 6868 7648
rect 6804 7588 6808 7644
rect 6808 7588 6864 7644
rect 6864 7588 6868 7644
rect 6804 7584 6868 7588
rect 10305 7644 10369 7648
rect 10305 7588 10309 7644
rect 10309 7588 10365 7644
rect 10365 7588 10369 7644
rect 10305 7584 10369 7588
rect 10385 7644 10449 7648
rect 10385 7588 10389 7644
rect 10389 7588 10445 7644
rect 10445 7588 10449 7644
rect 10385 7584 10449 7588
rect 10465 7644 10529 7648
rect 10465 7588 10469 7644
rect 10469 7588 10525 7644
rect 10525 7588 10529 7644
rect 10465 7584 10529 7588
rect 10545 7644 10609 7648
rect 10545 7588 10549 7644
rect 10549 7588 10605 7644
rect 10605 7588 10609 7644
rect 10545 7584 10609 7588
rect 5948 7516 6012 7580
rect 3556 7380 3620 7444
rect 8156 7380 8220 7444
rect 4693 7100 4757 7104
rect 4693 7044 4697 7100
rect 4697 7044 4753 7100
rect 4753 7044 4757 7100
rect 4693 7040 4757 7044
rect 4773 7100 4837 7104
rect 4773 7044 4777 7100
rect 4777 7044 4833 7100
rect 4833 7044 4837 7100
rect 4773 7040 4837 7044
rect 4853 7100 4917 7104
rect 4853 7044 4857 7100
rect 4857 7044 4913 7100
rect 4913 7044 4917 7100
rect 4853 7040 4917 7044
rect 4933 7100 4997 7104
rect 4933 7044 4937 7100
rect 4937 7044 4993 7100
rect 4993 7044 4997 7100
rect 4933 7040 4997 7044
rect 8434 7100 8498 7104
rect 8434 7044 8438 7100
rect 8438 7044 8494 7100
rect 8494 7044 8498 7100
rect 8434 7040 8498 7044
rect 8514 7100 8578 7104
rect 8514 7044 8518 7100
rect 8518 7044 8574 7100
rect 8574 7044 8578 7100
rect 8514 7040 8578 7044
rect 8594 7100 8658 7104
rect 8594 7044 8598 7100
rect 8598 7044 8654 7100
rect 8654 7044 8658 7100
rect 8594 7040 8658 7044
rect 8674 7100 8738 7104
rect 8674 7044 8678 7100
rect 8678 7044 8734 7100
rect 8734 7044 8738 7100
rect 8674 7040 8738 7044
rect 1900 6972 1964 7036
rect 4476 6972 4540 7036
rect 9628 6972 9692 7036
rect 2636 6836 2700 6900
rect 5212 6564 5276 6628
rect 2822 6556 2886 6560
rect 2822 6500 2826 6556
rect 2826 6500 2882 6556
rect 2882 6500 2886 6556
rect 2822 6496 2886 6500
rect 2902 6556 2966 6560
rect 2902 6500 2906 6556
rect 2906 6500 2962 6556
rect 2962 6500 2966 6556
rect 2902 6496 2966 6500
rect 2982 6556 3046 6560
rect 2982 6500 2986 6556
rect 2986 6500 3042 6556
rect 3042 6500 3046 6556
rect 2982 6496 3046 6500
rect 3062 6556 3126 6560
rect 3062 6500 3066 6556
rect 3066 6500 3122 6556
rect 3122 6500 3126 6556
rect 3062 6496 3126 6500
rect 6564 6556 6628 6560
rect 6564 6500 6568 6556
rect 6568 6500 6624 6556
rect 6624 6500 6628 6556
rect 6564 6496 6628 6500
rect 6644 6556 6708 6560
rect 6644 6500 6648 6556
rect 6648 6500 6704 6556
rect 6704 6500 6708 6556
rect 6644 6496 6708 6500
rect 6724 6556 6788 6560
rect 6724 6500 6728 6556
rect 6728 6500 6784 6556
rect 6784 6500 6788 6556
rect 6724 6496 6788 6500
rect 6804 6556 6868 6560
rect 6804 6500 6808 6556
rect 6808 6500 6864 6556
rect 6864 6500 6868 6556
rect 6804 6496 6868 6500
rect 10305 6556 10369 6560
rect 10305 6500 10309 6556
rect 10309 6500 10365 6556
rect 10365 6500 10369 6556
rect 10305 6496 10369 6500
rect 10385 6556 10449 6560
rect 10385 6500 10389 6556
rect 10389 6500 10445 6556
rect 10445 6500 10449 6556
rect 10385 6496 10449 6500
rect 10465 6556 10529 6560
rect 10465 6500 10469 6556
rect 10469 6500 10525 6556
rect 10525 6500 10529 6556
rect 10465 6496 10529 6500
rect 10545 6556 10609 6560
rect 10545 6500 10549 6556
rect 10549 6500 10605 6556
rect 10605 6500 10609 6556
rect 10545 6496 10609 6500
rect 5396 6428 5460 6492
rect 5212 6156 5276 6220
rect 3924 6020 3988 6084
rect 4693 6012 4757 6016
rect 4693 5956 4697 6012
rect 4697 5956 4753 6012
rect 4753 5956 4757 6012
rect 4693 5952 4757 5956
rect 4773 6012 4837 6016
rect 4773 5956 4777 6012
rect 4777 5956 4833 6012
rect 4833 5956 4837 6012
rect 4773 5952 4837 5956
rect 4853 6012 4917 6016
rect 4853 5956 4857 6012
rect 4857 5956 4913 6012
rect 4913 5956 4917 6012
rect 4853 5952 4917 5956
rect 4933 6012 4997 6016
rect 4933 5956 4937 6012
rect 4937 5956 4993 6012
rect 4993 5956 4997 6012
rect 4933 5952 4997 5956
rect 8434 6012 8498 6016
rect 8434 5956 8438 6012
rect 8438 5956 8494 6012
rect 8494 5956 8498 6012
rect 8434 5952 8498 5956
rect 8514 6012 8578 6016
rect 8514 5956 8518 6012
rect 8518 5956 8574 6012
rect 8574 5956 8578 6012
rect 8514 5952 8578 5956
rect 8594 6012 8658 6016
rect 8594 5956 8598 6012
rect 8598 5956 8654 6012
rect 8654 5956 8658 6012
rect 8594 5952 8658 5956
rect 8674 6012 8738 6016
rect 8674 5956 8678 6012
rect 8678 5956 8734 6012
rect 8734 5956 8738 6012
rect 8674 5952 8738 5956
rect 7788 5748 7852 5812
rect 7420 5612 7484 5676
rect 9812 5612 9876 5676
rect 2822 5468 2886 5472
rect 2822 5412 2826 5468
rect 2826 5412 2882 5468
rect 2882 5412 2886 5468
rect 2822 5408 2886 5412
rect 2902 5468 2966 5472
rect 2902 5412 2906 5468
rect 2906 5412 2962 5468
rect 2962 5412 2966 5468
rect 2902 5408 2966 5412
rect 2982 5468 3046 5472
rect 2982 5412 2986 5468
rect 2986 5412 3042 5468
rect 3042 5412 3046 5468
rect 2982 5408 3046 5412
rect 3062 5468 3126 5472
rect 3062 5412 3066 5468
rect 3066 5412 3122 5468
rect 3122 5412 3126 5468
rect 3062 5408 3126 5412
rect 6564 5468 6628 5472
rect 6564 5412 6568 5468
rect 6568 5412 6624 5468
rect 6624 5412 6628 5468
rect 6564 5408 6628 5412
rect 6644 5468 6708 5472
rect 6644 5412 6648 5468
rect 6648 5412 6704 5468
rect 6704 5412 6708 5468
rect 6644 5408 6708 5412
rect 6724 5468 6788 5472
rect 6724 5412 6728 5468
rect 6728 5412 6784 5468
rect 6784 5412 6788 5468
rect 6724 5408 6788 5412
rect 6804 5468 6868 5472
rect 6804 5412 6808 5468
rect 6808 5412 6864 5468
rect 6864 5412 6868 5468
rect 6804 5408 6868 5412
rect 10305 5468 10369 5472
rect 10305 5412 10309 5468
rect 10309 5412 10365 5468
rect 10365 5412 10369 5468
rect 10305 5408 10369 5412
rect 10385 5468 10449 5472
rect 10385 5412 10389 5468
rect 10389 5412 10445 5468
rect 10445 5412 10449 5468
rect 10385 5408 10449 5412
rect 10465 5468 10529 5472
rect 10465 5412 10469 5468
rect 10469 5412 10525 5468
rect 10525 5412 10529 5468
rect 10465 5408 10529 5412
rect 10545 5468 10609 5472
rect 10545 5412 10549 5468
rect 10549 5412 10605 5468
rect 10605 5412 10609 5468
rect 10545 5408 10609 5412
rect 5948 5400 6012 5404
rect 5948 5344 5998 5400
rect 5998 5344 6012 5400
rect 5948 5340 6012 5344
rect 5948 5068 6012 5132
rect 7972 5204 8036 5268
rect 5396 4932 5460 4996
rect 7972 4932 8036 4996
rect 4693 4924 4757 4928
rect 4693 4868 4697 4924
rect 4697 4868 4753 4924
rect 4753 4868 4757 4924
rect 4693 4864 4757 4868
rect 4773 4924 4837 4928
rect 4773 4868 4777 4924
rect 4777 4868 4833 4924
rect 4833 4868 4837 4924
rect 4773 4864 4837 4868
rect 4853 4924 4917 4928
rect 4853 4868 4857 4924
rect 4857 4868 4913 4924
rect 4913 4868 4917 4924
rect 4853 4864 4917 4868
rect 4933 4924 4997 4928
rect 4933 4868 4937 4924
rect 4937 4868 4993 4924
rect 4993 4868 4997 4924
rect 4933 4864 4997 4868
rect 8434 4924 8498 4928
rect 8434 4868 8438 4924
rect 8438 4868 8494 4924
rect 8494 4868 8498 4924
rect 8434 4864 8498 4868
rect 8514 4924 8578 4928
rect 8514 4868 8518 4924
rect 8518 4868 8574 4924
rect 8574 4868 8578 4924
rect 8514 4864 8578 4868
rect 8594 4924 8658 4928
rect 8594 4868 8598 4924
rect 8598 4868 8654 4924
rect 8654 4868 8658 4924
rect 8594 4864 8658 4868
rect 8674 4924 8738 4928
rect 8674 4868 8678 4924
rect 8678 4868 8734 4924
rect 8734 4868 8738 4924
rect 8674 4864 8738 4868
rect 9444 4856 9508 4860
rect 9444 4800 9494 4856
rect 9494 4800 9508 4856
rect 9444 4796 9508 4800
rect 5396 4660 5460 4724
rect 10916 4660 10980 4724
rect 3740 4524 3804 4588
rect 2822 4380 2886 4384
rect 2822 4324 2826 4380
rect 2826 4324 2882 4380
rect 2882 4324 2886 4380
rect 2822 4320 2886 4324
rect 2902 4380 2966 4384
rect 2902 4324 2906 4380
rect 2906 4324 2962 4380
rect 2962 4324 2966 4380
rect 2902 4320 2966 4324
rect 2982 4380 3046 4384
rect 2982 4324 2986 4380
rect 2986 4324 3042 4380
rect 3042 4324 3046 4380
rect 2982 4320 3046 4324
rect 3062 4380 3126 4384
rect 3062 4324 3066 4380
rect 3066 4324 3122 4380
rect 3122 4324 3126 4380
rect 3062 4320 3126 4324
rect 6564 4380 6628 4384
rect 6564 4324 6568 4380
rect 6568 4324 6624 4380
rect 6624 4324 6628 4380
rect 6564 4320 6628 4324
rect 6644 4380 6708 4384
rect 6644 4324 6648 4380
rect 6648 4324 6704 4380
rect 6704 4324 6708 4380
rect 6644 4320 6708 4324
rect 6724 4380 6788 4384
rect 6724 4324 6728 4380
rect 6728 4324 6784 4380
rect 6784 4324 6788 4380
rect 6724 4320 6788 4324
rect 6804 4380 6868 4384
rect 6804 4324 6808 4380
rect 6808 4324 6864 4380
rect 6864 4324 6868 4380
rect 6804 4320 6868 4324
rect 10305 4380 10369 4384
rect 10305 4324 10309 4380
rect 10309 4324 10365 4380
rect 10365 4324 10369 4380
rect 10305 4320 10369 4324
rect 10385 4380 10449 4384
rect 10385 4324 10389 4380
rect 10389 4324 10445 4380
rect 10445 4324 10449 4380
rect 10385 4320 10449 4324
rect 10465 4380 10529 4384
rect 10465 4324 10469 4380
rect 10469 4324 10525 4380
rect 10525 4324 10529 4380
rect 10465 4320 10529 4324
rect 10545 4380 10609 4384
rect 10545 4324 10549 4380
rect 10549 4324 10605 4380
rect 10605 4324 10609 4380
rect 10545 4320 10609 4324
rect 3924 4252 3988 4316
rect 3924 4116 3988 4180
rect 5580 4116 5644 4180
rect 9260 4116 9324 4180
rect 980 3980 1044 4044
rect 4693 3836 4757 3840
rect 4693 3780 4697 3836
rect 4697 3780 4753 3836
rect 4753 3780 4757 3836
rect 4693 3776 4757 3780
rect 4773 3836 4837 3840
rect 4773 3780 4777 3836
rect 4777 3780 4833 3836
rect 4833 3780 4837 3836
rect 4773 3776 4837 3780
rect 4853 3836 4917 3840
rect 4853 3780 4857 3836
rect 4857 3780 4913 3836
rect 4913 3780 4917 3836
rect 4853 3776 4917 3780
rect 4933 3836 4997 3840
rect 4933 3780 4937 3836
rect 4937 3780 4993 3836
rect 4993 3780 4997 3836
rect 4933 3776 4997 3780
rect 8434 3836 8498 3840
rect 8434 3780 8438 3836
rect 8438 3780 8494 3836
rect 8494 3780 8498 3836
rect 8434 3776 8498 3780
rect 8514 3836 8578 3840
rect 8514 3780 8518 3836
rect 8518 3780 8574 3836
rect 8574 3780 8578 3836
rect 8514 3776 8578 3780
rect 8594 3836 8658 3840
rect 8594 3780 8598 3836
rect 8598 3780 8654 3836
rect 8654 3780 8658 3836
rect 8594 3776 8658 3780
rect 8674 3836 8738 3840
rect 8674 3780 8678 3836
rect 8678 3780 8734 3836
rect 8734 3780 8738 3836
rect 8674 3776 8738 3780
rect 2084 3572 2148 3636
rect 4292 3436 4356 3500
rect 10916 3436 10980 3500
rect 2822 3292 2886 3296
rect 2822 3236 2826 3292
rect 2826 3236 2882 3292
rect 2882 3236 2886 3292
rect 2822 3232 2886 3236
rect 2902 3292 2966 3296
rect 2902 3236 2906 3292
rect 2906 3236 2962 3292
rect 2962 3236 2966 3292
rect 2902 3232 2966 3236
rect 2982 3292 3046 3296
rect 2982 3236 2986 3292
rect 2986 3236 3042 3292
rect 3042 3236 3046 3292
rect 2982 3232 3046 3236
rect 3062 3292 3126 3296
rect 3062 3236 3066 3292
rect 3066 3236 3122 3292
rect 3122 3236 3126 3292
rect 3062 3232 3126 3236
rect 6564 3292 6628 3296
rect 6564 3236 6568 3292
rect 6568 3236 6624 3292
rect 6624 3236 6628 3292
rect 6564 3232 6628 3236
rect 6644 3292 6708 3296
rect 6644 3236 6648 3292
rect 6648 3236 6704 3292
rect 6704 3236 6708 3292
rect 6644 3232 6708 3236
rect 6724 3292 6788 3296
rect 6724 3236 6728 3292
rect 6728 3236 6784 3292
rect 6784 3236 6788 3292
rect 6724 3232 6788 3236
rect 6804 3292 6868 3296
rect 6804 3236 6808 3292
rect 6808 3236 6864 3292
rect 6864 3236 6868 3292
rect 6804 3232 6868 3236
rect 10305 3292 10369 3296
rect 10305 3236 10309 3292
rect 10309 3236 10365 3292
rect 10365 3236 10369 3292
rect 10305 3232 10369 3236
rect 10385 3292 10449 3296
rect 10385 3236 10389 3292
rect 10389 3236 10445 3292
rect 10445 3236 10449 3292
rect 10385 3232 10449 3236
rect 10465 3292 10529 3296
rect 10465 3236 10469 3292
rect 10469 3236 10525 3292
rect 10525 3236 10529 3292
rect 10465 3232 10529 3236
rect 10545 3292 10609 3296
rect 10545 3236 10549 3292
rect 10549 3236 10605 3292
rect 10605 3236 10609 3292
rect 10545 3232 10609 3236
rect 1716 3224 1780 3228
rect 1716 3168 1766 3224
rect 1766 3168 1780 3224
rect 1716 3164 1780 3168
rect 3372 3028 3436 3092
rect 2452 2892 2516 2956
rect 3556 2892 3620 2956
rect 2268 2816 2332 2820
rect 2268 2760 2318 2816
rect 2318 2760 2332 2816
rect 2268 2756 2332 2760
rect 3924 2892 3988 2956
rect 4108 2952 4172 2956
rect 5580 3088 5644 3092
rect 8892 3164 8956 3228
rect 5580 3032 5594 3088
rect 5594 3032 5644 3088
rect 5580 3028 5644 3032
rect 9996 3088 10060 3092
rect 9996 3032 10046 3088
rect 10046 3032 10060 3088
rect 9996 3028 10060 3032
rect 4108 2896 4158 2952
rect 4158 2896 4172 2952
rect 4108 2892 4172 2896
rect 5396 2892 5460 2956
rect 6316 2892 6380 2956
rect 7604 2892 7668 2956
rect 9812 2892 9876 2956
rect 4693 2748 4757 2752
rect 4693 2692 4697 2748
rect 4697 2692 4753 2748
rect 4753 2692 4757 2748
rect 4693 2688 4757 2692
rect 4773 2748 4837 2752
rect 4773 2692 4777 2748
rect 4777 2692 4833 2748
rect 4833 2692 4837 2748
rect 4773 2688 4837 2692
rect 4853 2748 4917 2752
rect 4853 2692 4857 2748
rect 4857 2692 4913 2748
rect 4913 2692 4917 2748
rect 4853 2688 4917 2692
rect 4933 2748 4997 2752
rect 4933 2692 4937 2748
rect 4937 2692 4993 2748
rect 4993 2692 4997 2748
rect 4933 2688 4997 2692
rect 4108 2620 4172 2684
rect 3740 2484 3804 2548
rect 7788 2756 7852 2820
rect 8434 2748 8498 2752
rect 8434 2692 8438 2748
rect 8438 2692 8494 2748
rect 8494 2692 8498 2748
rect 8434 2688 8498 2692
rect 8514 2748 8578 2752
rect 8514 2692 8518 2748
rect 8518 2692 8574 2748
rect 8574 2692 8578 2748
rect 8514 2688 8578 2692
rect 8594 2748 8658 2752
rect 8594 2692 8598 2748
rect 8598 2692 8654 2748
rect 8654 2692 8658 2748
rect 8594 2688 8658 2692
rect 8674 2748 8738 2752
rect 8674 2692 8678 2748
rect 8678 2692 8734 2748
rect 8734 2692 8738 2748
rect 8674 2688 8738 2692
rect 6132 2620 6196 2684
rect 5948 2484 6012 2548
rect 8156 2484 8220 2548
rect 5212 2348 5276 2412
rect 9076 2348 9140 2412
rect 7420 2212 7484 2276
rect 2822 2204 2886 2208
rect 2822 2148 2826 2204
rect 2826 2148 2882 2204
rect 2882 2148 2886 2204
rect 2822 2144 2886 2148
rect 2902 2204 2966 2208
rect 2902 2148 2906 2204
rect 2906 2148 2962 2204
rect 2962 2148 2966 2204
rect 2902 2144 2966 2148
rect 2982 2204 3046 2208
rect 2982 2148 2986 2204
rect 2986 2148 3042 2204
rect 3042 2148 3046 2204
rect 2982 2144 3046 2148
rect 3062 2204 3126 2208
rect 3062 2148 3066 2204
rect 3066 2148 3122 2204
rect 3122 2148 3126 2204
rect 3062 2144 3126 2148
rect 6564 2204 6628 2208
rect 6564 2148 6568 2204
rect 6568 2148 6624 2204
rect 6624 2148 6628 2204
rect 6564 2144 6628 2148
rect 6644 2204 6708 2208
rect 6644 2148 6648 2204
rect 6648 2148 6704 2204
rect 6704 2148 6708 2204
rect 6644 2144 6708 2148
rect 6724 2204 6788 2208
rect 6724 2148 6728 2204
rect 6728 2148 6784 2204
rect 6784 2148 6788 2204
rect 6724 2144 6788 2148
rect 6804 2204 6868 2208
rect 6804 2148 6808 2204
rect 6808 2148 6864 2204
rect 6864 2148 6868 2204
rect 6804 2144 6868 2148
rect 10305 2204 10369 2208
rect 10305 2148 10309 2204
rect 10309 2148 10365 2204
rect 10365 2148 10369 2204
rect 10305 2144 10369 2148
rect 10385 2204 10449 2208
rect 10385 2148 10389 2204
rect 10389 2148 10445 2204
rect 10445 2148 10449 2204
rect 10385 2144 10449 2148
rect 10465 2204 10529 2208
rect 10465 2148 10469 2204
rect 10469 2148 10525 2204
rect 10525 2148 10529 2204
rect 10465 2144 10529 2148
rect 10545 2204 10609 2208
rect 10545 2148 10549 2204
rect 10549 2148 10605 2204
rect 10605 2148 10609 2204
rect 10545 2144 10609 2148
rect 5396 1940 5460 2004
rect 2636 1864 2700 1868
rect 2636 1808 2650 1864
rect 2650 1808 2700 1864
rect 2636 1804 2700 1808
rect 7052 1804 7116 1868
rect 1716 1668 1780 1732
rect 7972 1668 8036 1732
rect 1900 1532 1964 1596
rect 5764 1396 5828 1460
rect 4476 1260 4540 1324
rect 9260 1260 9324 1324
rect 7236 1124 7300 1188
rect 4292 988 4356 1052
<< metal4 >>
rect 2814 13088 3135 13104
rect 2814 13024 2822 13088
rect 2886 13024 2902 13088
rect 2966 13024 2982 13088
rect 3046 13024 3062 13088
rect 3126 13024 3135 13088
rect 2083 12612 2149 12613
rect 2083 12548 2084 12612
rect 2148 12548 2149 12612
rect 2083 12547 2149 12548
rect 2451 12612 2517 12613
rect 2451 12548 2452 12612
rect 2516 12548 2517 12612
rect 2451 12547 2517 12548
rect 979 11116 1045 11117
rect 979 11052 980 11116
rect 1044 11052 1045 11116
rect 979 11051 1045 11052
rect 982 4045 1042 11051
rect 1899 7036 1965 7037
rect 1899 6972 1900 7036
rect 1964 6972 1965 7036
rect 1899 6971 1965 6972
rect 979 4044 1045 4045
rect 979 3980 980 4044
rect 1044 3980 1045 4044
rect 979 3979 1045 3980
rect 1715 3228 1781 3229
rect 1715 3164 1716 3228
rect 1780 3164 1781 3228
rect 1715 3163 1781 3164
rect 1718 1733 1778 3163
rect 1715 1732 1781 1733
rect 1715 1668 1716 1732
rect 1780 1668 1781 1732
rect 1715 1667 1781 1668
rect 1902 1597 1962 6971
rect 2086 3637 2146 12547
rect 2267 8668 2333 8669
rect 2267 8604 2268 8668
rect 2332 8604 2333 8668
rect 2267 8603 2333 8604
rect 2083 3636 2149 3637
rect 2083 3572 2084 3636
rect 2148 3572 2149 3636
rect 2083 3571 2149 3572
rect 2270 2821 2330 8603
rect 2454 2957 2514 12547
rect 2814 12000 3135 13024
rect 2814 11936 2822 12000
rect 2886 11936 2902 12000
rect 2966 11936 2982 12000
rect 3046 11936 3062 12000
rect 3126 11936 3135 12000
rect 2814 11312 3135 11936
rect 2814 11076 2856 11312
rect 3092 11076 3135 11312
rect 2814 10912 3135 11076
rect 2814 10848 2822 10912
rect 2886 10848 2902 10912
rect 2966 10848 2982 10912
rect 3046 10848 3062 10912
rect 3126 10848 3135 10912
rect 2814 9824 3135 10848
rect 2814 9760 2822 9824
rect 2886 9760 2902 9824
rect 2966 9760 2982 9824
rect 3046 9760 3062 9824
rect 3126 9760 3135 9824
rect 2814 8736 3135 9760
rect 4685 12544 5005 13104
rect 4685 12480 4693 12544
rect 4757 12480 4773 12544
rect 4837 12480 4853 12544
rect 4917 12480 4933 12544
rect 4997 12480 5005 12544
rect 4685 11456 5005 12480
rect 4685 11392 4693 11456
rect 4757 11392 4773 11456
rect 4837 11392 4853 11456
rect 4917 11392 4933 11456
rect 4997 11392 5005 11456
rect 4685 10368 5005 11392
rect 6556 13088 6876 13104
rect 6556 13024 6564 13088
rect 6628 13024 6644 13088
rect 6708 13024 6724 13088
rect 6788 13024 6804 13088
rect 6868 13024 6876 13088
rect 6556 12000 6876 13024
rect 6556 11936 6564 12000
rect 6628 11936 6644 12000
rect 6708 11936 6724 12000
rect 6788 11936 6804 12000
rect 6868 11936 6876 12000
rect 6556 11312 6876 11936
rect 5579 11252 5645 11253
rect 5579 11188 5580 11252
rect 5644 11188 5645 11252
rect 5579 11187 5645 11188
rect 5211 10844 5277 10845
rect 5211 10780 5212 10844
rect 5276 10780 5277 10844
rect 5211 10779 5277 10780
rect 5395 10844 5461 10845
rect 5395 10780 5396 10844
rect 5460 10780 5461 10844
rect 5395 10779 5461 10780
rect 4685 10304 4693 10368
rect 4757 10304 4773 10368
rect 4837 10304 4853 10368
rect 4917 10304 4933 10368
rect 4997 10304 5005 10368
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 2814 8672 2822 8736
rect 2886 8672 2902 8736
rect 2966 8672 2982 8736
rect 3046 8672 3062 8736
rect 3126 8672 3135 8736
rect 2814 7686 3135 8672
rect 2814 7648 2856 7686
rect 3092 7648 3135 7686
rect 2814 7584 2822 7648
rect 3126 7584 3135 7648
rect 2814 7450 2856 7584
rect 3092 7450 3135 7584
rect 2635 6900 2701 6901
rect 2635 6836 2636 6900
rect 2700 6836 2701 6900
rect 2635 6835 2701 6836
rect 2451 2956 2517 2957
rect 2451 2892 2452 2956
rect 2516 2892 2517 2956
rect 2451 2891 2517 2892
rect 2267 2820 2333 2821
rect 2267 2756 2268 2820
rect 2332 2756 2333 2820
rect 2267 2755 2333 2756
rect 2638 1869 2698 6835
rect 2814 6560 3135 7450
rect 2814 6496 2822 6560
rect 2886 6496 2902 6560
rect 2966 6496 2982 6560
rect 3046 6496 3062 6560
rect 3126 6496 3135 6560
rect 2814 5472 3135 6496
rect 2814 5408 2822 5472
rect 2886 5408 2902 5472
rect 2966 5408 2982 5472
rect 3046 5408 3062 5472
rect 3126 5408 3135 5472
rect 2814 4384 3135 5408
rect 2814 4320 2822 4384
rect 2886 4320 2902 4384
rect 2966 4320 2982 4384
rect 3046 4320 3062 4384
rect 3126 4320 3135 4384
rect 2814 4059 3135 4320
rect 2814 3823 2856 4059
rect 3092 3823 3135 4059
rect 2814 3296 3135 3823
rect 2814 3232 2822 3296
rect 2886 3232 2902 3296
rect 2966 3232 2982 3296
rect 3046 3232 3062 3296
rect 3126 3232 3135 3296
rect 2814 2208 3135 3232
rect 3374 3093 3434 9555
rect 4685 9499 5005 10304
rect 5214 10301 5274 10779
rect 5211 10300 5277 10301
rect 5211 10236 5212 10300
rect 5276 10236 5277 10300
rect 5211 10235 5277 10236
rect 4475 9484 4541 9485
rect 4475 9420 4476 9484
rect 4540 9420 4541 9484
rect 4475 9419 4541 9420
rect 4291 9348 4357 9349
rect 4291 9284 4292 9348
rect 4356 9284 4357 9348
rect 4291 9283 4357 9284
rect 4107 8396 4173 8397
rect 4107 8332 4108 8396
rect 4172 8332 4173 8396
rect 4107 8331 4173 8332
rect 3555 7444 3621 7445
rect 3555 7380 3556 7444
rect 3620 7380 3621 7444
rect 3555 7379 3621 7380
rect 3371 3092 3437 3093
rect 3371 3028 3372 3092
rect 3436 3028 3437 3092
rect 3371 3027 3437 3028
rect 3558 2957 3618 7379
rect 3923 6084 3989 6085
rect 3923 6020 3924 6084
rect 3988 6020 3989 6084
rect 3923 6019 3989 6020
rect 3739 4588 3805 4589
rect 3739 4524 3740 4588
rect 3804 4524 3805 4588
rect 3739 4523 3805 4524
rect 3555 2956 3621 2957
rect 3555 2892 3556 2956
rect 3620 2892 3621 2956
rect 3555 2891 3621 2892
rect 3742 2549 3802 4523
rect 3926 4317 3986 6019
rect 3923 4316 3989 4317
rect 3923 4252 3924 4316
rect 3988 4252 3989 4316
rect 3923 4251 3989 4252
rect 3923 4180 3989 4181
rect 3923 4116 3924 4180
rect 3988 4116 3989 4180
rect 3923 4115 3989 4116
rect 3926 2957 3986 4115
rect 4110 3090 4170 8331
rect 4294 3501 4354 9283
rect 4478 8397 4538 9419
rect 4685 9280 4727 9499
rect 4963 9280 5005 9499
rect 4685 9216 4693 9280
rect 4757 9216 4773 9263
rect 4837 9216 4853 9263
rect 4917 9216 4933 9263
rect 4997 9216 5005 9280
rect 4475 8396 4541 8397
rect 4475 8332 4476 8396
rect 4540 8332 4541 8396
rect 4475 8331 4541 8332
rect 4685 8192 5005 9216
rect 5211 8396 5277 8397
rect 5211 8332 5212 8396
rect 5276 8332 5277 8396
rect 5211 8331 5277 8332
rect 4685 8128 4693 8192
rect 4757 8128 4773 8192
rect 4837 8128 4853 8192
rect 4917 8128 4933 8192
rect 4997 8128 5005 8192
rect 4685 7104 5005 8128
rect 4685 7040 4693 7104
rect 4757 7040 4773 7104
rect 4837 7040 4853 7104
rect 4917 7040 4933 7104
rect 4997 7040 5005 7104
rect 4475 7036 4541 7037
rect 4475 6972 4476 7036
rect 4540 6972 4541 7036
rect 4475 6971 4541 6972
rect 4291 3500 4357 3501
rect 4291 3436 4292 3500
rect 4356 3436 4357 3500
rect 4291 3435 4357 3436
rect 4110 3030 4354 3090
rect 3923 2956 3989 2957
rect 3923 2892 3924 2956
rect 3988 2892 3989 2956
rect 3923 2891 3989 2892
rect 4107 2956 4173 2957
rect 4107 2892 4108 2956
rect 4172 2892 4173 2956
rect 4107 2891 4173 2892
rect 4110 2685 4170 2891
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 3739 2548 3805 2549
rect 3739 2484 3740 2548
rect 3804 2484 3805 2548
rect 3739 2483 3805 2484
rect 2814 2144 2822 2208
rect 2886 2144 2902 2208
rect 2966 2144 2982 2208
rect 3046 2144 3062 2208
rect 3126 2144 3135 2208
rect 2814 2128 3135 2144
rect 2635 1868 2701 1869
rect 2635 1804 2636 1868
rect 2700 1804 2701 1868
rect 2635 1803 2701 1804
rect 1899 1596 1965 1597
rect 1899 1532 1900 1596
rect 1964 1532 1965 1596
rect 1899 1531 1965 1532
rect 4294 1053 4354 3030
rect 4478 1325 4538 6971
rect 4685 6016 5005 7040
rect 5214 6629 5274 8331
rect 5398 7853 5458 10779
rect 5395 7852 5461 7853
rect 5395 7788 5396 7852
rect 5460 7788 5461 7852
rect 5395 7787 5461 7788
rect 5211 6628 5277 6629
rect 5211 6564 5212 6628
rect 5276 6564 5277 6628
rect 5211 6563 5277 6564
rect 5395 6492 5461 6493
rect 5395 6428 5396 6492
rect 5460 6428 5461 6492
rect 5395 6427 5461 6428
rect 5211 6220 5277 6221
rect 5211 6156 5212 6220
rect 5276 6156 5277 6220
rect 5211 6155 5277 6156
rect 4685 5952 4693 6016
rect 4757 5952 4773 6016
rect 4837 5952 4853 6016
rect 4917 5952 4933 6016
rect 4997 5952 5005 6016
rect 4685 5872 5005 5952
rect 4685 5636 4727 5872
rect 4963 5636 5005 5872
rect 4685 4928 5005 5636
rect 4685 4864 4693 4928
rect 4757 4864 4773 4928
rect 4837 4864 4853 4928
rect 4917 4864 4933 4928
rect 4997 4864 5005 4928
rect 4685 3840 5005 4864
rect 4685 3776 4693 3840
rect 4757 3776 4773 3840
rect 4837 3776 4853 3840
rect 4917 3776 4933 3840
rect 4997 3776 5005 3840
rect 4685 2752 5005 3776
rect 4685 2688 4693 2752
rect 4757 2688 4773 2752
rect 4837 2688 4853 2752
rect 4917 2688 4933 2752
rect 4997 2688 5005 2752
rect 4685 2128 5005 2688
rect 5214 2413 5274 6155
rect 5398 4997 5458 6427
rect 5395 4996 5461 4997
rect 5395 4932 5396 4996
rect 5460 4932 5461 4996
rect 5395 4931 5461 4932
rect 5395 4724 5461 4725
rect 5395 4660 5396 4724
rect 5460 4660 5461 4724
rect 5395 4659 5461 4660
rect 5398 3090 5458 4659
rect 5582 4181 5642 11187
rect 5763 11116 5829 11117
rect 5763 11052 5764 11116
rect 5828 11052 5829 11116
rect 5763 11051 5829 11052
rect 6556 11076 6598 11312
rect 6834 11076 6876 11312
rect 8426 12544 8747 13104
rect 8426 12480 8434 12544
rect 8498 12480 8514 12544
rect 8578 12480 8594 12544
rect 8658 12480 8674 12544
rect 8738 12480 8747 12544
rect 8426 11456 8747 12480
rect 8426 11392 8434 11456
rect 8498 11392 8514 11456
rect 8578 11392 8594 11456
rect 8658 11392 8674 11456
rect 8738 11392 8747 11456
rect 5579 4180 5645 4181
rect 5579 4116 5580 4180
rect 5644 4116 5645 4180
rect 5579 4115 5645 4116
rect 5579 3092 5645 3093
rect 5579 3090 5580 3092
rect 5398 3030 5580 3090
rect 5579 3028 5580 3030
rect 5644 3028 5645 3092
rect 5579 3027 5645 3028
rect 5395 2956 5461 2957
rect 5395 2892 5396 2956
rect 5460 2892 5461 2956
rect 5395 2891 5461 2892
rect 5211 2412 5277 2413
rect 5211 2348 5212 2412
rect 5276 2348 5277 2412
rect 5211 2347 5277 2348
rect 5398 2005 5458 2891
rect 5395 2004 5461 2005
rect 5395 1940 5396 2004
rect 5460 1940 5461 2004
rect 5395 1939 5461 1940
rect 5766 1461 5826 11051
rect 6556 10912 6876 11076
rect 7051 11116 7117 11117
rect 7051 11052 7052 11116
rect 7116 11052 7117 11116
rect 7051 11051 7117 11052
rect 7603 11116 7669 11117
rect 7603 11052 7604 11116
rect 7668 11052 7669 11116
rect 7603 11051 7669 11052
rect 6556 10848 6564 10912
rect 6628 10848 6644 10912
rect 6708 10848 6724 10912
rect 6788 10848 6804 10912
rect 6868 10848 6876 10912
rect 6556 9824 6876 10848
rect 6556 9760 6564 9824
rect 6628 9760 6644 9824
rect 6708 9760 6724 9824
rect 6788 9760 6804 9824
rect 6868 9760 6876 9824
rect 6315 9756 6381 9757
rect 6315 9692 6316 9756
rect 6380 9692 6381 9756
rect 6315 9691 6381 9692
rect 6131 9076 6197 9077
rect 6131 9012 6132 9076
rect 6196 9012 6197 9076
rect 6131 9011 6197 9012
rect 5947 7580 6013 7581
rect 5947 7516 5948 7580
rect 6012 7516 6013 7580
rect 5947 7515 6013 7516
rect 5950 5405 6010 7515
rect 5947 5404 6013 5405
rect 5947 5340 5948 5404
rect 6012 5340 6013 5404
rect 5947 5339 6013 5340
rect 5947 5132 6013 5133
rect 5947 5068 5948 5132
rect 6012 5068 6013 5132
rect 5947 5067 6013 5068
rect 5950 2549 6010 5067
rect 6134 2685 6194 9011
rect 6318 2957 6378 9691
rect 6556 8736 6876 9760
rect 6556 8672 6564 8736
rect 6628 8672 6644 8736
rect 6708 8672 6724 8736
rect 6788 8672 6804 8736
rect 6868 8672 6876 8736
rect 6556 7686 6876 8672
rect 6556 7648 6598 7686
rect 6834 7648 6876 7686
rect 6556 7584 6564 7648
rect 6868 7584 6876 7648
rect 6556 7450 6598 7584
rect 6834 7450 6876 7584
rect 6556 6560 6876 7450
rect 6556 6496 6564 6560
rect 6628 6496 6644 6560
rect 6708 6496 6724 6560
rect 6788 6496 6804 6560
rect 6868 6496 6876 6560
rect 6556 5472 6876 6496
rect 6556 5408 6564 5472
rect 6628 5408 6644 5472
rect 6708 5408 6724 5472
rect 6788 5408 6804 5472
rect 6868 5408 6876 5472
rect 6556 4384 6876 5408
rect 6556 4320 6564 4384
rect 6628 4320 6644 4384
rect 6708 4320 6724 4384
rect 6788 4320 6804 4384
rect 6868 4320 6876 4384
rect 6556 4059 6876 4320
rect 6556 3823 6598 4059
rect 6834 3823 6876 4059
rect 6556 3296 6876 3823
rect 6556 3232 6564 3296
rect 6628 3232 6644 3296
rect 6708 3232 6724 3296
rect 6788 3232 6804 3296
rect 6868 3232 6876 3296
rect 6315 2956 6381 2957
rect 6315 2892 6316 2956
rect 6380 2892 6381 2956
rect 6315 2891 6381 2892
rect 6131 2684 6197 2685
rect 6131 2620 6132 2684
rect 6196 2620 6197 2684
rect 6131 2619 6197 2620
rect 5947 2548 6013 2549
rect 5947 2484 5948 2548
rect 6012 2484 6013 2548
rect 5947 2483 6013 2484
rect 6556 2208 6876 3232
rect 6556 2144 6564 2208
rect 6628 2144 6644 2208
rect 6708 2144 6724 2208
rect 6788 2144 6804 2208
rect 6868 2144 6876 2208
rect 6556 2128 6876 2144
rect 7054 1869 7114 11051
rect 7235 10028 7301 10029
rect 7235 9964 7236 10028
rect 7300 9964 7301 10028
rect 7235 9963 7301 9964
rect 7051 1868 7117 1869
rect 7051 1804 7052 1868
rect 7116 1804 7117 1868
rect 7051 1803 7117 1804
rect 5763 1460 5829 1461
rect 5763 1396 5764 1460
rect 5828 1396 5829 1460
rect 5763 1395 5829 1396
rect 4475 1324 4541 1325
rect 4475 1260 4476 1324
rect 4540 1260 4541 1324
rect 4475 1259 4541 1260
rect 7238 1189 7298 9963
rect 7419 5676 7485 5677
rect 7419 5612 7420 5676
rect 7484 5612 7485 5676
rect 7419 5611 7485 5612
rect 7422 2277 7482 5611
rect 7606 2957 7666 11051
rect 7971 10708 8037 10709
rect 7971 10644 7972 10708
rect 8036 10644 8037 10708
rect 7971 10643 8037 10644
rect 7787 5812 7853 5813
rect 7787 5748 7788 5812
rect 7852 5748 7853 5812
rect 7787 5747 7853 5748
rect 7603 2956 7669 2957
rect 7603 2892 7604 2956
rect 7668 2892 7669 2956
rect 7603 2891 7669 2892
rect 7790 2821 7850 5747
rect 7974 5269 8034 10643
rect 8426 10368 8747 11392
rect 8426 10304 8434 10368
rect 8498 10304 8514 10368
rect 8578 10304 8594 10368
rect 8658 10304 8674 10368
rect 8738 10304 8747 10368
rect 8426 9499 8747 10304
rect 10297 13088 10617 13104
rect 10297 13024 10305 13088
rect 10369 13024 10385 13088
rect 10449 13024 10465 13088
rect 10529 13024 10545 13088
rect 10609 13024 10617 13088
rect 10297 12000 10617 13024
rect 10297 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10545 12000
rect 10609 11936 10617 12000
rect 10297 11312 10617 11936
rect 10297 11076 10339 11312
rect 10575 11076 10617 11312
rect 10297 10912 10617 11076
rect 10297 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10545 10912
rect 10609 10848 10617 10912
rect 10297 9824 10617 10848
rect 10297 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10545 9824
rect 10609 9760 10617 9824
rect 9627 9620 9693 9621
rect 9627 9556 9628 9620
rect 9692 9556 9693 9620
rect 9627 9555 9693 9556
rect 8426 9280 8468 9499
rect 8704 9280 8747 9499
rect 8426 9216 8434 9280
rect 8498 9216 8514 9263
rect 8578 9216 8594 9263
rect 8658 9216 8674 9263
rect 8738 9216 8747 9280
rect 8426 8192 8747 9216
rect 9443 8940 9509 8941
rect 9443 8876 9444 8940
rect 9508 8876 9509 8940
rect 9443 8875 9509 8876
rect 8891 8396 8957 8397
rect 8891 8332 8892 8396
rect 8956 8332 8957 8396
rect 8891 8331 8957 8332
rect 8426 8128 8434 8192
rect 8498 8128 8514 8192
rect 8578 8128 8594 8192
rect 8658 8128 8674 8192
rect 8738 8128 8747 8192
rect 8155 7444 8221 7445
rect 8155 7380 8156 7444
rect 8220 7380 8221 7444
rect 8155 7379 8221 7380
rect 7971 5268 8037 5269
rect 7971 5204 7972 5268
rect 8036 5204 8037 5268
rect 7971 5203 8037 5204
rect 7971 4996 8037 4997
rect 7971 4932 7972 4996
rect 8036 4932 8037 4996
rect 7971 4931 8037 4932
rect 7787 2820 7853 2821
rect 7787 2756 7788 2820
rect 7852 2756 7853 2820
rect 7787 2755 7853 2756
rect 7419 2276 7485 2277
rect 7419 2212 7420 2276
rect 7484 2212 7485 2276
rect 7419 2211 7485 2212
rect 7974 1733 8034 4931
rect 8158 2549 8218 7379
rect 8426 7104 8747 8128
rect 8426 7040 8434 7104
rect 8498 7040 8514 7104
rect 8578 7040 8594 7104
rect 8658 7040 8674 7104
rect 8738 7040 8747 7104
rect 8426 6016 8747 7040
rect 8426 5952 8434 6016
rect 8498 5952 8514 6016
rect 8578 5952 8594 6016
rect 8658 5952 8674 6016
rect 8738 5952 8747 6016
rect 8426 5872 8747 5952
rect 8426 5636 8468 5872
rect 8704 5636 8747 5872
rect 8426 4928 8747 5636
rect 8426 4864 8434 4928
rect 8498 4864 8514 4928
rect 8578 4864 8594 4928
rect 8658 4864 8674 4928
rect 8738 4864 8747 4928
rect 8426 3840 8747 4864
rect 8426 3776 8434 3840
rect 8498 3776 8514 3840
rect 8578 3776 8594 3840
rect 8658 3776 8674 3840
rect 8738 3776 8747 3840
rect 8426 2752 8747 3776
rect 8894 3229 8954 8331
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 8891 3228 8957 3229
rect 8891 3164 8892 3228
rect 8956 3164 8957 3228
rect 8891 3163 8957 3164
rect 8426 2688 8434 2752
rect 8498 2688 8514 2752
rect 8578 2688 8594 2752
rect 8658 2688 8674 2752
rect 8738 2688 8747 2752
rect 8155 2548 8221 2549
rect 8155 2484 8156 2548
rect 8220 2484 8221 2548
rect 8155 2483 8221 2484
rect 8426 2128 8747 2688
rect 9078 2413 9138 7923
rect 9446 4861 9506 8875
rect 9630 7037 9690 9555
rect 10297 8736 10617 9760
rect 10297 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10545 8736
rect 10609 8672 10617 8736
rect 9995 7852 10061 7853
rect 9995 7788 9996 7852
rect 10060 7788 10061 7852
rect 9995 7787 10061 7788
rect 9627 7036 9693 7037
rect 9627 6972 9628 7036
rect 9692 6972 9693 7036
rect 9627 6971 9693 6972
rect 9811 5676 9877 5677
rect 9811 5612 9812 5676
rect 9876 5612 9877 5676
rect 9811 5611 9877 5612
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 9259 4180 9325 4181
rect 9259 4116 9260 4180
rect 9324 4116 9325 4180
rect 9259 4115 9325 4116
rect 9075 2412 9141 2413
rect 9075 2348 9076 2412
rect 9140 2348 9141 2412
rect 9075 2347 9141 2348
rect 7971 1732 8037 1733
rect 7971 1668 7972 1732
rect 8036 1668 8037 1732
rect 7971 1667 8037 1668
rect 9262 1325 9322 4115
rect 9814 2957 9874 5611
rect 9998 3093 10058 7787
rect 10297 7686 10617 8672
rect 10297 7648 10339 7686
rect 10575 7648 10617 7686
rect 10297 7584 10305 7648
rect 10609 7584 10617 7648
rect 10297 7450 10339 7584
rect 10575 7450 10617 7584
rect 10297 6560 10617 7450
rect 10297 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10465 6560
rect 10529 6496 10545 6560
rect 10609 6496 10617 6560
rect 10297 5472 10617 6496
rect 10297 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10545 5472
rect 10609 5408 10617 5472
rect 10297 4384 10617 5408
rect 10915 4724 10981 4725
rect 10915 4660 10916 4724
rect 10980 4660 10981 4724
rect 10915 4659 10981 4660
rect 10297 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10545 4384
rect 10609 4320 10617 4384
rect 10297 4059 10617 4320
rect 10297 3823 10339 4059
rect 10575 3823 10617 4059
rect 10297 3296 10617 3823
rect 10918 3501 10978 4659
rect 10915 3500 10981 3501
rect 10915 3436 10916 3500
rect 10980 3436 10981 3500
rect 10915 3435 10981 3436
rect 10297 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10545 3296
rect 10609 3232 10617 3296
rect 9995 3092 10061 3093
rect 9995 3028 9996 3092
rect 10060 3028 10061 3092
rect 9995 3027 10061 3028
rect 9811 2956 9877 2957
rect 9811 2892 9812 2956
rect 9876 2892 9877 2956
rect 9811 2891 9877 2892
rect 10297 2208 10617 3232
rect 10297 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10545 2208
rect 10609 2144 10617 2208
rect 10297 2128 10617 2144
rect 9259 1324 9325 1325
rect 9259 1260 9260 1324
rect 9324 1260 9325 1324
rect 9259 1259 9325 1260
rect 7235 1188 7301 1189
rect 7235 1124 7236 1188
rect 7300 1124 7301 1188
rect 7235 1123 7301 1124
rect 4291 1052 4357 1053
rect 4291 988 4292 1052
rect 4356 988 4357 1052
rect 4291 987 4357 988
<< via4 >>
rect 2856 11076 3092 11312
rect 2856 7648 3092 7686
rect 2856 7584 2886 7648
rect 2886 7584 2902 7648
rect 2902 7584 2966 7648
rect 2966 7584 2982 7648
rect 2982 7584 3046 7648
rect 3046 7584 3062 7648
rect 3062 7584 3092 7648
rect 2856 7450 3092 7584
rect 2856 3823 3092 4059
rect 4727 9280 4963 9499
rect 4727 9263 4757 9280
rect 4757 9263 4773 9280
rect 4773 9263 4837 9280
rect 4837 9263 4853 9280
rect 4853 9263 4917 9280
rect 4917 9263 4933 9280
rect 4933 9263 4963 9280
rect 4727 5636 4963 5872
rect 6598 11076 6834 11312
rect 6598 7648 6834 7686
rect 6598 7584 6628 7648
rect 6628 7584 6644 7648
rect 6644 7584 6708 7648
rect 6708 7584 6724 7648
rect 6724 7584 6788 7648
rect 6788 7584 6804 7648
rect 6804 7584 6834 7648
rect 6598 7450 6834 7584
rect 6598 3823 6834 4059
rect 10339 11076 10575 11312
rect 8468 9280 8704 9499
rect 8468 9263 8498 9280
rect 8498 9263 8514 9280
rect 8514 9263 8578 9280
rect 8578 9263 8594 9280
rect 8594 9263 8658 9280
rect 8658 9263 8674 9280
rect 8674 9263 8704 9280
rect 8468 5636 8704 5872
rect 10339 7648 10575 7686
rect 10339 7584 10369 7648
rect 10369 7584 10385 7648
rect 10385 7584 10449 7648
rect 10449 7584 10465 7648
rect 10465 7584 10529 7648
rect 10529 7584 10545 7648
rect 10545 7584 10575 7648
rect 10339 7450 10575 7584
rect 10339 3823 10575 4059
<< metal5 >>
rect 1104 11312 12328 11355
rect 1104 11076 2856 11312
rect 3092 11076 6598 11312
rect 6834 11076 10339 11312
rect 10575 11076 12328 11312
rect 1104 11034 12328 11076
rect 1104 9499 12328 9541
rect 1104 9263 4727 9499
rect 4963 9263 8468 9499
rect 8704 9263 12328 9499
rect 1104 9221 12328 9263
rect 1104 7686 12328 7728
rect 1104 7450 2856 7686
rect 3092 7450 6598 7686
rect 6834 7450 10339 7686
rect 10575 7450 12328 7686
rect 1104 7408 12328 7450
rect 1104 5872 12328 5915
rect 1104 5636 4727 5872
rect 4963 5636 8468 5872
rect 8704 5636 12328 5872
rect 1104 5594 12328 5636
rect 1104 4059 12328 4101
rect 1104 3823 2856 4059
rect 3092 3823 6598 4059
rect 6834 3823 10339 4059
rect 10575 3823 12328 4059
rect 1104 3781 12328 3823
use sky130_fd_sc_hd__nand3_4  _174_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__a31oi_4  _178_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _364_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1621208567
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1621208567
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1621208567
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _396_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3864 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1621208567
transform 1 0 4784 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 4692 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _250_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 6164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1621208567
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1621208567
transform 1 0 6440 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1621208567
transform 1 0 6532 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1621208567
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1621208567
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1621208567
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1621208567
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1621208567
transform 1 0 7452 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_67 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1621208567
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output103 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1621208567
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1621208567
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _239_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1621208567
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1621208567
transform 1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1621208567
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1621208567
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1621208567
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1621208567
transform 1 0 10304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1621208567
transform 1 0 10212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1621208567
transform 1 0 10672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1621208567
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1621208567
transform 1 0 11040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1621208567
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1621208567
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1621208567
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1621208567
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1621208567
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1621208567
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1621208567
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1621208567
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1621208567
transform -1 0 12328 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1621208567
transform -1 0 12328 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _265_
timestamp 1621208567
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1621208567
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1621208567
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _255_
timestamp 1621208567
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1621208567
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1621208567
transform 1 0 3220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1621208567
transform 1 0 4140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1621208567
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _328_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 4508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1621208567
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1621208567
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1621208567
transform 1 0 6624 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _251_
timestamp 1621208567
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1621208567
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1621208567
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _315_
timestamp 1621208567
transform 1 0 5980 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _316_
timestamp 1621208567
transform 1 0 5704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _241_
timestamp 1621208567
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _313_
timestamp 1621208567
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1621208567
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1621208567
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1621208567
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp 1621208567
transform 1 0 8556 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1621208567
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1621208567
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1621208567
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1621208567
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1621208567
transform 1 0 9476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1621208567
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1621208567
transform -1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1621208567
transform 1 0 11316 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1621208567
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1621208567
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1621208567
transform 1 0 2208 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1621208567
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1621208567
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1621208567
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1621208567
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _258_
timestamp 1621208567
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp 1621208567
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1621208567
transform 1 0 3680 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _247_
timestamp 1621208567
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _248_
timestamp 1621208567
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _317_
timestamp 1621208567
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _322_
timestamp 1621208567
transform 1 0 5796 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _323_
timestamp 1621208567
transform 1 0 5520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1621208567
transform 1 0 5244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1621208567
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_44
timestamp 1621208567
transform 1 0 5152 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1621208567
transform 1 0 7912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1621208567
transform 1 0 7452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _314_
timestamp 1621208567
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1621208567
transform 1 0 8556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1621208567
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1621208567
transform 1 0 7084 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1621208567
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _238_
timestamp 1621208567
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1621208567
transform 1 0 9292 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1621208567
transform -1 0 12328 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1621208567
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1621208567
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1621208567
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1621208567
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_105
timestamp 1621208567
transform 1 0 10764 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1621208567
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1621208567
transform 1 0 2760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _268_
timestamp 1621208567
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1621208567
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1621208567
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1621208567
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp 1621208567
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 1621208567
transform 1 0 3956 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _271_
timestamp 1621208567
transform 1 0 4232 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _338_
timestamp 1621208567
transform 1 0 4508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1621208567
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1621208567
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1621208567
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1621208567
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1621208567
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _236_
timestamp 1621208567
transform 1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1621208567
transform 1 0 5152 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1621208567
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1621208567
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1621208567
transform 1 0 7268 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1621208567
transform 1 0 9108 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1621208567
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1621208567
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1621208567
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1621208567
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1621208567
transform -1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1621208567
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1621208567
transform 1 0 11316 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1621208567
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1621208567
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1621208567
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1621208567
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _263_
timestamp 1621208567
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1621208567
transform 1 0 3128 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_41
timestamp 1621208567
transform 1 0 4876 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1621208567
transform 1 0 4968 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1621208567
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _246_
timestamp 1621208567
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _334_
timestamp 1621208567
transform 1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1621208567
transform 1 0 6532 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1621208567
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1621208567
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _229_
timestamp 1621208567
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 1621208567
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1621208567
transform 1 0 7360 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1621208567
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1621208567
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1621208567
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1621208567
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1621208567
transform 1 0 10120 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1621208567
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1621208567
transform -1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1621208567
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1621208567
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1621208567
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input27 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1621208567
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1621208567
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1621208567
transform 1 0 1748 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _278_
timestamp 1621208567
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1621208567
transform 1 0 1656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1621208567
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1621208567
transform 1 0 2852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1621208567
transform 1 0 2024 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _277_
timestamp 1621208567
transform 1 0 2576 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _272_
timestamp 1621208567
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_24
timestamp 1621208567
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1621208567
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1621208567
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1621208567
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1621208567
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1621208567
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1621208567
transform 1 0 3864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1621208567
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1621208567
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1621208567
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1621208567
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1621208567
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_49
timestamp 1621208567
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1621208567
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1621208567
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1621208567
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1621208567
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1621208567
transform 1 0 4968 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1621208567
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _333_
timestamp 1621208567
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1621208567
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1621208567
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1621208567
transform 1 0 6532 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _212_
timestamp 1621208567
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _213_
timestamp 1621208567
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 1621208567
transform 1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _234_
timestamp 1621208567
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _319_
timestamp 1621208567
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1621208567
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1621208567
transform 1 0 8464 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_75
timestamp 1621208567
transform 1 0 8004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _227_
timestamp 1621208567
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _230_
timestamp 1621208567
transform 1 0 9568 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _231_
timestamp 1621208567
transform 1 0 9844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1621208567
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1621208567
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1621208567
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1621208567
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1621208567
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1621208567
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1621208567
transform 1 0 10764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _318_
timestamp 1621208567
transform 1 0 11132 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _320_
timestamp 1621208567
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1621208567
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1621208567
transform 1 0 11960 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1621208567
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _321_
timestamp 1621208567
transform 1 0 11684 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _226_
timestamp 1621208567
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1621208567
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1621208567
transform -1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1621208567
transform 1 0 2852 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1621208567
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1621208567
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1621208567
transform 1 0 3864 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1621208567
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1621208567
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1621208567
transform 1 0 6808 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1621208567
transform 1 0 5336 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1621208567
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _219_
timestamp 1621208567
transform 1 0 8372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1621208567
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1621208567
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1621208567
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1621208567
transform 1 0 9384 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1621208567
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1621208567
transform 1 0 11040 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1621208567
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1621208567
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1621208567
transform -1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1621208567
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1621208567
transform 1 0 2576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1621208567
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1621208567
transform 1 0 2300 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1621208567
transform 1 0 2024 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1621208567
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1621208567
transform 1 0 1472 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1621208567
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1621208567
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _275_
timestamp 1621208567
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _280_
timestamp 1621208567
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1621208567
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1621208567
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1621208567
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1621208567
transform 1 0 3036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 1621208567
transform 1 0 3312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1621208567
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1621208567
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _208_
timestamp 1621208567
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _209_
timestamp 1621208567
transform 1 0 5060 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1621208567
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1621208567
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 6440 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 1621208567
transform 1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1621208567
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1621208567
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1621208567
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _224_
timestamp 1621208567
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 1621208567
transform 1 0 10120 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _223_
timestamp 1621208567
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1621208567
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1621208567
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1621208567
transform -1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1621208567
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1621208567
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_118
timestamp 1621208567
transform 1 0 11960 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _282_
timestamp 1621208567
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1621208567
transform 1 0 2392 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1621208567
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1621208567
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1621208567
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1621208567
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1621208567
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp 1621208567
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1621208567
transform 1 0 3220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1621208567
transform 1 0 4692 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1621208567
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1621208567
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_22
timestamp 1621208567
transform 1 0 3128 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_34
timestamp 1621208567
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1621208567
transform 1 0 6256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp 1621208567
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1621208567
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1621208567
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _217_
timestamp 1621208567
transform 1 0 6900 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _337_
timestamp 1621208567
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1621208567
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1621208567
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1621208567
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp 1621208567
transform 1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _221_
timestamp 1621208567
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _331_
timestamp 1621208567
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _336_
timestamp 1621208567
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1621208567
transform 1 0 10304 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1621208567
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1621208567
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1621208567
transform 1 0 11776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1621208567
transform -1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _284_
timestamp 1621208567
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1621208567
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1621208567
transform 1 0 2852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1621208567
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1621208567
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1621208567
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1621208567
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1621208567
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1621208567
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1621208567
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _203_
timestamp 1621208567
transform 1 0 6624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _206_
timestamp 1621208567
transform 1 0 5336 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1621208567
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_50
timestamp 1621208567
transform 1 0 5704 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1621208567
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_58
timestamp 1621208567
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1621208567
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1621208567
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1621208567
transform 1 0 8740 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp 1621208567
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1621208567
transform 1 0 8832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1621208567
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _418_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9844 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1621208567
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_91
timestamp 1621208567
transform 1 0 9476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _332_
timestamp 1621208567
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1621208567
transform -1 0 12328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1621208567
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_118
timestamp 1621208567
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1621208567
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1621208567
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1621208567
transform 1 0 2852 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1621208567
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1621208567
transform 1 0 3864 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1621208567
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1621208567
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1621208567
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1621208567
transform 1 0 6164 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1621208567
transform 1 0 8556 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _175_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1621208567
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1621208567
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1621208567
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1621208567
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1621208567
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _183_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9936 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _185_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 10396 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1621208567
transform 1 0 9108 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1621208567
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1621208567
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 1621208567
transform 1 0 10856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _335_
timestamp 1621208567
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1621208567
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1621208567
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1621208567
transform -1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1621208567
transform 1 0 11960 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1621208567
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _289_
timestamp 1621208567
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1621208567
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1621208567
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1621208567
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1621208567
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1621208567
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1621208567
transform 1 0 1656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1621208567
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1621208567
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1621208567
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1621208567
transform 1 0 3312 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1621208567
transform 1 0 3036 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1621208567
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1621208567
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1621208567
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1621208567
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1621208567
transform 1 0 4140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _300_
timestamp 1621208567
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _297_
timestamp 1621208567
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1621208567
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1621208567
transform 1 0 5428 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_52
timestamp 1621208567
transform 1 0 5888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1621208567
transform 1 0 5520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1621208567
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1621208567
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 1621208567
transform 1 0 5612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 1621208567
transform 1 0 5244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1621208567
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1621208567
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1621208567
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1621208567
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1621208567
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 1621208567
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1621208567
transform 1 0 5520 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1621208567
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1621208567
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _304_
timestamp 1621208567
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1621208567
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1621208567
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1621208567
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1621208567
transform 1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1621208567
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _308_
timestamp 1621208567
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1621208567
transform 1 0 7084 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3_4  _162_
timestamp 1621208567
transform 1 0 8648 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1621208567
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 1621208567
transform 1 0 10212 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _172_
timestamp 1621208567
transform 1 0 9936 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1621208567
transform 1 0 10396 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _306_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9108 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1621208567
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1621208567
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_97
timestamp 1621208567
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1621208567
transform 1 0 10488 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1621208567
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1621208567
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1621208567
transform -1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1621208567
transform -1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1621208567
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1621208567
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1621208567
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_118
timestamp 1621208567
transform 1 0 11960 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1621208567
transform 1 0 2300 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1621208567
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1621208567
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1621208567
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1621208567
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_12
timestamp 1621208567
transform 1 0 2208 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1621208567
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1621208567
transform 1 0 3956 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _188_
timestamp 1621208567
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1621208567
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _192_
timestamp 1621208567
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _194_
timestamp 1621208567
transform 1 0 5428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1621208567
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1621208567
transform 1 0 6716 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1621208567
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _421_
timestamp 1621208567
transform 1 0 7268 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1621208567
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _168_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9476 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8832 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1621208567
transform 1 0 10120 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_90
timestamp 1621208567
transform 1 0 9384 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1621208567
transform -1 0 12328 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1621208567
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1621208567
transform 1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_118
timestamp 1621208567
transform 1 0 11960 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1621208567
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _291_
timestamp 1621208567
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _292_
timestamp 1621208567
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _295_
timestamp 1621208567
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1621208567
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1621208567
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_10
timestamp 1621208567
transform 1 0 2024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1621208567
transform 1 0 2392 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _294_
timestamp 1621208567
transform 1 0 3312 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _298_
timestamp 1621208567
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1621208567
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1621208567
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1621208567
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1621208567
transform 1 0 4508 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1621208567
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1621208567
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_40
timestamp 1621208567
transform 1 0 4784 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1621208567
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _197_
timestamp 1621208567
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1621208567
transform 1 0 6072 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1621208567
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1621208567
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1621208567
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1621208567
transform 1 0 8464 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1621208567
transform 1 0 7728 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1621208567
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_79
timestamp 1621208567
transform 1 0 8372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1621208567
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _160_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9568 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _169_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 10304 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1621208567
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1621208567
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1621208567
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1621208567
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _167_
timestamp 1621208567
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1621208567
transform -1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1621208567
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1621208567
transform 1 0 11960 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1621208567
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1621208567
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1621208567
transform 1 0 2484 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1621208567
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _195_
timestamp 1621208567
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1621208567
transform 1 0 4416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1621208567
transform 1 0 3956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1621208567
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1621208567
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1621208567
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _189_
timestamp 1621208567
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1621208567
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1621208567
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1621208567
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1621208567
transform 1 0 5796 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1621208567
transform 1 0 6072 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1621208567
transform 1 0 7728 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1621208567
transform 1 0 7452 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1621208567
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1621208567
transform 1 0 7084 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _161_
timestamp 1621208567
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _164_
timestamp 1621208567
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _305_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9292 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1621208567
transform 1 0 10672 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1621208567
transform 1 0 9200 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1621208567
transform -1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1621208567
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1621208567
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1621208567
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1621208567
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1621208567
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _349_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1621208567
transform 1 0 1380 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1621208567
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1621208567
transform 1 0 3864 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1621208567
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1621208567
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1621208567
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1621208567
transform 1 0 5336 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1621208567
transform 1 0 6808 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__o21bai_1  _309_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 8280 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _165_
timestamp 1621208567
transform 1 0 9844 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _311_ PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform 1 0 9108 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1621208567
transform 1 0 10120 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1621208567
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1621208567
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1621208567
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _350_
timestamp 1621208567
transform 1 0 11592 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1621208567
transform -1 0 12328 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_118
timestamp 1621208567
transform 1 0 11960 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1621208567
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1621208567
transform -1 0 2208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1621208567
transform -1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1621208567
transform -1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 PDK/openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621208567
transform -1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1621208567
transform -1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1621208567
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_12
timestamp 1621208567
transform 1 0 2208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _198_
timestamp 1621208567
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1621208567
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1621208567
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1621208567
transform 1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1621208567
transform -1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1621208567
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1621208567
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1621208567
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_30
timestamp 1621208567
transform 1 0 3864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _345_
timestamp 1621208567
transform 1 0 4968 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _346_
timestamp 1621208567
transform 1 0 5612 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _347_
timestamp 1621208567
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1621208567
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1621208567
transform 1 0 5336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1621208567
transform 1 0 6532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1621208567
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1621208567
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _312_
timestamp 1621208567
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp 1621208567
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1621208567
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1621208567
transform 1 0 7544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1621208567
transform 1 0 8188 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1621208567
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1621208567
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1621208567
transform 1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1621208567
transform 1 0 10028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1621208567
transform 1 0 9660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1621208567
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1621208567
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1621208567
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1621208567
transform -1 0 12328 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1621208567
transform 1 0 11776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1621208567
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1621208567
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1621208567
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1621208567
transform 1 0 11868 0 1 12512
box -38 -48 222 592
<< labels >>
rlabel metal2 s 11150 14818 11206 15618 6 cfg_bit_out
port 0 nsew signal tristate
rlabel metal2 s 12622 14818 12678 15618 6 cfg_bit_out_valid
port 1 nsew signal tristate
rlabel metal2 s 9678 14818 9734 15618 6 cfg_out_start
port 2 nsew signal tristate
rlabel metal2 s 3698 14818 3754 15618 6 col_sel[0]
port 3 nsew signal tristate
rlabel metal2 s 5170 14818 5226 15618 6 col_sel[1]
port 4 nsew signal tristate
rlabel metal2 s 6642 14818 6698 15618 6 col_sel[2]
port 5 nsew signal tristate
rlabel metal2 s 8206 14818 8262 15618 6 col_sel[3]
port 6 nsew signal tristate
rlabel metal2 s 754 14818 810 15618 6 wb_clk_i
port 7 nsew signal input
rlabel metal2 s 2226 14818 2282 15618 6 wb_rst_i
port 8 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_ack_o
port 9 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[0]
port 10 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[10]
port 11 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[11]
port 12 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[12]
port 13 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[13]
port 14 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[14]
port 15 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[15]
port 16 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[16]
port 17 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[17]
port 18 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[18]
port 19 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[19]
port 20 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[1]
port 21 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[20]
port 22 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[21]
port 23 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[22]
port 24 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[23]
port 25 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[24]
port 26 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[25]
port 27 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[26]
port 28 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[27]
port 29 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[28]
port 30 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[29]
port 31 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[2]
port 32 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[30]
port 33 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[31]
port 34 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[3]
port 35 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[4]
port 36 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[5]
port 37 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[6]
port 38 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[7]
port 39 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_adr_i[8]
port 40 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[9]
port 41 nsew signal input
rlabel metal2 s 110 0 166 800 6 wbs_cyc_i
port 42 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_dat_i[0]
port 43 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[10]
port 44 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[11]
port 45 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[12]
port 46 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[13]
port 47 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[14]
port 48 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[15]
port 49 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[16]
port 50 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[17]
port 51 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[18]
port 52 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[19]
port 53 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 54 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[20]
port 55 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[21]
port 56 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[22]
port 57 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[23]
port 58 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[24]
port 59 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[25]
port 60 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[26]
port 61 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[27]
port 62 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[28]
port 63 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[29]
port 64 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_dat_i[2]
port 65 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[30]
port 66 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[31]
port 67 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_dat_i[3]
port 68 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[4]
port 69 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[5]
port 70 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[6]
port 71 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[7]
port 72 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[8]
port 73 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_i[9]
port 74 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[0]
port 75 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[10]
port 76 nsew signal tristate
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[11]
port 77 nsew signal tristate
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[12]
port 78 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[13]
port 79 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 80 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[15]
port 81 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[16]
port 82 nsew signal tristate
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[17]
port 83 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[18]
port 84 nsew signal tristate
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[19]
port 85 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[1]
port 86 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[20]
port 87 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[21]
port 88 nsew signal tristate
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[22]
port 89 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[23]
port 90 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[24]
port 91 nsew signal tristate
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[25]
port 92 nsew signal tristate
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[26]
port 93 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[27]
port 94 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[28]
port 95 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[29]
port 96 nsew signal tristate
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[2]
port 97 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[30]
port 98 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[31]
port 99 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[3]
port 100 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[4]
port 101 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 102 nsew signal tristate
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[6]
port 103 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[7]
port 104 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[8]
port 105 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[9]
port 106 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 wbs_sel_i[0]
port 107 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_sel_i[1]
port 108 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_sel_i[2]
port 109 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_sel_i[3]
port 110 nsew signal input
rlabel metal2 s 18 0 74 800 6 wbs_stb_i
port 111 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_we_i
port 112 nsew signal input
rlabel metal4 s 10297 2128 10617 13104 6 VPWR
port 113 nsew power bidirectional
rlabel metal4 s 6556 2128 6876 13104 6 VPWR
port 114 nsew power bidirectional
rlabel metal4 s 2815 2128 3135 13104 6 VPWR
port 115 nsew power bidirectional
rlabel metal5 s 1104 11035 12328 11355 6 VPWR
port 116 nsew power bidirectional
rlabel metal5 s 1104 7408 12328 7728 6 VPWR
port 117 nsew power bidirectional
rlabel metal5 s 1104 3781 12328 4101 6 VPWR
port 118 nsew power bidirectional
rlabel metal4 s 8427 2128 8747 13104 6 VGND
port 119 nsew ground bidirectional
rlabel metal4 s 4685 2128 5005 13104 6 VGND
port 120 nsew ground bidirectional
rlabel metal5 s 1104 9221 12328 9541 6 VGND
port 121 nsew ground bidirectional
rlabel metal5 s 1104 5595 12328 5915 6 VGND
port 122 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 13474 15618
<< end >>
