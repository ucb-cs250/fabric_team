VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clb_tile
  CLASS BLOCK ;
  FOREIGN clb_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 678.560 BY 727.440 ;
  PIN carry_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 611.280 629.480 611.880 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 619.510 680.120 619.790 684.120 ;
    END
  END carry_out
  PIN cb_east_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 54.360 629.480 54.960 ;
    END
  END cb_east_in[0]
  PIN cb_east_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 74.760 629.480 75.360 ;
    END
  END cb_east_in[1]
  PIN cb_east_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 95.160 629.480 95.760 ;
    END
  END cb_east_in[2]
  PIN cb_east_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 116.240 629.480 116.840 ;
    END
  END cb_east_in[3]
  PIN cb_east_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 136.640 629.480 137.240 ;
    END
  END cb_east_in[4]
  PIN cb_east_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 157.040 629.480 157.640 ;
    END
  END cb_east_out[0]
  PIN cb_east_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 178.120 629.480 178.720 ;
    END
  END cb_east_out[1]
  PIN cb_east_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 198.520 629.480 199.120 ;
    END
  END cb_east_out[2]
  PIN cb_east_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 218.920 629.480 219.520 ;
    END
  END cb_east_out[3]
  PIN cb_east_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 240.000 629.480 240.600 ;
    END
  END cb_east_out[4]
  PIN cb_east_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 260.400 629.480 261.000 ;
    END
  END cb_east_out[5]
  PIN cb_east_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 280.800 629.480 281.400 ;
    END
  END cb_east_out[6]
  PIN cb_east_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 301.880 629.480 302.480 ;
    END
  END cb_east_out[7]
  PIN cb_east_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 322.280 629.480 322.880 ;
    END
  END cb_east_out[8]
  PIN cb_east_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 625.480 342.680 629.480 343.280 ;
    END
  END cb_east_out[9]
  PIN cb_north_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.230 680.120 59.510 684.120 ;
    END
  END cb_north_in[0]
  PIN cb_north_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.550 680.120 78.830 684.120 ;
    END
  END cb_north_in[1]
  PIN cb_north_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.870 680.120 98.150 684.120 ;
    END
  END cb_north_in[2]
  PIN cb_north_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.190 680.120 117.470 684.120 ;
    END
  END cb_north_in[3]
  PIN cb_north_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.510 680.120 136.790 684.120 ;
    END
  END cb_north_in[4]
  PIN cb_north_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.830 680.120 156.110 684.120 ;
    END
  END cb_north_out[0]
  PIN cb_north_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.150 680.120 175.430 684.120 ;
    END
  END cb_north_out[1]
  PIN cb_north_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.470 680.120 194.750 684.120 ;
    END
  END cb_north_out[2]
  PIN cb_north_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.790 680.120 214.070 684.120 ;
    END
  END cb_north_out[3]
  PIN cb_north_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.110 680.120 233.390 684.120 ;
    END
  END cb_north_out[4]
  PIN cb_north_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.430 680.120 252.710 684.120 ;
    END
  END cb_north_out[5]
  PIN cb_north_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 271.750 680.120 272.030 684.120 ;
    END
  END cb_north_out[6]
  PIN cb_north_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.070 680.120 291.350 684.120 ;
    END
  END cb_north_out[7]
  PIN cb_north_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 310.390 680.120 310.670 684.120 ;
    END
  END cb_north_out[8]
  PIN cb_north_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.710 680.120 329.990 684.120 ;
    END
  END cb_north_out[9]
  PIN cen
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 631.680 629.480 632.280 ;
    END
  END cen
  PIN clb_south_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.230 44.120 59.510 48.120 ;
    END
  END clb_south_in[0]
  PIN clb_south_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.010 44.120 79.290 48.120 ;
    END
  END clb_south_in[1]
  PIN clb_south_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.790 44.120 99.070 48.120 ;
    END
  END clb_south_in[2]
  PIN clb_south_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.030 44.120 119.310 48.120 ;
    END
  END clb_south_in[3]
  PIN clb_south_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.810 44.120 139.090 48.120 ;
    END
  END clb_south_in[4]
  PIN clb_south_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.050 44.120 159.330 48.120 ;
    END
  END clb_south_in[5]
  PIN clb_south_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.830 44.120 179.110 48.120 ;
    END
  END clb_south_in[6]
  PIN clb_south_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.070 44.120 199.350 48.120 ;
    END
  END clb_south_in[7]
  PIN clb_south_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.850 44.120 219.130 48.120 ;
    END
  END clb_south_in[8]
  PIN clb_south_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.090 44.120 239.370 48.120 ;
    END
  END clb_south_in[9]
  PIN clb_south_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.870 44.120 259.150 48.120 ;
    END
  END clb_south_out[0]
  PIN clb_south_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 279.110 44.120 279.390 48.120 ;
    END
  END clb_south_out[1]
  PIN clb_south_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.890 44.120 299.170 48.120 ;
    END
  END clb_south_out[2]
  PIN clb_south_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 319.130 44.120 319.410 48.120 ;
    END
  END clb_south_out[3]
  PIN clb_south_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.910 44.120 339.190 48.120 ;
    END
  END clb_south_out[4]
  PIN clb_west_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 55.720 53.480 56.320 ;
    END
  END clb_west_in[0]
  PIN clb_west_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 78.840 53.480 79.440 ;
    END
  END clb_west_in[1]
  PIN clb_west_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 102.640 53.480 103.240 ;
    END
  END clb_west_in[2]
  PIN clb_west_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 126.440 53.480 127.040 ;
    END
  END clb_west_in[3]
  PIN clb_west_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 150.240 53.480 150.840 ;
    END
  END clb_west_in[4]
  PIN clb_west_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 174.040 53.480 174.640 ;
    END
  END clb_west_in[5]
  PIN clb_west_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 197.840 53.480 198.440 ;
    END
  END clb_west_in[6]
  PIN clb_west_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 220.960 53.480 221.560 ;
    END
  END clb_west_in[7]
  PIN clb_west_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 244.760 53.480 245.360 ;
    END
  END clb_west_in[8]
  PIN clb_west_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 268.560 53.480 269.160 ;
    END
  END clb_west_in[9]
  PIN clb_west_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 292.360 53.480 292.960 ;
    END
  END clb_west_out[0]
  PIN clb_west_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 316.160 53.480 316.760 ;
    END
  END clb_west_out[1]
  PIN clb_west_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 339.960 53.480 340.560 ;
    END
  END clb_west_out[2]
  PIN clb_west_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 363.760 53.480 364.360 ;
    END
  END clb_west_out[3]
  PIN clb_west_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 386.880 53.480 387.480 ;
    END
  END clb_west_out[4]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 652.760 629.480 653.360 ;
    END
  END clk
  PIN east_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 446.040 629.480 446.640 ;
    END
  END east_double[0]
  PIN east_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 467.120 629.480 467.720 ;
    END
  END east_double[1]
  PIN east_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 487.520 629.480 488.120 ;
    END
  END east_double[2]
  PIN east_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 507.920 629.480 508.520 ;
    END
  END east_double[3]
  PIN east_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 529.000 629.480 529.600 ;
    END
  END east_double[4]
  PIN east_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 549.400 629.480 550.000 ;
    END
  END east_double[5]
  PIN east_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 569.800 629.480 570.400 ;
    END
  END east_double[6]
  PIN east_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 590.880 629.480 591.480 ;
    END
  END east_double[7]
  PIN east_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 363.760 629.480 364.360 ;
    END
  END east_single[0]
  PIN east_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 384.160 629.480 384.760 ;
    END
  END east_single[1]
  PIN east_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 405.240 629.480 405.840 ;
    END
  END east_single[2]
  PIN east_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 425.640 629.480 426.240 ;
    END
  END east_single[3]
  PIN north_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 426.310 680.120 426.590 684.120 ;
    END
  END north_double[0]
  PIN north_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 445.630 680.120 445.910 684.120 ;
    END
  END north_double[1]
  PIN north_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 464.950 680.120 465.230 684.120 ;
    END
  END north_double[2]
  PIN north_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 484.270 680.120 484.550 684.120 ;
    END
  END north_double[3]
  PIN north_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 503.590 680.120 503.870 684.120 ;
    END
  END north_double[4]
  PIN north_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 522.910 680.120 523.190 684.120 ;
    END
  END north_double[5]
  PIN north_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 542.230 680.120 542.510 684.120 ;
    END
  END north_double[6]
  PIN north_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 561.550 680.120 561.830 684.120 ;
    END
  END north_double[7]
  PIN north_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 349.030 680.120 349.310 684.120 ;
    END
  END north_single[0]
  PIN north_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 368.350 680.120 368.630 684.120 ;
    END
  END north_single[1]
  PIN north_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 387.670 680.120 387.950 684.120 ;
    END
  END north_single[2]
  PIN north_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 406.990 680.120 407.270 684.120 ;
    END
  END north_single[3]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 625.480 673.160 629.480 673.760 ;
    END
  END rst
  PIN set_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.050 44.120 619.330 48.120 ;
    END
  END set_in_hard
  PIN set_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 600.190 680.120 600.470 684.120 ;
    END
  END set_out_hard
  PIN shift_in_hard
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.270 44.120 599.550 48.120 ;
    END
  END shift_in_hard
  PIN shift_out_hard
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.870 680.120 581.150 684.120 ;
    END
  END shift_out_hard
  PIN south_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 439.190 44.120 439.470 48.120 ;
    END
  END south_double[0]
  PIN south_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 458.970 44.120 459.250 48.120 ;
    END
  END south_double[1]
  PIN south_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 479.210 44.120 479.490 48.120 ;
    END
  END south_double[2]
  PIN south_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 498.990 44.120 499.270 48.120 ;
    END
  END south_double[3]
  PIN south_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 519.230 44.120 519.510 48.120 ;
    END
  END south_double[4]
  PIN south_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 539.010 44.120 539.290 48.120 ;
    END
  END south_double[5]
  PIN south_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 559.250 44.120 559.530 48.120 ;
    END
  END south_double[6]
  PIN south_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 579.030 44.120 579.310 48.120 ;
    END
  END south_double[7]
  PIN south_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 359.150 44.120 359.430 48.120 ;
    END
  END south_single[0]
  PIN south_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 378.930 44.120 379.210 48.120 ;
    END
  END south_single[1]
  PIN south_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 399.170 44.120 399.450 48.120 ;
    END
  END south_single[2]
  PIN south_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 418.950 44.120 419.230 48.120 ;
    END
  END south_single[3]
  PIN west_double[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 505.880 53.480 506.480 ;
    END
  END west_double[0]
  PIN west_double[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 529.680 53.480 530.280 ;
    END
  END west_double[1]
  PIN west_double[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 552.800 53.480 553.400 ;
    END
  END west_double[2]
  PIN west_double[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 576.600 53.480 577.200 ;
    END
  END west_double[3]
  PIN west_double[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 600.400 53.480 601.000 ;
    END
  END west_double[4]
  PIN west_double[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 624.200 53.480 624.800 ;
    END
  END west_double[5]
  PIN west_double[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 648.000 53.480 648.600 ;
    END
  END west_double[6]
  PIN west_double[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 671.800 53.480 672.400 ;
    END
  END west_double[7]
  PIN west_single[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 410.680 53.480 411.280 ;
    END
  END west_single[0]
  PIN west_single[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 434.480 53.480 435.080 ;
    END
  END west_single[1]
  PIN west_single[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 458.280 53.480 458.880 ;
    END
  END west_single[2]
  PIN west_single[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 482.080 53.480 482.680 ;
    END
  END west_single[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 653.560 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 678.560 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 623.560 672.525 ;
      LAYER met1 ;
        RECT 55.000 54.760 623.560 672.680 ;
      LAYER met2 ;
        RECT 56.940 679.840 58.950 680.120 ;
        RECT 59.790 679.840 78.270 680.120 ;
        RECT 79.110 679.840 97.590 680.120 ;
        RECT 98.430 679.840 116.910 680.120 ;
        RECT 117.750 679.840 136.230 680.120 ;
        RECT 137.070 679.840 155.550 680.120 ;
        RECT 156.390 679.840 174.870 680.120 ;
        RECT 175.710 679.840 194.190 680.120 ;
        RECT 195.030 679.840 213.510 680.120 ;
        RECT 214.350 679.840 232.830 680.120 ;
        RECT 233.670 679.840 252.150 680.120 ;
        RECT 252.990 679.840 271.470 680.120 ;
        RECT 272.310 679.840 290.790 680.120 ;
        RECT 291.630 679.840 310.110 680.120 ;
        RECT 310.950 679.840 329.430 680.120 ;
        RECT 330.270 679.840 348.750 680.120 ;
        RECT 349.590 679.840 368.070 680.120 ;
        RECT 368.910 679.840 387.390 680.120 ;
        RECT 388.230 679.840 406.710 680.120 ;
        RECT 407.550 679.840 426.030 680.120 ;
        RECT 426.870 679.840 445.350 680.120 ;
        RECT 446.190 679.840 464.670 680.120 ;
        RECT 465.510 679.840 483.990 680.120 ;
        RECT 484.830 679.840 503.310 680.120 ;
        RECT 504.150 679.840 522.630 680.120 ;
        RECT 523.470 679.840 541.950 680.120 ;
        RECT 542.790 679.840 561.270 680.120 ;
        RECT 562.110 679.840 580.590 680.120 ;
        RECT 581.430 679.840 599.910 680.120 ;
        RECT 600.750 679.840 619.230 680.120 ;
        RECT 56.940 48.400 619.780 679.840 ;
        RECT 56.940 48.120 58.950 48.400 ;
        RECT 59.790 48.120 78.730 48.400 ;
        RECT 79.570 48.120 98.510 48.400 ;
        RECT 99.350 48.120 118.750 48.400 ;
        RECT 119.590 48.120 138.530 48.400 ;
        RECT 139.370 48.120 158.770 48.400 ;
        RECT 159.610 48.120 178.550 48.400 ;
        RECT 179.390 48.120 198.790 48.400 ;
        RECT 199.630 48.120 218.570 48.400 ;
        RECT 219.410 48.120 238.810 48.400 ;
        RECT 239.650 48.120 258.590 48.400 ;
        RECT 259.430 48.120 278.830 48.400 ;
        RECT 279.670 48.120 298.610 48.400 ;
        RECT 299.450 48.120 318.850 48.400 ;
        RECT 319.690 48.120 338.630 48.400 ;
        RECT 339.470 48.120 358.870 48.400 ;
        RECT 359.710 48.120 378.650 48.400 ;
        RECT 379.490 48.120 398.890 48.400 ;
        RECT 399.730 48.120 418.670 48.400 ;
        RECT 419.510 48.120 438.910 48.400 ;
        RECT 439.750 48.120 458.690 48.400 ;
        RECT 459.530 48.120 478.930 48.400 ;
        RECT 479.770 48.120 498.710 48.400 ;
        RECT 499.550 48.120 518.950 48.400 ;
        RECT 519.790 48.120 538.730 48.400 ;
        RECT 539.570 48.120 558.970 48.400 ;
        RECT 559.810 48.120 578.750 48.400 ;
        RECT 579.590 48.120 598.990 48.400 ;
        RECT 599.830 48.120 618.770 48.400 ;
        RECT 619.610 48.120 619.780 48.400 ;
      LAYER met3 ;
        RECT 53.480 672.800 625.080 673.625 ;
        RECT 53.880 672.760 625.080 672.800 ;
        RECT 53.880 671.400 625.480 672.760 ;
        RECT 53.480 653.760 625.480 671.400 ;
        RECT 53.480 652.360 625.080 653.760 ;
        RECT 53.480 649.000 625.480 652.360 ;
        RECT 53.880 647.600 625.480 649.000 ;
        RECT 53.480 632.680 625.480 647.600 ;
        RECT 53.480 631.280 625.080 632.680 ;
        RECT 53.480 625.200 625.480 631.280 ;
        RECT 53.880 623.800 625.480 625.200 ;
        RECT 53.480 612.280 625.480 623.800 ;
        RECT 53.480 610.880 625.080 612.280 ;
        RECT 53.480 601.400 625.480 610.880 ;
        RECT 53.880 600.000 625.480 601.400 ;
        RECT 53.480 591.880 625.480 600.000 ;
        RECT 53.480 590.480 625.080 591.880 ;
        RECT 53.480 577.600 625.480 590.480 ;
        RECT 53.880 576.200 625.480 577.600 ;
        RECT 53.480 570.800 625.480 576.200 ;
        RECT 53.480 569.400 625.080 570.800 ;
        RECT 53.480 553.800 625.480 569.400 ;
        RECT 53.880 552.400 625.480 553.800 ;
        RECT 53.480 550.400 625.480 552.400 ;
        RECT 53.480 549.000 625.080 550.400 ;
        RECT 53.480 530.680 625.480 549.000 ;
        RECT 53.880 530.000 625.480 530.680 ;
        RECT 53.880 529.280 625.080 530.000 ;
        RECT 53.480 528.600 625.080 529.280 ;
        RECT 53.480 508.920 625.480 528.600 ;
        RECT 53.480 507.520 625.080 508.920 ;
        RECT 53.480 506.880 625.480 507.520 ;
        RECT 53.880 505.480 625.480 506.880 ;
        RECT 53.480 488.520 625.480 505.480 ;
        RECT 53.480 487.120 625.080 488.520 ;
        RECT 53.480 483.080 625.480 487.120 ;
        RECT 53.880 481.680 625.480 483.080 ;
        RECT 53.480 468.120 625.480 481.680 ;
        RECT 53.480 466.720 625.080 468.120 ;
        RECT 53.480 459.280 625.480 466.720 ;
        RECT 53.880 457.880 625.480 459.280 ;
        RECT 53.480 447.040 625.480 457.880 ;
        RECT 53.480 445.640 625.080 447.040 ;
        RECT 53.480 435.480 625.480 445.640 ;
        RECT 53.880 434.080 625.480 435.480 ;
        RECT 53.480 426.640 625.480 434.080 ;
        RECT 53.480 425.240 625.080 426.640 ;
        RECT 53.480 411.680 625.480 425.240 ;
        RECT 53.880 410.280 625.480 411.680 ;
        RECT 53.480 406.240 625.480 410.280 ;
        RECT 53.480 404.840 625.080 406.240 ;
        RECT 53.480 387.880 625.480 404.840 ;
        RECT 53.880 386.480 625.480 387.880 ;
        RECT 53.480 385.160 625.480 386.480 ;
        RECT 53.480 383.760 625.080 385.160 ;
        RECT 53.480 364.760 625.480 383.760 ;
        RECT 53.880 363.360 625.080 364.760 ;
        RECT 53.480 343.680 625.480 363.360 ;
        RECT 53.480 342.280 625.080 343.680 ;
        RECT 53.480 340.960 625.480 342.280 ;
        RECT 53.880 339.560 625.480 340.960 ;
        RECT 53.480 323.280 625.480 339.560 ;
        RECT 53.480 321.880 625.080 323.280 ;
        RECT 53.480 317.160 625.480 321.880 ;
        RECT 53.880 315.760 625.480 317.160 ;
        RECT 53.480 302.880 625.480 315.760 ;
        RECT 53.480 301.480 625.080 302.880 ;
        RECT 53.480 293.360 625.480 301.480 ;
        RECT 53.880 291.960 625.480 293.360 ;
        RECT 53.480 281.800 625.480 291.960 ;
        RECT 53.480 280.400 625.080 281.800 ;
        RECT 53.480 269.560 625.480 280.400 ;
        RECT 53.880 268.160 625.480 269.560 ;
        RECT 53.480 261.400 625.480 268.160 ;
        RECT 53.480 260.000 625.080 261.400 ;
        RECT 53.480 245.760 625.480 260.000 ;
        RECT 53.880 244.360 625.480 245.760 ;
        RECT 53.480 241.000 625.480 244.360 ;
        RECT 53.480 239.600 625.080 241.000 ;
        RECT 53.480 221.960 625.480 239.600 ;
        RECT 53.880 220.560 625.480 221.960 ;
        RECT 53.480 219.920 625.480 220.560 ;
        RECT 53.480 218.520 625.080 219.920 ;
        RECT 53.480 199.520 625.480 218.520 ;
        RECT 53.480 198.840 625.080 199.520 ;
        RECT 53.880 198.120 625.080 198.840 ;
        RECT 53.880 197.440 625.480 198.120 ;
        RECT 53.480 179.120 625.480 197.440 ;
        RECT 53.480 177.720 625.080 179.120 ;
        RECT 53.480 175.040 625.480 177.720 ;
        RECT 53.880 173.640 625.480 175.040 ;
        RECT 53.480 158.040 625.480 173.640 ;
        RECT 53.480 156.640 625.080 158.040 ;
        RECT 53.480 151.240 625.480 156.640 ;
        RECT 53.880 149.840 625.480 151.240 ;
        RECT 53.480 137.640 625.480 149.840 ;
        RECT 53.480 136.240 625.080 137.640 ;
        RECT 53.480 127.440 625.480 136.240 ;
        RECT 53.880 126.040 625.480 127.440 ;
        RECT 53.480 117.240 625.480 126.040 ;
        RECT 53.480 115.840 625.080 117.240 ;
        RECT 53.480 103.640 625.480 115.840 ;
        RECT 53.880 102.240 625.480 103.640 ;
        RECT 53.480 96.160 625.480 102.240 ;
        RECT 53.480 94.760 625.080 96.160 ;
        RECT 53.480 79.840 625.480 94.760 ;
        RECT 53.880 78.440 625.480 79.840 ;
        RECT 53.480 75.760 625.480 78.440 ;
        RECT 53.480 74.360 625.080 75.760 ;
        RECT 53.480 56.720 625.480 74.360 ;
        RECT 53.880 55.360 625.480 56.720 ;
        RECT 53.880 55.320 625.080 55.360 ;
        RECT 53.480 54.495 625.080 55.320 ;
      LAYER met4 ;
        RECT 0.000 0.000 678.560 727.440 ;
      LAYER met5 ;
        RECT 0.000 70.610 678.560 727.440 ;
  END
END clb_tile
END LIBRARY

