module \$_MUX_ (output Y, input A, input B, input S);
  sky130_fd_sc_hd__mux2_1 _TECHMAP_REPLACE_ (
    .X(Y),
    .A0(A),
    .A1(B),
    .S(S)
  );
endmodule